`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K7UK20KtYtnttkXS6lU/HOF4tijgui0zStIRFnwn32o/nJy4DeiF7UrgVMrJTVk7+A/ofPKJFOl/
CV7MMBfZVA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h4IOwO8Sg9A8HxCiUHOwGIlocLGLtuMFoPsY08yDLz8P6G4iVP4wCZCINiI2Ovcy2s/BKa6AfejN
Z8uk4GH2Nb+z180AOljbvsK/28v6p/OXvProHdG7ccqkWT2JsQtIg0PITbcytIUGHdaE4/WfQf5P
dDNP7LLaryVR5VEPDS8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EhuTeEDxaJMTNBir1celk26YZXo7PkcSsJs9NUOhrIutY+aa0VEh7UpXTDCTloUIwVuV2TPlW5hz
RIL1cappTaJtYxpvVfHRBnRTR40TAyoVQbo6UHSRG3gMllC/anoxorL/DGJiib1w/JfXGBdpNnZS
dh+FMeaaJWiGrPZNHGP3j1/dC8zZNp23xn6uNQvlwGcT0b5xEgOcBu0YBh2OAl+do8fBnYORv9NG
SOtzhHTU6Njr9qkvbdwlRShMklfnRPTFuwEG8IzKf8GDzOOQIBqFGNx+CWONzVvAd/HnNJPWDhWf
rZJ1BXfAieMyQSm08c71zRUNaWgpPVYSx426aQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cSSIgzW3p3+9i5undeYqqx+qF1I3mDoYc0yUQlVRs2rl6wBAbEjJqYbFP1ICH6KQqTBM1GmqqZjF
luvWJKGwvvgwrOIcnxcSj+M51LeVXnNxbzqjVasSzMrci0dxhQ7Ue5TNdQdP3nVkm6QJlijfBxVn
UidP8b6S8Qa+lTL9nDs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a/rb8apvM08/cENnRM4KjBSgIf1TnMy9tJi2x9IU1FuL1BLy98OJiPVKhir7wCq8XIwkzgezxN2p
rymf80w7KXDfJGd84a3C+JOgj05kTTST/fr8TAZE6b5jwedG4eCa65p30dzOt7h1WWN3OmpoXpTb
RWCZbQW7uB4dliZOa6P0rwZZD2MJ540cMt8FlzA3MLvAzuWEUfDxZ0rPn3UtLDC1RLWRBhirCSJs
sA7wjyHGaa+lO8qfQjxFSXNmibhYl4T5AT8nNu8Rc2mFror3Sh0JmlRxX7P2jbrKpXYrxLHDmc07
fWQz8yIs/Si3IZTOlYxAZNOdUH615EkP1RsYVQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
E/BcPQTM9nz0M44dDlPOhrv2gPPw1jktZOFR5CDVOYhEeb3XrFzXRaoZFb+UZBrbgwXbvx+a4tB4
8DFKxNb6wU6pWt5yky7YCL1JnleHw3Cy0QZ0XRvMmu7fhf+t47d1aJW0OsFbcUYqP30u1y+xW4QH
fyxvGou/YADJK5uAQ/2vHtQZzugitNwo3aGOKXGGBF9eo3vEURDvdz9hh7QhIBsd8gWA/d0meJP0
RZLEYGuK1Dcs/dmT1CsIxOcGot9s1yE4VicGRVDjaiCKTrZmhiHjkShNZ7uhvSKslweJLa6op5k0
cGrpp1potAm/Dv1EIpOF6Ew6Id1Yw+4z91nlAihwhg8UKy8u0L0/nmeXWoYTFomoe+2R5ZLqSxXt
0nAhdyT9u25TT9r8WEY9cNqZyGandw9w5JlJOPTeoLlz5eAKTKjjmuyhUYlpnyiMlyhB8UYE6uOJ
i+Zv5mLCuBvdZBSMGpF5kY4+eXuBvaCRmnk6hpeFeEzgPLIN6w85ngIQyamcO8TmPmTm/ljzQx1F
j7rVTOc/g8VEBTKa+ogrYDhYE1uMpx3aeEpNRdOSYq+fHt/i3aInOgLk1gpqzujgi+fafQ5K98UE
XAWpzNmp0f5WIJy3IQlUHSfD/n2Jzh+3wUuNgapFHdFs9kOhVnHIw12BF4tZp/MTTj+vVuEhag9Q
GSCJfOEKaPwO/eTlEaBYWO17hHeCvnEc84mwl5Ns1tW4Vf/f7jW4bMekDEw0cshj/NY2Q31YxKnM
xYZbM1hc4/WSZCld/hkBNirFJhQ6Jgn0f4HGSxRJh1EB0DzD2YEzMRx3lonpDUC8CU9NrLzr5LD/
RDu1Vdhw5nmnhizzF/oOm8zBpOdirYDKOpsQTfov79EB+RzqFqrNo44dDyDBGSZrq9Lrst70hqP+
AJQ6J8vqKaZ9ptt76AnSyN4y68tYjVVRnUG+uTNhLrPQMLMHCLx1srqgPe+fvZX5jRUNWS/Svbcu
kBAhQBtjshmcho+Jb2V4L7tBNT2ILfZPrb+n5Yu1Ua9nEE1a6RbvXNNTnCjhk9A8WPay1SDg6RFL
lYWakF+NhzYhDXv5c2WB/58K2SsiyV8mYvYAUn2sCCsBmel6fovb7n75C/YhijkijGXSD3StW+/D
GaaPBYvaKML3aFhEUyJlOa3TINLoEiQVIRaqH0J2oE9tcVk4RGSQN5yIcIFDFGsJF2Pg0Nt2MP11
b4GY9kB5qMnUsKr2DyUVBa4Ebf2WhQ2Lm9JNg7nAK3MinF4S2pJ8RlU/5yu9A5VFuCr/G7GhgwDz
Ac4KUBoA4kNakoOtEewYhDRZk48CVkMbDxoZ6auJ3Jnc84jLnOwn2K8zQt00kum0sUAn16QDGKvE
Qx//+EFw5VsSkIZo8w6MkAtOZPZU8E30y+1gPPgQAhMp61/wbwyC5jtRbSym75sB9Z2Em6i63Gvh
0iObDdbKB8CDa0aQ0bQF+n6+EZ4XUMS8ZSWwhrLkKNEmw6a0tnB6KbpAlaj/5vvam0ucvzpbYoJ+
16PcJtvcq81FPHdV6D0vwRwJHDGtxVEvHZKeP6FPxTPwDrcCAEw9sWw/HY90Gtnr1EjF+dpU4jfZ
o6qRWOdt6q6sA1tH6dkghKBXXulwpVel4HAzw6yTgzYFScYnpWl+1aExNFB9J0e6Clelra0XWYIM
c3PA1Nu5ZjFwns8qLI/nVpOaeFp6rFa+97rcmM0O3m8Pn2SnOWnaG/t7Eyvffu43MVsBqZYX8AaB
LBScercCqB/PR2erTgP4HzRjGVQIfF99NpjZFo0+DfUWYchAiRC6Qb+ROmARlMl+GEiq6yJ2FPFF
r+KMwDZ8Ey98LN+FRwiOYYVDG5TAVSsIxN7KU4tMq2JOhp6Y5G0z0a/fLEoURYw1YSCaainbtXv7
HSfFOgXbKP2lH961c1DvPbgSaNRj6WAIpWWdRWIY/E8Xif7f53vxizVT3rOrqF7bpS/cH6LrzcR5
B8bK4yJeziu6U1pgsSgMuo7QeZI5VM4WKj5iacGdVt88VEW9AyfJJUtUz6au8UM1A8t26Dsvg/sH
nRF5v74D6Q2jYXRWIHIsaKGd7UOfpaRYKBafrg+b+Yv0s+8LCn9pi0u/nM52Pp+jp/Fd6B+vWtXj
oCD3HXGE62D9rIDqpfHSftORDYCex76zyQLprL/jbgeF9mUMJdpPBmp6w00eKKCwzXkWp2G/qCvs
bb7gSIhRYbxb4DEfuIQQII9QsmliKAQrzHJjl2q9CIaC86ipqopXWWQsB7o4fFh6KYZ/WIClk8Zr
JiOMmVoYsrRkc+TQLzuMqnLpblbL0X0GZ7u6OhvZe6zanwXyvB+loFLCeJQN7ysRzGC2zOMuHNXB
dyBdqonlm7c9hxZ1dm9s9ZXh6IvnV08q2QXPsZSQzwuPjGpKlE3F3YpfJ5GxDypw2DjG57B8M7Mo
7y+Yym7i6Yi9WJAl8mFdu3PZBbvul1rI5uwh3kPKz3pu8CAjIyl8kNQavi/lamIq2n+QjCmUeXC9
8A7FOS0SUs7Vw6AcjROWhl5XFBJMpWHaimH1uIUdfZtc2mWVOkJWlhYWIgLofdKSuGnu94DQHaay
dZbIpIBWi2DQstofa2UX0s1bzggWhaVw22JWlW0jkuxdnJAy4RUbcbDAkhYxmdL5akhNsXcOaTfO
E3xGd2O4zVHtwYIxF1mu6dI0iyjD9zedVmRDxXd+AHoi+SbOR4AYr737mQVHIu6Glq7UulyHgjPA
TKvs0ws0raoskFoXGLxU4AMwWIhDZ8KBB9OyWLcLMzsypYF+n9MVRcJJr5l0juyv1/6MdxfZlYdP
U7kVcx3ytaGmpGxa2/h8daqEjHNpgCZW+QNJ6oGhfxAeXCEkpnCUO50ZrvWri67zAoCzBzrKvs3F
ftDtk2zi5a8D+CR94/9tZdPuXtmkMvf/GD/H7+GTau1qnKnq3XOtyNFkWPNLe6RZR9MqVW2rs05A
pJZeXbmVN9rIEa+yP3IwyHbTGapjekKwtxuvKrtYZfaFxICOv2WNDA9a+goalyOTSIEspFH+vsJU
PxzidcI5m/n0WJBxchxBJdLzrHEeVW1oGO37drd55HVPY/nfzp0WasdQ3FAZ1y7aRWSUSOCVahhr
yp+n/SpTl8g9GIH9K9AzJ0PGYnQnoyaOnDxm1ZyQJS/7bbIyxkuH+RlmFb2TC2ywHn1KjzAf1uj5
Ph1LVwRBwLCFR9+RHFyqlNWE9S0fNvZ9dSB9SLI/c3X15RDm6NulNIak3dwtHVGqZZtIGe0YOpLz
HBfFoPdjEF0WkWVPBbg2dddHanO50584yGqjLz3PUSjyeLNuQH93+meptITqK9gmbQ4RekDG6Ccx
whEo894q/dwxd8GtY37hiCcpJUb1FkCzFbPeIw87O29D/XSi9sKANxVQ0OOfHZs62iWUxiJHDmpB
h6IcRDMWW7rWTBk2Tj5+dnM9Nv7P8n9PYomNEjKogpuO1V+Q7aryYnaj7jesC5VkCvpD08/MXQc5
VpPqS4yABn061A6/UPeguDNJraCe4jMiKpSTIade92DQ1CwRjILkdtFERH1gFWtq7PrNYoH+keVO
SLolPoTCAhim9ZM3UNvnLvBBfVogXbB74dH7xyq6nRkOaN8PAkt3vlYFjqZiSAHVZZn58bvU6k26
sA6eKf2uKiF+js8TZOBIyKppH7dv3BlsNvef1Q1hzgm+HdJUdXoeH3SisimweZn39KgC4WmSZ0oi
3R7jTToT3QhCEvSE6MPsgi5j62rmQgEQIOTwokjlSzAcCtepdE54Fu+fMCmUkdweuhS54ciPb6Sj
JwllihB7qcRhCGq4nexmIxvBY4pDy/ZNGlDekKFupL6AWVqx4styKBYbUj+kXQQaJ/xuuym9itT3
dg4s4YJc8VvFNAzH7mSdkW0tKskla8flEtKw4iQqhjYnmS470On2hGXes3KTheTtXaSsiY2DRKMb
U9qdX+Di0LP47LX5qWiyIFp+7c8AjuGEaBJ8JuZJ7PUKob6J1MXL0jowFEh8WgzTD6s0cygX8KvH
K3dZHf/wrCVXzioLw5hJF8B2c5ZltFmE9L2bmRVCg+hiN8g470MfpDVYDM1+Y3wo04TlKh372Hv+
gxKAY3s3QjoEwwgESuBn4DA8jfeychriJpBaRI0Iku2I2YjDdkkrYihuhoil8uOFpJ7A1EW45j7/
PTiwvQstti/PH2c1P0GqmgC5eA0UFb0P8njmIzfvLzSl6Gy3vBMqcW016S8XUR1AzGT3+iU/QbxB
tyc6oRTnN/p4l680d0Q6GgSYC9J4eDYqUX0kM7C8asaqwzXl7DjI5ZfUJqcqWXTGdVDM9epjJD2I
mdKq6kQeYgEO3DRyWkAuhczPbx4Gmt7S7zTp5G6GGss04rA1MtLjmZbUBi3YZmQyRlV4g+iN+1+M
bBJndoKW83szWqyGyp3/TY9poIUQNKt39dj4kSzyuVolqEG9gKGHJvXRKrpJQe/Asva7sr1AEYHm
f5IfBL/oGDa2Duph8iYOd78i+q64L2FZqFD2hn1GPKQZ/J7udkiKp/ZNVuwUTRHbodzn/AFdSCRR
mXcYRlaAn5Q748QvcldbDm/iqG+RuJnpRdyjMDlkjdFTB4DWOuk5K7HjMX6ckDqGQJfmXZECgdeD
3u1TUj2CiXhjL5gPNQrVRq1x5SKhfi0GUuqEr9c6Uya9mCD9g8n1JMOVL7HNf7NV9m8teBE523L3
CRApHnd2iOZfZak7p6JStUmwjnmwNn4e8hJHxAY7V1x5BpA5ZqnLRFwZYbCxCXhWndRwf30F0jTO
luLjDj6ViEFGJNR8zPCcrmWG/m6hrL4/QhkFcjXBznXvWLn7D/CGvGHhaJgX0Jy0gsAMW0IsTjcr
X6557NoJZAZki48CdFQSPWfYFssqI3+GLW0wojb02pW4RFBmXfVwUSv58ZkqDaHdJ9vxvwnu9ZIv
jThm0VRwVXCLbVpacDu9RtR3TrvPKjw2KuBqL2Z9ywbQ7EIhsMSrZhmJ9j9L/O+yQYNBDB7bKrIH
xgNirFeVSub6lKEa3ngBb1vFjBq6NWMsv7tBia8GqpLAyLfYKRxlnbkDwOCkJJhOGhqg0VEI8pA+
mLOOSsX112iQSv2JwBgYOxosn/ZdIGPQMuDLB8el5ULLdZXO6znVWEZOQ8Xcc/s2Ll7/gScRFtYd
3MdwB1PvwWtt4w0c0GD6OXv95yCNEOLAq3zXisNDI0n1X3o0297TCrgSjBSxy5zJG+M1I0TDxCo2
eVPMn/wjnrSsSvFKzGAhoer1j1HLgWk26YWLu9Ev9P/++HTZkaMu5EZ4ZTqJ8FprSIJSYa9vLvlc
EcrAvh8QMWl9Vu/xM/8FaXO4BxOLbss1G/Rd5p3uEZbVhVoxLSzqlUarHR2Pjj57+ukY9unNu3X6
mRlVDDFcLSlVME+L+B4c5ZBinllHVdtoAOdVq6SjL9j60nKJIZpOhF0yThLcAQujyu4dnuYz45FF
VKefHr0UTtkSU4EqlpW5XZlElbpvGC6YC6OVZ5KA2dohPTkuchL3SKm3fR6MXWgLopErihu7JMo4
xhT3Ztu52psKyoSDziR/mvopz1kWY6WuIUoY5Qt/x0PQ5KjimPZ1o2FdzYk4c5R3UbPZTwjPBnlA
QCUCOVCey3r1JYa/hKcb+QUGx2YEtND3sc4WK/I2JRPtLoCRjw6EXsRfwh3rThPjPLN6M019CcxT
k/A6LYWSbK7LcOXrR/damDhsCECmu+bmaKuWrLOPoaJ2xBaNu2krbLw8ZT/NDgI3xKsoRGlHkAow
O85ai+GNMf1R5XETwj0k60OTaeNV/UGDOf/tLlJzXM5kejG5Za2XmcYVpwr4BiUpXpN1hL1VxQ6f
DIoT+dFXiosG30ri26ot332KGF0hvdcX8x8rQKJ9BViBWXIM+zOw6h2wtfIOYFK3Vd5Kb9cjw/I9
JN0doHYKux4088P0NpUeDvPAw2lvf2sRW6Gtz2ghANILOvUl9dznDJOG2mwWNbZVn2E94avLCPwS
bas6BGmimah/ZiBseDtRfD6LP55ET2UTVbGgCSPeK9SKjSkb00hcR3N9MGm+LADnAmsp5UVLbWu1
lganayOX5J4qgWsEDnLFAMTwNY1rJr0tpqggs7aHMDK/CrJCq4dt4IkdQ2ut5HwFgAD0+xNmiQQV
qe1XJqSeOQ==
`protect end_protected
