`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KyfJu81pgUAHlvzi3aEasjHSuBkSGb5D0FA6uzvVMaRIjVZzqhPU5B+p4BPDbnm4/uklhfT9akv6
O7ZwjvoE8A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BlApESOjgmO8NSqY6OV/n0ywYhgUOHl0V/VzlkzJt8+T6EYmO9wqY+yha+1UXffpxZM5WkrFkKXL
BBtVMduncX5Jhqm/tdehp9YL4gr4SWXHfpuSzBUbjkeu0ZOl29mPEzeovD4yyaRnEJNn1AfmnCmY
+VMq74Bm61Yh05bKE9M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KuHkREdcIG5X316TfFUuKN0nnXGwdSnJ+WVOKOLBar/5QrXMxq9gpbCUM0wP9C6vY8+shbtoG0Uz
MEm3r9Ixag7zJCJKQEqii8xJEI9VlzkmX8ZLew/Vc1pN66F2DdMgZ4pd/rLFaEdBv+a1GLnbNG/d
ve98CHIQSg19gNG4Cjbi7WAWUkp6yd3N3ELIiMr0gfx6h9QMtbHXgkiRnYLh72t5FbiS68lFINU0
F1W/Nm9X0mSB3etEErPrIp6ebJi6lWofb9Skj6yf94j9ShgRvX79HLsC3R/VLGCOhgZGdiNaFZn3
8TF+J9IbmIE1ikmlCohTHDcEgCEq0jCGxY/azg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hkMFfpc6MUVNUopcWOgurreIQUqhQBxlUiz1anTLVqxe483foZQe0DPXIMkDMIwP8NWmWRDxkszK
m6aHuplyWkc8NgYZOsLw6uw78hWmc6IGL1j3x0egdtaYzxH3iQPIhJYui6kIbq8sMyccCmp/1IXK
c089H/SubKVp0TOPLjA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pvJOBQTk+B+5JKELSQ0kGPNyoSuapXq2V6QRE+/vv2WxL+bjgtFN3TJb3+Z5qMmKMnNRmxb+/Yui
3iGPWEKONaDsweoAVLTMXGb5lRbFMU5Yrb9rwAf52hWV8dYTp8gc2msctj2QR94p7q+SwbY52jLj
ZVBmNmlmjIEtwwbMVpUmF1laxHpB0cUfs/Rk/EN0m8smzO8QN6AqpykV9obhL6vHIDQbgdIJ9wwO
g49mc7yg7OGJqUzzqXkFQDLNPTL7Obf7pNL8Aau1iSZeZqiwvmm+JJIivenvZ70syH2dJhsotO0r
TwFSa6PEW07m8xNW3Gy9otU6PFl+gdMAQWqnHA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4608)
`protect data_block
9KmG6Zx/RiS9aO9X5Yngd86h0OlAlPgDnFFnfpsEueLVKiDcjzDdufcIoa+nCEnbhJVmbbsY8hNi
c41Yz1prFZ67p/fJ5iGSyz8P/V9WktG4GgTuxR7/+uUyP1T8JYESvLvJcs+WcGRerh3wHtsqmVYF
IsHDH9UrNN58JjUBlNlBIXXK51G5xpBoj/NHkb8kYRK+te/g3tP9btrcpglJi3H+xj3xVtIQd8WK
F9LAMETnTx5+ti/awHxH1S4zj6VRp4K1nm9N0vGnIRvZNJEewjy+4hdVIG+qzZ+FWFNBulNee4id
xR7wyGdel9xNb0Y4zhHnwYGsMeE4SwZSyHy35+U1IeXMRURNRaaZGJecAzyloK81TjFK8Ga5m+5q
fB2wq8oHvJA9szUw2T99ptFpaa6gwCpLo8KK+n5NJDRTUKLUYM2NPTScBb3Hk1NvJWBw/xuAgCTh
OaQ0DKSiZYm9UNHxrfID9fkA2dAJ1IkFwglFX+UZZXvmgAUMh2U4tnMDgvJ+VpuomV2uS+yrapPD
nDHD7HHjKffsTvnSURQBnVdTxQM4PCfupRLOWs8o4rsRRC+49ngeeAn/ADDkxmqAWtW5Bo+uZWA3
XPoLypBzRq/Z7uCJwRwHoV2mbyIXdU3lvRDhs9kb8QteDY8J3IjNQfaQfo+3nqWM1a+wWY5Z9Wmp
+nytDF2mOcrP9OGU0GcB1pZ1hUvrUr6zSaahZgDiA5XRLByAqSbcN1TTcgDutTquF+sgNkcU/BJw
tiH2NgTx6Qp3UCpF5UHgNPZRil3bKtLGNcKVe0TzCKssA5AhHjZyVGrR/4LNy0W783tof5K0eGxd
fwUVlnHWYhY+J97tcYicDzEK82fNIJ9kklzr0gjupn8kOZFnDewToLskCTR2/4n9DNpSrPb8GgTD
E2C5cO+bj/wsd8AvWlw8LmpY2O3Upg5X1QmT5jw++NKbXhf9C5n7uCHQoOtx5GByS3wGrPwoSUNy
HPF3YYekoENPSiZY4VWnawONDwnn5AEONU3sqwfh+ZPdZCO+/iFDaoz78qqM0QORYrjRWMi3LtjG
dWPD5lBUz+KM+mm58e2/x0Z8aHVUB7ej7S5ldlCKNctdVUDXf6CblKGEU/4xkPaDFL7XlGoi1kNP
BxOggLIL7Vt0yhgZd52ttdgvkazsIhbfhpkNvumj8j3QfNZAZWADjWZryWRjbSK8HtOfDUNQ394I
DaReMl/WvmaCVmSUbWzuLvl4StzdsvqHd3geYRfvyp7DcJ03gAb7GIDtnqfr8Jp7EN0roLGki4OS
2yqWKQpeTQmxw/Wgdpsy59rPgCz4EOeCK9T/0kp7S9SaHMeBNNhmyqmKlpFydURWfW5UvYHRkYNw
PQQ2OHrjxzDW0cpmtklJPeWeKlUKl3Xkkj7UyRhUsWVdM0wZ54WVEWX5NforRJDJtMAd4FtNwRcl
gRxN107mu81cKwU7O8lXVeZW1e76du2JxJUAb662++HiV7Nx062TcNpkREUTetzZ44IjhkemPLxW
xl143l+nu9yXqlrXQd27HLIfrTsnY7WXUwYM3a0/sGqf04Qn+CIUPA/8enFz8smPQ6NFl+Q8wrJz
GXOUSiLFSV7xqEpbS9b+7J8y/s7FGcK8JIcCw4L1dmRlXLz67Nd1KIl8v0SGlGaejXRlDh37DKrU
hO+dGONvcxiQFJxxwckjVxFd7N99zo2dX1UuxP0hltcrrG+ZJ0VF48BvKEOoOwrGKGqG/eNQzOs6
DpdOREgVE39HWJTOWTqUNv3R8YTn8Wh99inSfwcdtG+b1ir/Ijuj00SW0QckF4ZQ6EYkC8YaHDYl
YxJLhHRQqmZee72cLX8jxEqSvyiouUCnmEKKEvHRgxiIkq5QIk3AIz+xgorvwrQMNHYjcfSnYZ/D
frUyQTuP/wYbyTSUDwhEVHMo5MvdRdqniDI2WKjlC5u8ECzsjiIu6BrCekAHF9/vtHWFSQX1zZwW
al3Jt7txYTIQhuK32DtLinQdDEPZX87/QnzwK6m4Fpg5bHEaP5COCb4xpN+3vz/4GIk6ShFPu1Rp
IEuLNRtgFTXP+tgdwHCS+MC/1CeDPhXLPCf+v6Wqyw2IVD/2llPpDC4D+FVd1U91pyqotXY7uUR8
ISxtciEPg/5WPogKln9ysCL8KPi54Zv8cH4W2CHt+9Z0jY4j68v8tyZpjPj2AUav48MByrhCh9j+
fWiVX5ITX7j4NcWN0ECLmjOYvooIqLyQ9zsDTK8X/6uMmP3OPWDbdNPFUuInLnAD47Zf2ZfwUO5m
ACCQ0RDrJZzoXEQDjl/0cEuS2B/m3eaoE2kEQ9h9gmgFh9N/yjoBfzvOnFbjykBmghWINNrW5E7b
vcGc6Jnr1Hl4B8eYWZoQUt+M338FJQDWnLqS3OfIcYYZ3/wxURbCvGyG8pyamzZ4Tmvo32zNb+CO
Lf5nZapltrJb+PWWos4koYB8JYV+zUyCRZWUbnHZr/0zpNh7rZPIpJ4AMNss7HlskCqP1YslWiRd
Ze1pzlpsoP0wbQo5Nbo4DVXHxQ3dR5dG19PcbJkuErnjP8Rq0oJlpVKctGwV/SO95/vSogsO1hi+
Xd8fmGQqU+AwkrVm54gFzAeVpmToamQ0JGg0BXeo+2qo5teFj2iRIXzp3iyCwrf3NMMKFiASuQTB
VFYLd/fSgE1xlQ8Rfpc++g5i8jlkkl9hYvnBZpdIhamZjIQEhKRPSyRoQbBFiEBX7ZPBMTZ2Fj06
c4zVAKiMo5p/8Et7R5SYSHVn5zmGtBfptYLnNLHxdwUtdsiV08/q3v2pbSmB0prvhU3qwJzjc3dn
M8QtMg+YvSgUWPyuBKe6sQ82MO3VhAacA7cTYtTR4gYA4wMn8zt6gqiAgOZcUqJXLmHEATbxZsWH
IKt3D/miC/hvoYJQSSb5FA3eT1XtaTH8H3Cto8PdpFHO4wXqwLlRjhSO4HSWlVt3zyMY7K8F5UEW
QHvM2vwVhuaKqEQ3L/0gCom3+9DEZpKQYrkJWyOxhjDcC0Fu/H9YadgHnu2+3LcQc/7i+ndM79iF
VYaWg3zZo1S67YcCjc2lZPPjibgPH8RQ1HpGr+DhzeUO1+QXiS5nGurLRdIRq5JeHK2lUc9rt/7M
aL4uGN4pkqrLc85dLS5bvXfLnvZGVppSsCIKBcftF5TTuFAiYIpNGUqaBlPNaAbTKeTHnNbN+Jan
5Hs8G5QvdQwA4/3lGDcmJGZD34XONnSUcyF2BDFF4IFcT/WmxqEj3bSs+sPxwxQonGS6j1WMDP1v
P8+cAJFg8JQCwpwlP2HrQ3eEFDIUAxlw2SbPxHRvRTjeBDgnbpMQsvhtzDWPOStFVaZ6vIMIOymc
uTV4cxyUysOQBgsKSzlnl3ORCvYvA7PbVjVQcqFj+t595Sh4B8aohm3D4AzkQ7fB5+mriNRwXho2
VuOQhCx2yqJONScTQMr32z1Y8j4vDcmgj6D/nddpnUh4T0zYq/ESLl2wnvagUlWhnfMjw0tyvcly
4bmPm3HWOUCUxvErUeByGYc6+ohJ8xfyEySnMbtujOzLXB8GhTAXYr/UJZmNCW6l643v0O5QPeOD
elfSMTNsNJGeEdkvkgNmkVavCi4vsUCWhqINkvAXYDbJ4u+d7irpYU/sMR/HaSqH/jpHPFfqoqwx
oORmDhvOXkONoySsjD78QJTR2vMQofcbM6KKpHIz7jNPJDWUDk8cSayj+hfoD3Fufup4M96iT8rX
BOT5lChYG4eGxatsNn633n618LNqzSzdA7X6irARZQEYy5qjDE1t/p3cuVklhfyX64jnLdjgOhF4
FYp4lfzWrQrcpHdZcfVoEGVDk6Zb6UEE+l+o/ssPxQRh/CR6uCatjrI90FKE4Eaht/P1s4YQ7BKG
Tp1yJLRuaYSwxp7zmfaMt8q+jPIlYr6UKvl0pSfzgK+od8otjOebYAIFBu0yAwRLr23x86ttAsd5
ONAqL6+rCHfRd1Z/4q714EMg6/WQ7itKvUfVVngHu72BkJXp8P1QQiSG+LHhhpsK5i9Rs9PZ8F+A
v7NVGT5kPYsgvVikVTJjjsALEat49NKCTyf9+vtQelpcumlYNJ6r2lN+PDz3yFxWWrrFh9MoHiHe
cB2gcyrimS3TuapjTI6Cpdkaidajm13lFWIKj4TC1yMNbVYQ/E8fIMw0dDxeGSTqJ9yS6R8NnaFR
35IwgKFB2Wo+ifT6E7BClXK9twqoB/LKCwJLKrPzr6KSaTgtrtA3AXL8Gq7WVq9zPgwWaQROzjpc
DLZRoRxsgODgD9J2+LfHJJkUDaA1ri96WyDgKYAgHKqyt4HKSvxLMZRR7a9jqhfwPiQ//EK8Sqyn
ayT0zr3VNBASuhpOv0aTxh8hht05wo3BgpIrNeRr6GDZyMy+bfX4zinwd90jC/j1ZrL3EPy+5n/E
VDhcVoTBBar+s4Ge/SnGor9oJwqlEnIq2sPW1jwFd0LkxZrlUlWh20ztHodCl2JMvuJjGisE39Dl
4TQFY9ommhqviOvmnvQf/6WWRfEA/5lKGxVL8X1TnAyn7XScWzDKhrWQASZ9PXd/Zr/qswM8EC0a
xTQ7mbJuaugD3lg18i0hIXrNpn65Oy6+/rsA1UaxjKzPjFyzpIL1iSy3cJFtrxZ12YJO8NH36yEw
w97gcNIuwiEhOcQKHW5u0xEP9hKkVg7eXMet+TcXXgfU9XTAQ6d4sjKEM3pO57U98dJMR3yg8LA/
t9yMM2gpkCosoP+a3OH7/u+ZRiQP1WgnJh5aAFqYVc3LjM+Yf0UMKvDC6uRC7XhqkuqAQhJPtqXe
RC7ffOURj/EOJF3Ko/8ZF0HHsgtKF43KU702eWv0Ndx0uO3CAP8KovSZnrVa6Jh/XOp9+TUPWl3u
q74Pka3cvQekfvb8zgSjSw08s9e0DJf1TcTGQhVU05jLjypDzl6imfgAaJox/43ybCFa1kL+loj0
TrREfL6ifAKk54rTQARG5R2ejolW2feZ0+KVXslwoHjjI4stKGRyJRMF6pnnkt9ZjdA6iw0sybei
lFUjXbAGrfTvhuwkBEG40O2xWBHituyRpXyl5WxIA9nrOu9Dm6w9hw3FxUuRF+U6t0NNdgnEP5aM
yh+80rou929y7aDkjBv2k43keEB8wEVkRLEgwTOj14QFfbkWZep+APRkMHgH7McT5l6bRsvrXHzY
/B4yi+2cMVOo1wWy7bb37aOIO8XMl5myXbJxJSI0vSYHHHBe/TmIpw0oJaTC+sRGlZUTFtxclvQh
XckRB35KbTLow5o6q10BL6JcYW9Mo0EZxD/4yeehOD/OKscWDcBB2sRFN86YOctmeDyASzBDy1/d
6siQLbBSUJy/cvn+zMS1bYuFsiQAIlGW/PrWGbCA/74+L5Vgu1nvCzV9jyYghekkRCxeevVNMuoe
djOexHdJD0Ov1r0CvI/5IagcQyuxKxHIAV9Ku7e3SjqrWVHLVxiO/n5R0lgGVQo92w+jSR0bnTXS
BflHZmeKFuaIP/ATjaHShZyBsaWoO2bRE3567gezzjwOFLeZ+Yl1j6PnM/lahEZJRjHqfK4CVUId
LOQ72gE5y1jDkpxoBLCBqenJKJwuxd18AiPHs/Lzg+foeDPIRUN+dScIaYC4IBxFQjTH5tkHNeqU
RNxlmNFVjE/K4yiirQ81MTfBNyZcQE/9X7qIJf95wSnBUaY1+1TG3CTsEcVkQUaracAnaU5O8IiO
nDsX0nBmnRTLTt2G8D0xp23h4u0l4cQExtR4108EWfyCnHXBmp6GJnHUC1IPwxru0Gq9/s7686e2
A4O2IQTnznKD0xbEGtohFOaRDm6BgXojOemA9453QLawZYp+XWpMzbZZXEcMj1QvbMl8waypGVbN
GISGlWIbNcuKtXD5cemch4Y2qTkJe2mNL3On+NdPLd+V0Sn7W6Q8ezbvCJsMtZaS4X07RHXCbj7u
vz6w8/bgDxQeJU90I7aLaB1wpp1tGsQBWigtt7JNMpE/r9dWDIzAnj6RLPyn3bAZ//W/65ZvQ6Fy
nU16zIaZINTHASWEZNfKEB1ZGKD8jw9lSve+hgi2eQyCoMFT71qSHuMO/xC9VqIONP9geJLp9khy
L5l45UIMgVKDesGeyDQTLDA4rp9nVWoexEn9w8cneAFKiti1PCDtOH6jA/H56x1R
`protect end_protected
