`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cxH0Am4zBkP+C1narCZLijksiL8klkxAgC+hKFB4tG2W4rk1gpT/pNxXbk/Bb6VWbKS0yYbElig7
kQl3EWjo1g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFx+ePuBfDCUvJqJJm4CTzrdJYjHmkqp5EWxpVH5z/wO3wotmQ/ZyoxCPZTl5TNO5yya14onLi0F
6IdnxbX7SWzzPvZq+zY1BJSUOo8Sw0gJLSnfRxoO/hQsFydJ661Uexi4ZY+gv4JRkvQz8Pqn2MGt
RKkWs99YRL1lXl8jMqk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I/STf/85I3N3vIZLXFcsdtm9WL1pDlnvafm/pFOWv/peTQCcUNzloUz1RHah80baKyemGJp4cqfn
r5QF6yT/qt3FY8YeJw1S0+iRVhU2dAQWvt4JIQNiSVZsl7aqrXrvZzJ2SlCvL+kPtcOmL4Yf29ES
uAIayrnoCJVAiwJAftFFpjg9B+OjZtyMvQeI4rCnAA3IY2bP0hkw8Uq1dfPiumSIY43ax5DXpZAX
qY7SttiTjeZD/Ca0XgmSGNPopnckbeZQqIck73JjRQLR4aIYeZasDzqFT/2rG41Z8l8CnZPl3NQn
CL3G9b87F9edrEQ9/jO2MbDd3IwwmvfmvEeGNA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bh8Es+1OGPj47kwixjD3thSY3v0j334BVYGfk9zRw/P0IBIHvNGvr/v/n1Y3Q3d0nucjcKTizgza
zXvOiR3fyVlhO60y4AH8JrrZidNMp0WMnstn7dNCtSTOSh9NGY0z+k8/jAXksTkRRHw3qq6xxSUn
5shRFYfk1pT27PEBRec=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WZFCQN7yeiF4TjMUb6/Fblff2REsL4dtOcpOpfjBJiu2yzSKHZpdP8Oza9WDMQn3HKuOgBT6w6cv
hol9x1P4RxQh+0lINRR5jGs05QZdzgBcvPqKzwNo5fG9xEuvV/UxEPSIBrEMHNTR58t6W7ESfJ9z
01/Rkc0f6xUyRSCVq77jEOOzeKnpTj1Q9ku9D/5yvkmYyow66FJFskLQmCUQymXprFzqv/ui81pv
7qsZtYtoZlmkWpDgI/cCQyJ7XEAxXvaamkoiDTZ90xfGk/QhLs2gJHIIruMxCk/jVpswppVv40iF
8IU1LXfqwqOGxEVTOi2XQBcaz4n0CQxy/r8kdQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6208)
`protect data_block
S0jLAU4aAcWQ0Tj6PUC6Bz9hCOvI3ccMTjOtT0rtynHEF0GIFohhtsMmOz1NuGBbosCaN0d/aDyn
3kJ/rxUBqZsr5uPsZVhRnzZKvoAj6VA2zEAXwKmasCv87y1fCHXX91hzTuC2fR7n2Am5HYZjz49z
cHcBgV5KskCCXLo14oyZOQ4I6EKJuCGXpUiaFvAtFVTVnEiuaxMVU1sGAqzYQde3yHMcHZKx9Eg1
c5Frv5aAAtO7eeoVfZMVfexkUpdjDKq1Q4guFdgkUXvGYTuoLuUW7IGBtwKc4TNnSH1MFXIwDcRx
ZiYqS38mQsk/aCMk0EPJN3Io9OuQOciUXlLrg2vlGlmj/s/wM5Xsh4ZXXf2xrZJUppe+UD+Rcc5y
rspYkQbuSdfumZGPFwx7GN/fldzVqR1hGsG7icdlCWwAhd7kEY9QxmLvPuDrMLZnuTMPg/hH/kS2
7yDGXgsvVpi/xvUELj2jTsA6Gy1VlGdtY0o9pFTN9LnO8bmjEsnJfYJnLqJRHeAYPrbbiWVUIOQ9
p16aN8OXzdAsbL44VLqpR/b5w0iKeaJaW9MhcSk2R7c3Ww9kPVS0AjM41GyPjuAKlKSfSZguxyIK
PoPjGqpLJk9jYDsNyKpHyZlOdgHqvm2VjJZApLPj5mYS0YpU4sbYuBkO9dRHC2v4Yv95bC6qlar1
63f3Ky/U7ZpLeOophWoR62WN1i3y5w7DN41Oy4HlgRSy22CRM4sG0yOmMuYxajyo4rRHolVrAdUt
NMH+qcjJ/UGIDs5OEi90CmO9fp1TEEvh+z6geOFpv3BBoUF3sneoPKMoptpdIFWUgNxx0Vldd9iq
mh5KxeBwQ+Pr2lBUYqnHeGQIrAIziT0n4UT5CyAhE/ook7rj0VSiI+WWJIBxjWBWKukOBsxaLHE/
zCcEoIehd7Ifb+Su63v/0QtxCnGmyGJ7uEKDNhuWxDX2j4LMBuLGWagZgwnpXthHRBod6Q1EfoWs
+NGrKJBSRrki0pDgY9CFiggHuIt3gmXz5ad6oCRXip1o86ZcEPsG5Kiuq7PeuPvOaWmXozvWxwjb
IyerGPt39G8k/JiUSS8GACB6xiIaSLVhHP9tQHTs2xh1aj6Vb7eN/ieV7RomuiuNN+Ed/Ml24MKU
E9/pQq6fO0USepg4+sQf+1Qr4lZPGf4kASouGIeg2VhnUiDv/Azm7QiBUCte3Dk9n7EyQwfkGB6C
4k8/R8QIquFxVbSsqms3K7bwludQAcZL03gPFkNcGPvhoUQY20dLNks7bb+iqcU6ueTw117PghII
vZE9NTcsV5c36HBlpbMnfaXQhfTakpY9rT8Nb+0ll70OqKK3jnKMVMIO1tqGGyqIgBNUUezy9YO4
P+bbQ+xqIRLs7uA2hqnv7oGYu0i/kVZlZ12s5Gladl/p3XrGCF3yy7NotrQasKXDZ4rc+GDX2Fyh
5jl9JQ5ewfaggibMUtirVraBSfbYNhAgJTHU7Vsq5P6NMBoG5+FJgRTW4l92Rj7mHYxRnVBFB5+n
N5fyJXGEz4E/bJeCRT5JtbSm+HNG4g3IEVRDyUpS1TNu8dE1POG1Kql4Gplwi+iDwtNJr6yNj5O+
sBwQLo81Ogi72j6wbqXhMgOt+u91vJgu2y9DST5uIz4WDEUg5a2k+JY4+6H/8j+zNv91XLfNGQVH
PpOe0wU4088nzQexDkWfGhOwbeJtJhgpuvVuWClRhpsFDf+CFlXyF7pXujmErTIiViNhWTg+RPGF
sOb7bDNAGKtHO1JzN2izl4LOQo2gi4rPffn3CekPGE1d5qGvmM+VTwAoTFsEqUsv7p9VCWlryVnb
W9hjrnj7BStkjZP28heVKSN8yvazwLE8MJvhyu7W+yNoFFVvs566Teku6ZQGYIPz9MXrT0xrMjfx
gGOrHSmueCsndhzIE/ffk33JHZSrdfx5KhduPOmTKkghfvk6XrvkyFNL+4wyKOpBa36xFgIXO8gQ
OnTIk/tHsLTqFhuxsSHIgiw18dc94/964WXeW9sURM5NlGdxAij01/fBWy52XlpEHuifRz+zMSF6
nDLlRg29+1BLZ4l30X+sgMcGw6Urrc1S6qDxYGO5ionCLzhdZU5S1RgEJN5dJG/D70WIF7frtGlK
L44UuJ10K9PJMJ0rVLLnfx2B1lS9Q/Jp3Rr2OdK75SUM3WV2utjhkdBoQAl4gvG0HXagKjrmHK/L
vsTiKEFTuYmboIn976MmauLJdpgK6VeGyh+odOkAreQ8FONgLUTfOQl0n4dXl405tqp1pvazUw5i
0ijsRUQTS+p/Hx2ZFPuisaL/RGY5KCOfj101OeE+02AR1fvaNm2uV6z65G4dYmYbCk0dxpqyAjOC
Fc1WecS+OvTFCDXWWxr+vzCAH8JG3kU/XW7AvhrRdzauICUc+3iO/LG8I4J1xWCY4FFreI65+au9
X4+3AlcUqYgvsVKAvfEFGI5MvBtm5Uoqy2nkuYYSAnR+xLdP/hwiHOT4QKc3AboPEzDfA4MBODA/
mLkZQZlFgyBJY3nZBDoq7X/mCofzHzC/GicxjqateHku8hoPf1aXi9i9YBpQlMZKY4j+2xT8c8AU
UkrpVTA2JVMEbSGLF6pCmtW1QvcyHltirlCM8sKBA1VQcf30katm6TT1VuJo2RaQm+9sxWAvQJaM
fHUduXJUMKln74t3cU6mQ8A7sYuhWOHkZuvEa3ntloezlPWGFaK98sD/rXl04K0K7z4bNwmr6uOW
Pf+FppEyEXcJIwBaH89ur/S/61soq5fN86z5jZxut7WgtiqllzM1H39p3KCnvGpXKcuEhgetDeSh
UvpieZ1FY1SrLNbHw69lUbZfZzmEqkiCwJ741GZ5IdG12DsRx0Xsg/VQkCsjZpEvdLX0qFLJELDd
9cffty6yP5DbfQkHKGv7RTJ2qi2DFajT0Itro6A6Hs13YG0/Wz2hUc322StwbEiab5dEVWXnlklU
3BGAfnaLGnTSmxAIeCqpMopHTU9c3Dn51mSPN6PPCTQ4M5MfYdpHZRZt8Um4VjT8Nrr7zuHo9Kup
Kc9sZGTAEP1X9/M8PBP/MJzb3ifTE8zW/02YWzGw9mlC+m5ViuXNUKcv9rcvMyovEogIWbpEsUxM
GP56w3VVl1S8oqUuIjhsw2aKHV6pV4t632YWABvVUVW8IvlfoDdmE9178P5D8nWuyMRsVjF/KBvN
lD/fxzz8MT25vBkq3XR+hjeRNq8ulu30nw3N69ElbLgPrR8kA6sbNPRksf9vOl2+5+eDiqoayLIp
Gpl2lP1ZosIZtU+E2eVgwu5n0Y3SE/A2l8jz+hP8jS+k5GCOu6EnVepMsM7nrMFVuaKJaHW2xcHT
mYrEUTFLTlVlm2+1IZpfUIoXayedvcRSPY29sHxCTwyPObnNSFyn1/M04ntnL4DHiOlpdeOmRX4e
82mqYL3XKdSKrrwEGDSkAbYx6Kj0ogmR4JdWi+eZtm8Y1bh6BRnKiRuEL2s+yo0Y3m4QSq6u6JXw
IdCyh7RK4f/fTbLz1HYqo++n3NREbq3rf3zAK/KFbZFqUtUIjK+kgd+2fine+JWNSriBrQZsD8wW
kR7nwC3upyUVam4P2q59aEpj4h44ZDzfpUVVKkRt11L1naZDdSLFmNBuXkxk5QExSPfw1nKJ4WVz
JLA8Tq2HnuoeT3oHPcmjFlD7Aec0wUzYXP49Xq5m+1yQHe3dtu69sToIMcFh3h53YwGdpNmR7ytf
dw3bL61fEnBjcsUzG0VBX5teYfbZWppLK8ASuDtw53PHeDTIUadd5o+sqq4V1pBJeBGiqU8hsUbx
v4oNRDXOnNod+WvAM5E2a7aG9pOl2mcFWQ+/M3kVQvfiGF52RCbkTYZm36TPOsyMtWUvDV+f3/ZO
1wk41caaR7jHEmLLkMt7pXDJEtvsrKo0InH5H4MY1TmlAB0po0cN0BcUFpDEolG/bypbkrqshIpa
wmfUoRbwVe6RzJpXDADF9+diQYOSZ1s2XLDAcdQ/zYR5uhig9soPUSwoZEougoPFpNisEgG/416Q
E/oc6hKHxVcHEVP34/nBFBO6sby9LweepB6sTGU+PrLB7wAakA16UpMCWdqEBoN6ZJzkTWR910Po
pzkU6mUi1/ay34688d9snX1Aw7JBJpN8LRZGVRefmCdh7VqXJPTk2ZJc8TDKi6s381NeNMysgqlC
/KL2GWHnyk+1lk2gPtirdhci2yrVwlBXS6wqI0XcD0SyVgSwi2gd7wIkn5qJObJqi3LmFtgJX0mV
zSE2WCaaGMTYlxJbkL4cxeke8a2MBqBw5H43VWT4Zkk64LtvI5o/LfpfvM1EFtdthMkBrj3dHtsm
x0wY7F1VrgvaAssElb87j8J0ABNwMrsqQd3PHNSE7/D7Z9p6+3CJhLRe/kBAaMq8Wl4l/fIQttgS
oLmA87C/z1pahmzCH31Pm8Gev2YwzPTt/jzCQ+kKacNz2eNErhtEiEh9NngW5wq/5D/5sPQCfjNg
b4WkuEznE15IUej9BZInP3H3jj10maFZ5liuVmCxGT4N8+whyEvxwnym31vBbl1ZC3cL44RkMOQT
VfnvotyI1yQSUmfH1zQ0MlN1hxEyGFBJ2rXiaPwUSzKevy2vDIx4P5kyTI4qXHaF4MlaPsSB0ITP
K1cf5kk8CCsIgp2/2b4oEwlzKw4fuEj5fzGAMzS76cj31JlqAZFMM+NNTVuHJ3wNrqFi8kNO/gqj
FboKMsw1TdfB4+a+ESz0fdyisyXAow6X5E48VgfJZDOV+OJ3aIO1XK+SHqLut3PDRazJIBnqqh++
TsMV6idYdeJnmuQ0zilwoKZlRKSatteznxf5pnGZTMUURhrOTCmJVeKubqZ3j3+0UwOBhWRryo4+
rTq84QG9U57dX080wd1C/XQiwB454NWueRXFHgituTyLZN6fxObdomSdiYWK3VxmLENdnMXBChAu
9+7Yq1us49jFU37tjwOPoCzo/95LrkhmbDJ0sdAKQavIT0sR2Y1DbVj7dQLRodRFrraaAdLEDZyY
0UKhR+I6AqyJWbhAEEuVDFI4U+QzIoesstFAHnARl6CnoAd6vzJ7zuYGxW/BraC2/vkZtRWxX0Mi
BQDCeovtlhWGVVl0z8tGdmiTnkdsFXV7LmeJqVD9Op5BUgd4/ndbKJ9e+HHAueqDroyItFD8UYvr
GlIlHAEjLTo92FH/D8GmgGwXA4Om3eTYfphbVx//WCXx3HGL64NiD0a1kavIXhcEj5ed9+bIOEgk
EiF0Dy3HvRqfm/I98o02VChlXqaG2CKlpXixIpmubRR9tmHe7krbGzXg4De5o0PYtRqyKsYVWmvG
IFtUct6GqA/XqLH+MKBc4dNeqgSgg3gTagzjJ+djgb7JH691DWkU/FRifXudsIrq/Hu+RAgYt6BK
nJGg2cdj9tj9t5iynTv7X5j8TrA+9L14xvuffro7KCw/nd/I1RDdoixlwm7aT7jwZr3mgfTUQ9Qr
XBkodFTtXh2GS+CFtciMvkczusHycbgZ9Q24/s+Yae3XmAY/vYvck0AKch4v8HTKTmUVEn66dBKm
VIEsA+20dEaU5WjHamtcAAkXrxgJUJL8Evnya3JxWL3MwUAfFooO9W87x9dCVWsYohgRALk01IxU
uDhTc0GWLb/lXftnOBku/K3tuE4/iAC8rnbMgoyax1/UqYNOhkOVIC6jogjFvdsVcQWhiHZSewhK
FVGAeGUZWGMAjsT/RKKnznnhdbu9fNxM4tj+Awc7EMRNNAfNOUAkjhHAvbkcvqWk/v+wQO2ko9SX
S/PhrUY1l2APzNGpEeG/YRnsNEp48xpOH+QGWdwYfnLa6uD3b9ZgkXOnoqfQun/U5KNPTQNjUbIK
8MPEri0ZKJJZS9uhXEDiHkorfdliBMUIUxcij7Bp1SGryAejIQqM7p1giEsLM5D4AmSD1+qEtuuX
rB2m0umgygR2hFOt4W0F0emsTBVqbonaKFOYNjgapcIRueR3AwCu1PAm91q3LYV8b8tvRLjxdG0e
psDxoGyB0mX8mYIiM5YpHVtJmlYJ8SW/kZBvPln/x7BPOSgdXiB/k98kEllJb+6i/8x8xWeN/cRe
T22EIxB3USte0PH/fptsphUpBzBkORwfEFlDmF9h2kpl87hOcOT00An6eix4M+X8jl+F7cwaK+ZP
qongH/G+KIISNqGfHBEyXiRIr+RcApRK89u4RqVwXmI+ESLALtuwKgehWdynrQ1TFHgddLC+1QNm
W9/vBG98Ca9aBj8JwwaHix3kTbWmS2PNiK+UCzKn8AWbQU6JJR1zS4YA5AL4I39QKgpfFHmaKyIF
FyR52Lc6hgyZ1QlGV1AWsT626z+CuWREi+TSu8kfYpNOUXqBX1OnA6blBf/nuN0ytjW51KxCltvz
wiRmjmCl9CPodZde86QVyoRr5BfcxWX98E8/js1v/QvYnL2NOitLgSc8FsEwVm9/jFAkEdsVbCCU
6/vkdeJ4j2DjSD+fk96J/1MM9z+vc9VZo/x6vQA3hcg22LkBTSsVcRaAT19829wCbvSb9mqW83SH
z9XrEYBzj/LCasiKkDL4TX7DVXVPVKKR1M0Eqne92m5U9wuoJR8VswaMn050PBcHaruzqErtrnvS
OoD/CSCxbqJSFaFHt1eoKnP1zFyLbsQ0jNMbEF9MEEpeBgPohS+XTbK609P29UCjqY0m6kfSMams
8Y2Pimu59xoSnnX92igNcm4kpcFw6DLWrjmI4qBUph3UwLnffah3FYTJhMHUhpya0+fCiEv6RMOS
qVZOb25mAg/62JV9z088ivlDqk1Ues4DGdIgpzYcuYriTfTSKvEsdnH6Bt8/1RfPrrI2O+6x+XaB
zPMjlhOrZOKyoSgYCMrlHz8TPuge6A+/iDwMIc1lXgrRc7iNuEJK5IaDg13+XRDm3LudJTi/JJhH
eS/Zuy8GWNHvWN17Zs619zYn7z4QaEXUIZYJJd2w/UoIYU1Ws5VyevZTRPeh2VPAMtRKjOj7eEV9
yzq0WHaamO1pS9A8FkBsBRiEShLN2AkeGGX8A9UPFIV9l+CBswzUnVF8wOK2nR7LZS3GV9fP3j5E
gveSwCFyoOWgzCki2IJnxEy22f52sKMNJRIlKpZE2+tN+vb3NlrDVqilwhyP4scW0eTJsyJeSNl/
yaBJ2SCGgpKPcBQnIcyeYmgLov5TPyx57IRE9tQ2W0ReAOcOGrPzcA+tHpGYagFsx+LY3Y5kOBPR
0rY2eA5EakIGVMmihs0zBtC80WDFjZwbmbuQgoyLTcXxdeTkNUnngl4RMmUhht7HoBjaVa0pf7+j
cq/HjaLNr9/sMPRKQx8pwlO2dWecxbd0P/DpUF2VCLso8F77XvSHLlD1wyLrTk4OenPTTM5noqlu
fx1DsOVoK/inkpiEdN11/lSzK9yTG3uUV/wKcJxo8MtPaRPGhIcDTCzFuUsFwxYqL5NwjUr4Vd8f
lifdmbxZZJxWYA6ysXcXJpmi5WarMVbaHpEMk/bK0wZlWvwf0uW+6djIgigLJ4xZ+1+n8EkpwIUm
cb7sHDLjFNBNuudbhuRz1iCR2EnxwND3/Ci917Mv69rv95pmeNrFQg0YdEFdfS7aQ2+d/JSED7lj
LM9fUkNJw1pQMeio3Hl2nwLp2OVrKkLZTSBWyAND40+AO2xMMFa48kp2tiyM+cWLAwyefM7nzTzU
zLehKVIhAnxraDk8V6uelics0bzBt0HnubortbPsBjbYQcOFgV3oSzDEHG2uBtKBa0G9Krv231bZ
PcNEIWdnEDz/96macg3DjzwFrm0EOLKJSA85g0Ix5zpYdKkjskII+b/XslyiTL6KqeKCcM14JNmC
VL9OKiIy0AJITRwSZQKvZfXGenS9MuR2RtQ4wHyfElFplmgV+OP67jahHWwNd+0R3Ix9O/NNYtGD
14hI2Xhh4CeIdP9803oK4s2yPBhm2vPoZBf3O4QWkU/gC5AA3cAulwH5Ma1C9KTBABgQu2PTCmus
uNTZ/V8lzPVS+totysivPxKbg73tWp/NTJNhfelLq39O329Z01j8GkGcTczL4acqytpJHm6bcpBK
sizPe/RCPPPHfPJXwOWCrI2rtvGje4HpR3wG/pKN92AfNbQlofyv6fYcpjnxnt6SxFCGcc7k3bOA
Lmi8gARp/C5BqaKKOh1WizWHiZdI7gYGBpjtyMXPxOnOieUb9+ER1+bOipuu0sC7sE3zHxcDdBWW
l33p39nQ4ehK8rPB1O2QVinzRFRZyyK6oFjd/yOuFXtz4SIaTuNbYYGGvmSli2RfjHt+3g==
`protect end_protected
