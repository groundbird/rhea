`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CUGUdRVD7FXtBGvg1Rll0byA7Oy2SPp9xIaTqV/t3zof+Qz16YLRRFewNukTQ3m9/p2zYRyJjlBY
0E803DRrMA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iapk1SvR6Pf4dAuiUKfpsIGATS3bMdqkwLWgmcDWKH/FT2cNQ/GSUdd1sh8zmVpVyBRaTuqwYTTA
ENmWCRaLp+EbwvaDQm8dn0/Lsirn3ocVqhLCZ1A9mn7puDUKnK1vnXROJc9/8gf0ISkuh7JA99Ez
/xZ8wHGJlTcGkarupTo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c4qOXa+eYiBjBcBRv3cdNbDJ7cCY3r70waoTcG10beabxu5qt+AUtwL0DBEijZ85mf8G83q1PZp6
VVgCxvTJTc8rEerQuFqek0GT6SieLTfTiBZju3pNQ1J2vIhzztrTcXkfEkTdvH4LIqfWq5E4iXX6
3wRyOHGXqLoRWB82Vyad8i5FvCF8dItlcxEFTdvbKXasXDVmHe/0EaFfpLI0CXYYjf7Pjt3Y3vZ3
FIauOSBlerRoBV1r4Y4Nj/CWV2mhUiilPBEqfMM+dg0KEqvv+UhWB03J3tsA6RamG1MyXiicMMup
MVAVXRX4gNYvqgOcBy2zJJzYaZ/bqirSDU++ZA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HIzsd79n6waeEwGnyKO1eFrE0LNhKi3y4cBBSppzOumawbSsoxbTYIt/Mf9VhKc8tSXmFs1mYiHP
kIk34065k4GQ3kwUo85cM5qn+C6vIj3vDu49NY52VXIl9bTHliBHsrgSi1ypREDX86n2S+V14pKX
/aLaoWLj+Ubi45vfmjM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YctimL+sYLCf7oANveKVQ+oaTtZbMjky/qMDvLle7xGfBWlxpUik9VkfpQgo4dovpI77ynimYRx8
slpWCCipfb4lviFHdXMUlj0QQ2FTlb9qaZgHcCwrsXwv15GTi6M1utNnpBgKgW3U/9QgAyZPDqTw
7ULX4uYPub2E2aCLlU1aBhZBBBT7xEkGu/JIdgSmvbWF7MV0Krf3hKh01FHPlxnzD9E5ii0xS9pJ
3xB7sUYYfoNIN/07vFeuy7JFXndd203scNBNDvCQ9XalDPJHwmDOLSM5cU7XkDnJtk+lQIJ3kj7c
qersb7OvoouwraGE0aZQbkf1rWBoSvRiAl9Z8A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7200)
`protect data_block
QzzlrSpnCE2f/NOlXdM3vRV81ajp0+n6qI9r9uYTV2jJy9h4Y2KD2WLWTc07JcgcYfXqP7zJEtNI
/obPZn5i+a/YJbamCoD73ionws4ftrX4Mom+3yV0UBTpMbFk0fDIAxy/oiW7tkc0yUQipcaiE02E
VepK8syk6VRjur532ComFZkk2JVuC4PLNIrMkzoASj6VJcWEA0ZkYIvzhXwKrjzG6y8G7WHpu3CF
zAHIdLuxlHa3sur17evWKV6AGyNIlaR2hMW4pPgoIUQxdHWOeA6OLx+z9hi6PqjCZd+lt81OtuKL
TfGM2wNes3qR0EiLXf5rAC5thmUyQBnHHAWZat6ECSrNi+HCVuMn1v1bG28s3XML5lQoEUmx1dV0
2NJS4vVoG01ZwIazCiO695f87seYe5gmm9YJnNKZdhUFs/17J0LM5FhkUa8zLx47gbJQx4E1HyM2
4bYblSPq/3fkJsO44S9ImbzHPcW5W5IiHTEDFg2shARGql5E5AP8HUR6TN/gOTZxbpqZvX6eE123
74rRfcdsO56/k2mfvi8K74BC09pZmdt2N5n3TVbcrJQgRIyFyiFcaLxH9ArUnWfAQadAxO0S60cf
3138cCiWTgSeo+NZVDUAsveDV/ogEnTqPnGwZlYrerKM6aGTx4K9uN14BBTsv8RveOF+v45JdHgP
naIg9a4XEOtgt3EJuiSYEUXC7OEgkgf+FwD2e6RMPVabGt6Ro6sLSPQe8dBzVwFrfPUulH1BIPCZ
d2MFYs61ol7UxSlBs49+etc+Y7vHU5tJodco0srpgFbZnWbWAG38kTv5cXtzjlDkaaksLUC4Igld
+ezC4CnM/oRnH0yDQR0ZI60KcSAYmIRv2psw5326kFSoofXnq065SUvjN5ry2bxh1pMw4MGTKMef
BczoghaEwoPW2/ot8NhfB5D2YAWnnwHiP3lWu4KIKtrsA/YlCcRCYz/IL6IqFzFWHg2YuScEw9G8
iGepSOQNyFwmQTQf9lYAIKyBWjB7vNhnqSyrHU/kpQGOzR9Ae9ijnEJaIFRkV78+Kw/E1wWql7B8
vwxW323zmRK9iORtRKM2z3zbQt5XEku91Qt3flb5R+pP3LVgJwqtU3EATXbWwj+Fua/CHrjlycRf
IdPxCUuevqai1YXSTiEX9pmpUj5Soo8ezaSGrT13YDatnX660oOptwn5pVCSBAXnNJdbQWvlaBJY
YJn7sHVSYxjiBe6xdtn3OfbdKeWBnD2XFL+sflca6QmjsizgVzFKrxnOr0eMEfnhe5t4iHcWBytF
o8yYVP2kcW9p3IlVcSfbKUp18kP8XRpCbi1VpW4XoXOvagXd9MXdj9TJ+u/9QUsVCX8ZWbEtvo97
AJn/2Imn7jK+WKnGha79I5bALnvgtyfozkuKkNbp/ARepxpphW2nplroI9ZT3ObRxzI/yY5q2Pbh
XA/DAGU1Xedo8BOrOefyXeBVXakL7kv0ZHcXh9b0U7INN2HkHaX24aky45AMfDHej22Pa5ZIonlu
fIeJDQ0U1++IVyA3YMa1wz7ValUP/nYTZx4UAS2zB4pBrMyS+EHVqPL/eSDDHSesx+MQAglJA0j+
1Qerl1lWLStwVJ3ircyQcltRRo9d3BYnbNtSaC8KfyzpH7PggQn6+TZL6MDWn++ozFVtcNk3/++5
wOLddWWcrSVJqKlTZT8WM/dZz2hr0MYhKIWMC7jMgCkUbOI6ciLYKI+3bZhiMjAa7xBiYKFQqT3V
CayjJFuOzS12E84CzBsRyu0YCql+ihGU3jZoYo8e+ss4Su18Y5wqxUJwfKOOEwgz2ujCVUfVHd7U
LcliZfcEJIZv/gmreRohGAhF1B/f5f9z+627qeOSd0Hv8J5XGGPq08lPf4M1KobCG9siejTV0ozn
LRrrxDRpKndmE5IFqoQg133BoneqaisjGrEZzI9QpmP4jdsMoLF5/d+DPEFV63x2g4iVDYZRbXDb
8yHxMiZMsqC4ThgZpnr2XAMq1vEHH23+2K3Y8Ldm92i34E2OiCW9B1D98kw9vgh131wJlbbOzR+G
cJpi+oNktAGqQ2duliEY+2ov9qRfhkadDEvkRtuYdi+28F46Z3Qar1ATNaOHwQZ3ob6r0dnvQDsy
HZmYauftx83XrR6p+DfR4zcmOQd7gp5yRbVmi2o+nNhHjrWy8dPbrJ9JU3JK3PIySXWIKBRU9vaw
h4C8UTjcs7IOso6L/K0bqeGMHSdRTBSnEXpSMUVGRfsGYLtJ30ATUvOJZfrVDb4m+U/tVWwMmMyi
y9YCXdoChyvbqXAnc+wG6Y5mDjN/xSxUfwcQdxiU/3BgnoTTK1gj7CSoq4yS763IEh9m8JmA6OEy
VTN8cdkWlvL9shGPr6HQpzzZPWnyRtPHR5k1HmEzrT3raF6YX6hZUj2SYwVqHJrM8DYVaGcto4P0
qtwlg8aqPCGS5JFvoMkO+n7I+uapr9idg9+Tx2qfge7VV92a2+764uqRpQZskq8/njmhhLnjkmYQ
c/EOaHNGgAmeRBmjZrAOOZI46ZgiGLSpo0rOVfI4JSvQHfHUohkGIRycFFoB88Ok4GbaYRZYRxuS
Pdmc98bVqTiM3E0PmxlR2Aa/qBIH0rEtRbdH0K9QuKlna0c4B8vy7a1sajBg8OIA9x6JgxsOvhBr
XlB5+zF+vzL8Rp2yjxfr4TFVdm+q5f9dykEXmgOgaumLI1kOuKYO59tYzYnrNrGonmHkbGNB68pw
jSU/T/SyDvzJKbCuKl1PUPZTNs8YP1YDKEfSARMX2dJpdj2hv1pN1+AWWbAQWWH0xHMs5Dp7ptD0
Ii9OGe+1ldA5cLSpN/rt8BmWB45aQ9iSj/emQGMKT7yCBqrKR6VLzc4wt3UjcgBdIfFShGqQY9e/
9qM8bXHzICojBDVq9NEMnThyh8IeqB96tFmdxKuolYXVbOx3dm3EB0PKVCLeFzX+WWrd72M3jtpg
dx27akXobv76sIP9uSUlW+9sJjLKDREqvs1uD17gi6ttcTTAnOHYTZyATQMbcftGZizr7Jkcs1Hy
/1gZ3oEVkyOdjClVCj4dX5sC/e9s7aHo2o3fRtat4WQrbB05AVYSDg97nPsUtKs0ihhIfc70iSK/
Ucysrb4vUd1XJZ/Jtq0l0M8tX4inH4zYT9DcxZ4ZLI1RVkpxtwk/Ch5iB8WgpihDiBwu32RRSKsM
gBOTSN77QTsg+1GrVg17KinmKCo74Uc1rWByxVlNgunNphEY1dcAffD6+DGEJScsJUGvmddSNL0i
NpYBFp3SkzoGv/DRp8HupYb4dd0PfeLXoTBzA6NOJx6xg8xfen+97TVRjr1ELAyVSw71PgC6eGCT
BO02w9MKULn3OaZabTud6CIhfSdDOhPEYX1eD1fY20SwGDkjMwZnPTNUIGF98Jq7rAvWNFYbqR0H
hCoHygCdZ6MBD3oqKIngVYCGrVqvw9eEFYf8Bfyb1SyGu4/AOKACIEpomCYyusceGk7DyKtK09GJ
+OsHVSyzMfAPnZQpr1boygb2vxTpd7Q3Zy2QQZiZVSLP28XQw1pEJu/P5g5CvxpcwAtpEGJodbJM
l1oqZxwI8zwgAlPWmfT4ySPdrJnbwHpXX0dKBS8L3cdxMg0Xu7C1qleTcZKXRSoHtDHlbpld610Q
hyVA3b3KHmxx64VvnJpbaiCcNlr/Xt2ogkcEbes3miy5i4lKF3jQR2UlFkAUBN4u/eIxb+yDrTjr
2JkCDLD854FLzMvH+zTzQY6axVEdKqMx8LW64cCIreh6LSBfIuN4E66zALU2PO5WGtqaSZ+X4CyK
aA8EL610OMRJVtyftqDAKO+k6HVgDciuSw1dE6hvwDizFzeolBIFleha/y+TU4li5NnMBqFXnYXU
45sy/1zVAK4c174utMNBkSiwiLQPijwzqOXR00Rw0a+fBvK7JXbe8ykP1IQAbwHWQGDK01HwOBpt
9xaUgIB8hW2caiVn8wyo80901GyR1q4XwM3D7JTDr4tzkzzXdV4XQM6l3utFfToVRdMDCz4H9Gcj
DryAQirpsFFBG0wlwost1/yrxUbIgUp0k+atVhAcIavBZR2bAvjN2/uJMXo7PCGzZ6qr5KVtKrhh
HuugnHk+qTuvt4/5d7Oxwg2C08nvUOllcPbnqiaf1InXdyBXxIpGc0PKiqmXiAC/tR41CmbabYzq
6NChqqSAnG4rkHurSBTv/Q1EW95zg/P1fHEuFOa+f9QanHb7r1BiTbqbJS0A87BwDoKpygrvHfWq
C+6NrpIpdjFCVsXIcz/g1BcSc25d1QEfQuAQp7W/uFX11eht5CtsLumTQ79YiMNPzM/6gN2dlz2Y
F3d6EKmQdMC2Ox9cE97YN53EhFz6xHkt7NUclpL5m4dmxip9aNEY/a13vsAo5mp6VadvqEs/lVeo
LPwQXqE2ur5etrvNtjnbZmfrZyCVIyMLnoeSMJ5S+oYvjID92veCymBjgNTNYCeUKKJt21nbRuco
0bi4oza/hUnRaqOFh4D2YELQIBsz1mpFGreWw04zGrpaXyg2jI+mFpBx1t9U6T3MFObLWCUMHLaB
cxjoH/lgTZU880nbAoGkkI0qkvXr1sX7YKgvwfsxlnYrRz2XKqsx3L1f1a83xNKIZ21zcxbx7bc+
o2w3bUDacO8xDQ7ITlpNRGqgVPYX5dXxHyjgc6XavoLnXM91SjMlta6L/kskKg8PQKp43yFwUA/G
C1XqdAnGYBYzRL6soYZLmKQGxa+O62gymO+VLXa3veCzKUby200c4uPLu/hQyEKLa61jg+1BtSQj
+E+g+Mhp0TKwtbxf5zIcEzsVTO4vTORwdFSbO57gj+nmvaZRvXQ8/Qu6lKLrFBuQ6BFamWat4Ta4
0XOTWYSw2DA3HdOfEjE7Xex4nkaHavYw+8paRfWhvA7Mjzu2HXWyvBqYu6zxvqvgd1Vx/sygF2g+
bSvSo4whXeAGA5Eb7TafvIZW+VupyC3RRUlD3ErHtWKFv46ECZUIHHNu0xdHa0oknK0CQZDXFZ16
6hIkXTUsjv+YQUxTe6/dcmmQRCHtqDtfqptDSTA0xIAqmFGm5p0/8+fKDJC3ikLzXrz/H2p5KUYy
CCfIt8qNwyHio1Ch7qSQz4x3kVc+I5rqLV6q5bf5uPYFoLUocw8UzJfrXzAyrWJrZhgijlOXIos9
9xLxOxDPCsLKtuAWn3eXk+y2DmbdH3Pmsbsg+S7S6KRYfuTSsLcGUeo3c4xsWw/jLlGwrPOJZxdi
/UuXLeuuoKFQrUgVEZrznQQMhgxmk0GhX0FTP3mdgrV1An3BaBjBHSrRTVmi0WARQDoRnARMP5Io
yHQKqpP4TwAaOsdn4wCUi0uzUrzf0AFyVYaanLQYCA0nY+p9Lipl/OwF8jtj+YudU1sGkLC9Uoz5
+gy4RgLqjz8ArKxQB9Q2vODS1bGenoLwQz4yN9IIMLUPuvlDo5zsXwFgRAAaS4ZQPq4siN/PKEkc
oc7QHPGY5DQqfPSXlQTdIExR5Vasjj1e/m4KrBTOfuQ0cmAEXG/OWmrCZwJBR10fHSoE/tFxn0So
jnYQAueuzHmJgbq8V0lAGxS/5WnU1YMMih3S/Kaxy0OaMfwYSjBgIE4wxJEuhw/Rp81r/GN5UO52
h9O8TsQV+S6BlV3oVrRVxmOVoumrfxJu7cRdbOWn+BzbTkgM0/q1P7nwUtpsK4vyQ4pBVW8p9BN7
Od3MJLnFqBqERgvNTm8p4aYrKJwZf8tOF5cGHNgPiPONLqIIPaBb7lrGcHXM3JlUrtWb/zliWK60
fIxOhKHR30HxI7AWqUB+2weYsy78oTESuXgWkwW7f0MQNSRsAEZzeqGg3JKEojQCoDDchp97OafR
f1b7z/I/478htv+Nop38praIfE3pHUqvyJDDeRTsgQKQNtqQvy1Bv+9MM34q6KbQmiN8h9C93p5t
pk++kKgy27FkZ3NhwYv0nEZXVxHaH08CNuikFgZhYsSxB1DkD8LQ62SPufbTikPVA3aYTrmfb8P7
0LvciKeN3Aodo1Dm7BoUjfBupuSGcSdHvJBeVwhk/Sw7+0xLcX9iNiHETf2ZocojdfzbIvtdo1ji
3fIAO1Bq3ak2dqJOurdILfysQ/B0/9SuNny8E5n8US9+TMeTQ25QuBRv3j7i3U/Y2mGz31vwQoX+
UuQThNQUIzMdJa3BJKEHGzgwBUZA3FwHo/l4BSyLt7Cn5OArBjKEj3BMS2je+NmznQCgXX/Hw8l5
jGH63sjADgv9CRpWwuIeMVm1xv6qvwubqZ+cHTeoPv+TJyw9GsUdC1ftrLHfbZawlj8ymc+h31NA
bdsxxIOe/zGj+yBgZN6ZN0dLYuqUD6CbzX+wKHwvucb1Z58bFi4ZdHf8hbwqidA/Jeb37Kt2Ztua
3FINxOo33P5bhPBpmeYbLrh3Z8QfE156nel0Kk+faogdqnmupQgdhhyjpapIKVczDLQ5iuWoIzK/
EpFNkOxp9DNYKdLmYnn8sIYKDr9FQNgD6yqQMVQL4iM6PBArjRL5qHJiB+dhqFXrxL1F98Chg/qB
pyEs3wonatBN8JOPZ5GSpTpmP48DC0H9KrKpVbofXfEH6J4dVZyCn9+kwB0JjCMrrVoICJZAB1lH
UXIrnez5pHDKuLrqcPm0F8NevBrCmwqS6iW0oT1kH9j7AEODIdqK5xFvRCbv8e5X/hryvnzA4w8+
1qACvKfFiS8zYItCa3OR9mhHGPweeH3YXjKh5wezqRCR4RG4oStSRzD/Da3i+SszYKbiO4V5AP/f
1e8FudKrYEb98Vi6CXIsiVEFDSUg2aE+WgwX0NIq+dPWrhl8mNlQZtlktWLph6FD5VSsRsmoFBVh
4DCknLnjSPBsjh0Li9MHiuBROueo1ep501T8lJxXSxAqRdOtHDqh0YvAxrE7J6KiAYjudVUQm4wh
RbexkW7sNU1/gYd2vkkIeQr4qKYk+F0oM8I9eWGOn1Cpeke8VKNcsIdIcMgvP1P02Yk4tnD3Umew
W7zfjYLyolilt5nGr5Z2ji+49vI6dvEb3t6+1TL+hsy0RkQ7jauBh8d2acghXfgtGZj3xvGtTpe0
0mM7h7JOiTa3/GsN5C7n+sNKMP/8byvUjpc99lO23Rax8kTAyKQCf4jmKV2C2e4KUdUcAITn0xYt
7Lbf4ZAskyp2WvsvHr4HQJFOW7MucB432bRJIn23smw+DEeSQzfHqxYDNm6iJqUBKhyM48vyqry/
+UCElBt9YqMHzEYQ4rbUWuljaZXvO+LFldpuVc5dzYan7ky/kiyUJ6CdDOnRfcTuym8lJxj3JMlK
f81ALiwFh6Nh5nGK6z9F8aqlOiaNP+qXXjy3GH/fQAsMVkIVs9mb7GJ1VTWx1ohWJW9ugSK8c9My
ixQeVJRiAPLaw9rvwl+3SxdoC4ON4y9iR+u1NSHZZ06viBvEsGBieRXwbXfeEVIUGflfZGtT9N3q
3a9YZgxXFYa+u3tCvPQStHXCsHs58Ps9miISFPMTsIeRB5x8a+nkDtg3DL4F66gJ/hKikYL8MCQ+
HZvmXdfspuanVkvj+yqlXDi85/NUj3IZVpw5mHhrNmH+P/KyIftLrPAcwHElg27AES0wUavv0Ao/
pxY9kEfOo4kdZ1YEcrGjS4ikcZsBVnloA2MlbDcrQiKyKxlFpkSH/B6vyPpVCO05bF2luZ3oGZnM
wKF/2wv8H967uDjIj+HDNlwR+/EM1UPlI0lkZy6becfIzAm7jPFdimSnySaPPcGLTQbm27NNabEk
WGPR0XUI0CN2f4CuANOENn7cPmjhWHf39XuurMVVGKpS0EbeAu35viL8oZbwlAfJtkgHqNBxveaE
5IAX0r1iZ6QXNAqQsyhyJJ2hUdwxr/xwwfYECL4iV+nvwbWaEIDlPTjeNGQ6Lx0vBkFpwGAj2cF0
Lz6YgVC1thLfqFjwjmCQzuyqQvb53oJelT6O1nTpE9vTQvlEEBhMWV1ozcF/0qrNzDzfKZ8ZPm/X
N+5dZ70XaUMixvWKrrINQrJZMGwNDMYqvXdNbDQnH/MM9EYESZ+7otRbDjmzd6oTw4m2fdDyuyiX
4f6sqq7IekH3MWdpfTs5c80nrMog2mWQ77HRsuh38UC21+zhZxASed5vw6TKsP5OY1pTqISc9OG5
uF/BPC8cROcOs/202Zerp0qlqHY6J/yyuTHNoRzAVetj0Xq1xt2XiqRJ84cqaH88IglC746cyzyw
iFFEeb+9V2lF3I3dwcoK1JVpf6W2DGTnMRjyQUq4Gq7cYiH5aMRv0h3R4zGXb9AhN5jgQ6S8vbFn
dOjTsXJlfcsW+c92W7YAcW5CXHfhuV9J5w0jqxJVrfwKYaxCxcsZELBsS6crb5LAYxpY1NlbXXk3
IO/HFeYo8ciZrjHBwwAg9cZyYIQgvH3pqb3Yscvt5q5JJ9ZCSZDmRMtGrFywwHRwbSP/96impcG7
Bdno2jHg7K/aC5oA+qkhLaf4dfgscRiF2CBJcZ6omtvmFQiqUyOJrDsSjN992FMhaoZwBm/jce+w
PUyoEUgkJDClgiWhayBD7/B+ozMHZXNn/ncPBajmSokWoTpGT6FGRrWFXVuGZday9G6X42YYVEsu
Bf1vAU9vt9TI4lBCVAQcayobMfATeF/Kno6xtaNk2XInec1PCeFqDSGzOwHtIBxkvBukpc28pTh2
QMEsycZ7CdAuWroTJk7JCHD08OjG4NNCQNjb1ay5i+wPG4xjw2lVsDRb7ZdFEBxLoFsPhjH4uSee
InxjJ+au8ixyiemSJUEi1rwtY6puxlzTtumxAFU3HafMiTwLg4MIVitTx09gdzIYlEB+0BiRVG8T
qaoueLUCchNNJIZsCWvVva336h1zitbX7hIbQeKVZISJtkJ9vIW/3Tm7YiCfY/T41DTOnGCE2Ec9
DCGMPSaOubA0teDmQw4I7QOq194Oeu4bB/adqbuz/i+viOztQMHRh4daGnOOwm+C9O0k6dxFqAWo
+1lfPNqUcG7E4Z5pbvgLOubOzWPJtAInJ1L8I3DpapW6EvADg5jcHbRHn97bHV1EDuythk+t8erc
95Z8O+ZBRT6sCRszhBxMeWJUr2S7aQMp8RhRNrUXbp8HpLCkkYAszfAR4HPvOuxsKtUGs4T+gIJ6
RscpyifkDDzm5tjtA3tYNVYjCMnzzie4VrlVkCqT44fFtCfAFpCddFCdo7EguiTyxlLZl27gnD89
5eAGAYAOvcYUX9JjdbFscKT8ZYIZjqDk8DS66soDLfpd+rerv37YK5WUD5TJHrafSkN+cUKJQmQD
1GsW981ivzF8pq1ASzkiH//rsh4/nCCYZoROPFUHQBg/rbau2LpaOdSn/rU502aot0Gerx3wzsNb
nsB+NkFLiPS583dBZokMLHicCe8maPq90ErJP5LcmCzcFdGLowXz6GD+6eLy11RpNykXZytlFSzv
bEBdQnMPkY5S0ZGKiMQJKv2XXIkW6WwNYMxL2/wa2igXz44CQpwiCAeyQzi3YElalE5o62Vi59fQ
ZbtvKnnhP0Ry+DT2KlARuNgiX7IDGamSbSzBH58E+FFWQxS9WV0xa/7FWMvznVt1V0Wf/HwdJ+pS
OJZhWw4jfThJ77CMAiBFM0sQ
`protect end_protected
