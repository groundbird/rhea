`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IhVqKYTaEih4PFXkSsQT2fL6Cd62YJyCkrLg+Z5h2dOTXFv2TbpyzTfsVF1TUje/bHHCm4NBzbNq
jEwIcNN0uw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VsLHX37wAHGF3w43roFVu4uIlvgDCzsirLrNC0Aye4W6JjU9GDFHBSWjGZB9+20csH3IFHZlBMe1
Dv/q+nS8p9PUujeT79tJriAyL69tZzvzks9w60YSBR2MOoc+w9Zht9zo3kBeiWtdxk6Fh2ZHGXHv
HwbgaRi9ebH58vNnYxw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AKe9zWeu4UwoZI8MxUMTWC1VLDqEnc4TuUcw9BTLhBS5XnOhYQvr/kbAxghbcoXKuAoQ7E2eCl5f
K5RGCAkJyy649bs3MaZ03P9ZQbNN3GmlZZlcg66ribVHOnhzoNTzsHTnWxRNoIpi/KB2FArI+0yI
IXLJSpv/JYDewsFetZSq1wI54GnVEIeuAq/gHU74lstXUKQC9gzo4Kwoxtifmr+44k6WCweofSci
IDSgWP2Xw4hGCDFyagZie2f8k19lOd7oMaufKgUFJ/ekOMf5lk6xWfchERcJkQs9fQvxUIWzCEV3
wKKa8wzX/XrLIPK90RC3eOfua7kPN5ba4RU0RA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dD+wBBLi5LaoPZ/V+DWe0Lo9jGJOJgQYS565lPp/JS2mfCL/sUBY0FDPDjZ+4QfyDKFB1ObjmTI3
g6nHxgcBOeuuYcBAGWy+aAh1iMvhq96toRTXfEVxFtbBaYySARtyY1h7EYzRaTmTX6Fd6w8307VW
40GL58RTl05ZKkAaDTE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSTUxKnO1UmpxfBKXCDLOqxLVrJWZBzS4Gr1H245Okw7/pMBVTYmNBYR7ZGIXPAyr3VnJMn5t3jA
uxJ/qnI9dJ9gIklZCUWz2jdkondG1P+fHeNwT+YtXrATstEfUKB04Znpt+62osUS0JmvJhxp5Q6u
Qzaqs1F5JKtfkTnu+ENI+Gjoyk0L8GxnYkBRRdXyvz/GDeysGkvHLV4mt7yI4dh4cAdFaSgnSh8W
q2pERZp56bclHRXQEfefs1adQtuKReHsE5W7iRPWuJZshBM1BR0u6TodNpYm/fMx//T7KA1nec6I
mHWK2eko2358TpnfX23WrEhbVxPbtju086L0bQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
m/xedYEUb54VmzA8q3B/xFIHoo+n97xBfesB440Ls9fujw4U6HrfZteb2aL2JgFOiv5Mt6st0D7P
2YaylPUsFqRsIGi0d0I4SrIfINxD6C3N5NwnWbjuxtwrVWP/7vtKdA4FbDpDYCpI6vEKznKUIVlX
CrJK34usbvIL1YmZ7vv+BIjQsFuvsJgylgT+dkyho0a0wQ9POF64erAjxcyrTPbgAZrGArdaQPMa
3Xip3pW5o4YT2+H0VJZxq/6cwkwxf5aaN6gGcu3+rHWcNpLf9MkBnvi0Qyp+feclT6HTVRsuVIZ4
2bU5V77tmuq9ElBzPTvO4p8oopFcBAZjW9Obt9XDtXLkOXrNRsYqJFLbGstXmaNYp2jU1gnhvO3S
Ake2q0YU3HplkRpvKRPydRKsQOtJMnJIYVy/Xbqf0lHTbUeyoLd6cTZiMVBaiimK90VAYa3cRPPG
/85tIW+kEpwBUWiRyegTUSSVeWcwTq+P1/aR8hygv9vu3A8anWteOQi1Rv+/VL8s+SU2ImcwIPl2
SPq9rdc0eZjCGNOQrRA+rmGWyNFxgXtSF0H9Z8BkYj1IY6F6QWtBlkT7eUyp1CZBbE2HbP5yhzI6
YzOxdEJD6v6SaAU4Xon7vIIrW54BNYhBC54PcHy9M8mwU9Zp9bKXrc+INmub4bXIfuCLVBRx+EpJ
4x3W/jx6XpfSAUClNKtnkEn1ftpOFdi1u61bs0pnSEZnuTiMXR+ihmeUrQMtypd6kWYk5Mjd25mF
7+G78VSs3PLLkwr4HnF54P9leeFw3tRlJcZM323S6jzKmS9eE6S2SnekFz896XUL1sXJ0mvvnYZI
c6oIyJ9IEAnY37C42cPBJcbDhKo2ArWBOYZrjzd60xSup3/UByky+Lw7n+7a9AqjpQrYMi/LpJnz
beEflduZMIKLvbrzZ4u5G5VIEnMcA8RP/khDZfmhDylk2Fu7tubBgKAs7K8zNK/Md7jaOstoWPlY
g3dZMShQ3AUAlGO8ODEWJtjj+QVxoECF5mlGHb/fZWjndKXDaApLVtZe4ERDo5LNxfJhvlHx2LOR
9a4k2p2pAiMKKCW1ekpZU4+EOzcW6BPME23wQcqND3M+79oybvqtKxws4X+iCus/oY1ZLEoZd/JI
3sVXQ2+/1vV3NYvp0RGKt8oMEhIHrpX3yxqVAJ4hbAXpnvXQ5hCTc/tQsDAfbo4U65qBtcCAPVJ8
iGQ6CRqqTSwH8hAUEnrPAjbooElaTYvc1pDcxKhCtVyUOYm/ZSUDcUSm+r9dn3vgmXsNPKKqqmZm
qbD2vq8t+slw8Yk+Sg8QUazhQL2/zhVMUwF7BKAIH1XJvmjx8HtH8qbpDIjphZrGy4gFFsSQCfXZ
G4Gr3cFgl7sawcWbEwfaH8kYq4GARYpL8aC1VXxrctahP1gN4ZyMxB1UAnZcsgnsNaCjylHd4WoF
hLsMiUonqRHsxcjeiAuDKpWBCCZYJGKO3z//oh/ZVBsJ93fFig9TWBJRicrToXRpsDo0RrttxxSJ
wScl62vowRlk3rK6jv0gCs0cPGiS/kx6hd7+9jsyaXr6dGZ61yrISsXJxASQw6vRw/SkR/yhEp0I
HFG1LGjTEPJAGLrf1gPcyz2pZ3dxhzTHPKNRCAvhSV9fdQ6sPQ9b43rWET5ozZ7phr1OZ5KQuF1d
T2ZO7Pn4zeJiAdDMTmiKLxApDQldtZQFNf3otGq7vzdObl3543/YVddYNFi0TuAusPZ4ZKyR3T1K
VbJMj8seiDkKk33oRSDBB+go2dgUN6cw9g9zLyCeGk7FNMPmAqMqIz5A+a5MioVBUnFgybct5ZRX
ppOQCvaki72gXl6mYMRMizZ/TOTgP40Ou09bPvF03Dmdu33uMGOqIVODo3jtRyci9A+YMoS8w1jM
8exYJrFL1bLgY1lqymPJLs5DC14XjgnXXsUATAeBjFYO+Le/8A9JEWPQ8R/NzdhxkdaCkJ+KC5hK
yXsy3tCiRjtO0gY3Pl1Y8AZPLqE5EblJCebt2D/18GJcJPS5pWNy2W9bPYu6xqG4AgtejKn64/4R
eXXa7k2Rk9EhtRgIS3y5czDj323oc+LFDBRnnSlbBVJ5Tv8ABZVVq3YoUlVfKGN7QIzCkaBnnYbi
CsIAoJhzplJPwdp8Ihtk23Y0jbp3L2S6/q4K9mKrC5KqxEqKdoSpvqj4pYc0ck3Y230RphKEaP8a
dVmYWX7w74QIpM7Pv0Sy7qOV4AjNPc5jQKc7j4jtqLXFbd4zX6TCAkLKf/gzYdLwAnaT+DBXtI6R
0BIMFW0f6fQHBfDl7kZ9AYG77eMOsw7Uq6JuDrsBYZ572gAj7hx6W3ez+oiAq68vAJpPXk7mD2Kf
jsm4G1DhLAFmPXLpHkravDe74bgljmDT0M7mdYRKIvQhwv02WN6vis4z6pkA1S7+wKrRYujFExjf
EPz1YdLOW0SPnaPB31cyCJLGVjlJ3cu6rHhzLdtrDu9J2U74bEBHVdvbaMFH1+pKP/9v1xkSJDSy
M90WIv3rfiNgGDBcSn7/FqWTV9FedP4IpQeCnzpZgDbiOJWvmDj1nXIkfaUnrGweyywhjq9hyZcJ
5R357pNur2c3sQOOHVStNuVfUtGRF91El+Yp+JmYcXwJrBrpywj4NXsGiH851/oPQUQJcuVcL3La
/04oXqEdTCBbyAr2yk1wlcbxB/1Fy8A521vu5sR7Z5slD4TUIG+Rw8vskABtaIt6+OylTAQiEJMx
kzXHUbsWrvv0oxHQniqVPwkxrbFXfJcrRv61Tj7oO4uJP5KnIOx6ii7iH/fjLchgfnsaElXcAH52
r8tiq43+dP4yOQfGNSWrI8dz7Nw/JXiytuOEHaCP0HzNYgmPM5EMzNHb51gmUXDAHg0wLEUVd+Rn
+tvXMrREcDDWRkWey8LntVrd2PmlBpGNWmAKrUpglQ/0IKbv9PHrWptvvyBxfwNezmXDst8b8RO4
3TtgKoqJvNtNlG1hp8UAAT8Iyeya0UVMNHFasrS8i8/EKB/gQGK/MyNd8zPROcyjENbi6IN9mrTQ
TX5/3oSxS/5Zl+ae4CnmNe4h+IrZ4kAxAurkhAY38yK6Goqt1DlbRD6KJSsyhrdhHWRcwM5f9R8d
zVRVujKmRivFHXS1fD4wY35ZrQGBR0BrvpqPwbMNCoPAwum/Q+A6Xp63pPCdwsfcytPj+ewlhKJ5
+qx9yhrQo3Fn1gG1sUV9Wn74HPb0g3iSmWZnrg2dnhtdjDBd9LCk3QsR1i+0r7s40kWAjRqaljeq
LFk8zAZar7pP4JNHCR34hNxcAGD4hL9ElqD7VPYVVMMjIn29Bg70fe+gyJgZwHHI9vnJfn6qsot7
vRfjtLlbfKnV77IDR927nwhdIU7jLH8j2wW6UCxGJ7l/co77GB0d9IKJv6Rpx7s440TvtW8E1tAz
zQqh+y6lfBhZpGEGrYy9oUvQkT95EMd6+4eJ1d+lMiEDyMjEc5U91sbmC+bydNcdIN5/imqI2LIh
C0YDkLb04XgGEc0TENiXjsEMO/XciKqTwLWO3elQTMEAmjChAZ5OdYoJZhvvfcyacLBdJJV8bV7v
dclmAhWCGRlPBjAnrftvYG4NxFaj3Yz60GtIthBe0nLpze8zZXCZe9k0NdN7V5T8W75R5DBj2mzv
YFJHnToNOpB+1Yxiq6iG1KrN7dys5Mt9SXAGBUeGgz26oZ/sbcE7mI5TGOTBq5tWw7MYgdeF9yDT
7DfT9bObEYSWjkltkiw2CjXq0QjxZUEW+qmqNFfst+YNNNuheOZVxB41PKVbfD2e4J5pVEWaGifZ
dDQmKZmPTi85afzrP6vytsrWLs+oRQnlhvVFdpWdOmWNS+A3dcNvkH1uYbcyeA8J9tz+TYbQTiEZ
5hDn7kaU65qUr6Rt10oGOnGtK+A2V4uykpz/womPhdBLSjPg5ccwBFftphn/WDhOR3jKJBw8Rsa9
CiVAY7Y+6GmkINUFAYiRu2WUXixYqMK8VXRels5JQz64+03nWltQeim1jQ6F4nIDapmNHXr+3hZc
JNAMoM9ypJmFCtqk/tx30X9wQik0Arno6QzKZfqmibiAxPiyYJFkvVR+IFQdbBYZ+unTCELSoKqZ
v/IpyAF+fUbdMQCnGFGzGoGeWnQ0FcqvNDYA7X8QJIPNbr4Hyo6Nmzcs03PDAHRMWzAncWtfgMev
5Ak+tkldnEGQezeM6eB7GiJsDcW8nP43T3vweWPjo2lSFoC6rYTU1j20JhU1otoU5zN+5jUubXea
QDaZWYC4IIQIcF66xHoo5SgEUJ1bJKVBLUHJfohZnqnBCU2KLVRrS2EWx19nQT132sL7GOBL2ebZ
mqCHmjVfIlM5LvGFepLT4m6FCI2ffVSwmd2oizj6PxBCLfBtLRYko10+IsI4riYrUwWe8rDeyxvK
QMxDt/lYz2t2G6vJHecAQEciPrJmCD0p+vOxUfk2DLXPhXBB34ujAL2jiORJP+/+v9BYXxrsaKuq
uof5ImEf5DCa/zvFgqZHDjCPSqXO2lkPgVqs/TsrBu01B/3XDackbhI56/vd7/MbN7sffqRDLQX+
Mqo7UzrdpAOOw1wiqB7HteQRO3ZPoKxQARAYJqjYob856eQDNqf+dBUmn5RMf/WQZWucrj9j/9n7
3SNTImcNSlB72e77wAJn8D0mbPJRbPrJekLx1/MTEJ8xSVVr2ToHwlwF3N8px34kenBkEpLGcGij
YIS8wVgwnHJcnWjJBhNxBxQaiy2YgJjuSaG+Kb3gmucZSS/1P8JuOr8Yh8/LusGftfHwbIMRJV5T
Uc9GfGppKAQy0Lf5n26miTO4ZlvYyg92otBVH5RVYCE/7RmefuFw55GHonGTNFP1+PXx5kSupb5b
Vc6amliSXATc9U2oQQ+iJmxkEm6PNgEJLgXmrKkpsQ9OaH0NCT1fnFrmTblpNSE5jZieIanQ+vfR
+i/vXSsa3AOStwbNP/y1hUf9KZsAQY3CSaP3tJUg1aTZ2DA9uosb4gstAdBTDn70No48rGXByF4L
0YGxftkass7EOI1bjDcywcCAvRhcpaO5ZToNzvsZTO3pwHKSaVG1y9SK2W0w3hTPgy1adBdOlVuS
Wsb0wnNo72EVGHxqShKr8aPVipg698S19NSekAnkJFVO/E1x+ZK/zqr/750gESuzxBcazYkaUS0e
V8nPaEhHCR3tqI9oh3zQ/NmA/YwlENGoYHkhJHJEYnCiSyOHVBTuAc/WD8ooGGbbR8BZwOnJwRn2
Hu4bAarp29Ga7jX3w/Q4XRakj1tFEVWE4mAlQMaPnwOjkkoXH3ecD42SD9iAI7GpHK6uJbwN5+Va
BLEch5N5nm6fWDLHSth0dBO9UjsiagGqDP8=
`protect end_protected
