`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VSnujw2zIGakDZtn+Isu9FyJeHx7Pz8U2bDtI3TDO63118cT4lX4GS/uUF69tsNeIYdtqQWMa9Sr
G3SXfw8DeA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M+UNyhXCe1hknfqmZ0Dmh/RIXszbZSHisHMiBCqJB9Z6PJMcE60LpusT5tCtdf6W5KhXoY6v3h0Q
amycXsXtaQyVn6ZnxhICH/rj0VMpqktxgfErAHe+0hyFYgUz5xFWC27RAbPLw2oMiGOks4VVe0nF
ELLVNDS4U3svrFtI1nY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EXfXHlFt7UAG9nwAKAdyJgyFpGU7WG54+x2bp9UMkt5mRjtv+A15WGAITbQK79Q0NpyxscIazDIp
vrfAF1mbrMzzg3wngBLvsc8GDIVElgZ5A1A7PZB13VyoO5H7qo5OK/xanPESIxFNfkTQ92ENENe/
cHToIJ61p/3gAmJwuKg1t40skfoLrJOHVpqOYl5HKIzxaER2xHKnqMJN/lpDHDCT88bOl/rJ4NJ3
WiwQGwMkfdvzwbZrx8nOTHC++BtESrmxKPgt+QxjXnApACHr/aBzgYaELqyFCZ04Q8WVJbFdr2KP
s4/cbGZOkZSUXsiLPz1es9PBaSw1IU/uypt48g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sfBofOCMECSFGZnGCAwAX+n91KylIDX7mACGkt6LCBWJJZ2SGnoXy46k7Av0mlNF3mrPNm04mCs9
E5ee0TCpjDlIvv+QfgLVAFJMBsgo7QXoBn4JKb47gO0arxdCt+aacglAC8RfEHuQpTEbFWvSfMbW
IpX5Gq4FkV+pMLRH/ZM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pnUMY1e51hghM3aJ40NgTx2kb6S+CLun1HjPAkgMG63GP+mGipqD7mGB0G10Hk7/A0Ugl+/rgah/
XvEvJcUwMwQxSULkpuDHQq842d5l7WIG4Hnoy5kcct0yo2yv9n06RCq+ViCMoQQzrk10ZMyK6s3A
TPYi5n5PVQ2n9lNCr5MAu4eUDBTCPsIHBXJ4jT6eZQfmnWTwYq6I+zxac3R39Sm4tqnWpQQlz/20
XwUylcTkjZNZEU2nMuV7hJWZ/XixLw7DwlEWIiC4upQAYZvOLS9jtf05SChws2EOjQKFSC1uMPNM
UqA9RSRhhG9miyhCMlWOO/EIBgNXxjDOgs2VMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 95680)
`protect data_block
lbLQ/X2y1BhIjtpsI6iSYEN+FpLN+E2GY5ULIpG8+o8EM7sTeOXmwKmKvTMuNCL52wxCGZJYGmb+
FS9fHn9il29VHWdK5Epz6s62czwsB0GxECW6quWlRGUka0rwRo6xn431qoHyq5Of6oGCgCcThfwt
pjcokpQihlIemOYmVKPJOtKGN4E5xqwf9qNsvhrN3F4uwRdPhK1CWwh3w1rmKwVoy76CqaYCDins
cyFQUtHXZHoeXsITMAreFOargjyrToN2246KuUSGHEbyEzviTpd90TJCkoqrF3JuBCxa632jA+3M
ttL0ezd1DpqO7DMALMFaxqjW7YM6vx5D7yO1ewMnsDRdM/Q8NoVlJjnRSQvFIXl7S4Lqkn1C2qYw
5ZxyL5BB4VPn0Gd7utmXLxzzyG3x0RKmoe8rCHA2fOkgg+usp9IMpJeqIIIlIoN1zOTT+r1yjWqH
C3o/jl4hdHvhfOT4ekhNNRgccuyGSqC79PqOQNvZGAIIlpxj54yLg5jZZhJnA14czi6iEzBwq82s
BMUDDI5helAWQ6f0NF10TNQyqMEaxJoUIla7IfQBp31aj4CJh3tiq+cmkk1ZGEOodDWX+de8K1S4
GwS9iiCLSN3oVrrChb8Wb6gB/xA67qsON1otIBhyz3JSz4Zz9sPTGSt3Y15UMSi3y5A7I1Eb1yE8
X6RgGU6g4sSkA0/n2NPmYyWJghRE6ET2IhDkSD0ye48FvL3GChNOc6+UyZK9je411GzoeSxLF0GH
L0dXyvmk4b42FoY242nC3fsXIDupPcdAcRkWpZT1gglunniGXdLhYdxtqKUeh919L5WRWWNaisXR
xMnZO6l/n9ZhQ0tFdg+pVtShtP/V0Z03a4FNR24XteQS/KiEUpIci1ivguWAIgGwh2ppOQTGN02L
aZTdtys9rcwAdDx2IqgZp0ZagbFUvWtHKHbrxeZ2p10egKulU+jAiIoZoHzJsAbxMqAHeTZwckAF
EL2/LnSHJqkWUxRW1Jv8RzkUMeT2Wq+X8iZTJbz27B+8k5MpLzMu+prHkDEnGXF7plGzjCKhKy0w
UtJPZ+4/3yFqLILrf0lRgKBmcSre00ARGGBw6bVrf6xlkmecUzQ/yn9WjHFXMtlTsoWMyNrln+r+
b0U8VbgbqCjXsaj7cYSj22/FQknjx4pxTJmdc7HXvd0IpMKklqe0X5AtIFQAsjKInOtAr9hBIVks
8Ei6i/ekvigzJggsMPCvWsppuepjzqMepDRNAuxuslOcDgLfhU0f7ZfSR5QP1q7QN43Xr2fgfxPZ
Zk1zkJFquZZ2m6LfWN/3WaEQCIqio+9quPCMaxyhH7Xy2QzR0xy/x8I6/DdDv6x4hicGRnsdNfVl
HdBokB/hZ7nmEAK7c8IEZFJnnubW3rUzADnl0ay9+M1bTCLYdg0fLBfqS5klPpb0iNSoMwnKw/5k
riUUFpVDApzjRAnLVTYb8DpXpdvawyPN5+5lHI/9eIJd4Z0U0xrI74HBeEggKl+lr0CPeN3i8Tur
SrnP0JwVNE4ZsQmlFfakgjU/9Kj/Ry0dWngeSpSd/ewDmiS3iurCISyJoTN2KCViSNLKHMoapohh
TVKKlNgiDoTe0y0VPwGGkUNk/HXJbpEtmCoDWAfBt6bAYlIxsYVDv6nPE6Berx8sQl2BK+VM7g25
VsqCTC8NTeq6B8t70u5rlZgEuOlBYKQ8l69T9Y4WJzf23OZcVulBX51G/FlzYR+8Vjq1wVbn9rWJ
D4rB/Pruto8zu5t5q5vbOK7QOxxkPsXbP0C/7QwtYMDazdcC1TOm7PQypORlFvZ3izLQrADwzz5x
4ebB5wysCMhJeoe3LaB2rugi23YJoauHrpr+YVkJx7zC07JSm/vcJAnEHGBlmt2JBUSSDLMMAb3u
9fLp/IQIFqdF8DCIzdjkD1RRfZnxnOr5sJ54Jr/d+hPYjDTXHjyQ5EDFtNrINantHS9QPiU6dCkC
v6RI4xq+qqJzeaVJxJ/P2ko8odohPVEKcGSayhLxdW5VwwNem5iHeqsd8xocOJa6ZVJODljNQsTE
4ydDb3jL+DDuoycGwEAyw8eNi9BYa2iy9FcmoClZ1ZyHVbMXAubo2DTGvdxBGTrmYZifcsMTuxrf
06TEf+L/q4nV/Uf7632UFXpdfDRIaujwciZS7PadSOFdOW+juzPexwOfxwOsWPzTVG53tyVpxx5H
T+hlFJGiGs6R+rNvmc51B8C5aVc6gmw8UMLV4HLI5njSYb39VHW6Nq0Zc4P0bW/ma+TinhiB9RFJ
XMScMPUEZ7CpNNaeQ6sqAeobhrhPIa+QIKlFSpYD+6+IzP5nYzh4bxGXmgUw3Si8THGVy00iq+Tt
qR9WdfVBzfEZaoX+6Hj+26wcI0XmQzD2p8DccakCbg39Cvuk2YizqMorDYtDa5ju/CGT9GFD4Fx9
rPMd3mjXGBIPYTqH1Key5uPR00yr6uKR1UJ431bipC51UGH2B00GQmqfUK9fMN+Q7nXQw0AIgsD5
zCZAm1s7+v+uxWpQG6owIO4QhI+8UXNqCndHzJFHar1CH+2xMqW+AGp3gC2CacJTUFInahPmF2wk
aHpgZjGHfp7/YKbuRW8QssD9lKv4U/PNmV55HJDCchxRzZaS+tQWg8Q8sL6yRnhfqciYyher0/wE
XD93DO/e6+Gj3rzcW2sc3O/9w+Wom8N2FRj2OBwUX+i9RxdMtcAWo9bxjpZn/gJRbxMH92j7J47/
vRAyIbpB5T7wScE12gWp9En/SzeJnDxzgNYdBxoOuclSXv4m1oHJEZLe5GzC2pvUkBQeYR2cb2ix
pWRQcEiIR8fGJNglNE74Y3Lu6SgbzaS0EUi7mZkVHLIX+jBL3lgaInbM71zuzRxO3HqE2eyIyDzq
Ge3X7DccZI9DPDnWLLuNVEjm2MrLaf0JM2QFNH0fvqTQE6ErnL5pRPzl2m8ozUqJeQjisJw1huGT
5C3ILd3iNEEqGZvUI20pBJrO6LnEP6EVpwGCy0GLMhYM69ffG3XonoElQAl4wy27XOlyK7H8xpnU
VSGIKs7rGs5ctNcAw3q+qP6iX/shIgFVmEXL2hDu7WP9F5TTCANRH9CWPxcB2Vw/9V0+2sGv3bWB
L77cdKW/CU51sVyjr8n0Xk+r2pn5s2zZwg5k1II9Z2iu66U7WLFmHvsap8M4MwAIvCtqYu++GimW
DSrJp3IBLZ02ul+miqmsMDCCJR/dw922gjKcEu4AyT8yR+EZfQauNFlbPF+zsD+KTRmVmRXs+5zQ
Ih+/zprLcku8arcs8aCagrxrdwH2ksUrHQACOTFf0t0BkEdgMnovJgX+egbpg+vnRbXq88WJG7Ma
ra0JBr816+kjRpfwW7M83D/VU/kVTZLaYqK2pObPneyW01WGa5gausYxPnNEpXbgT1Bkd4jaVT9G
jGUKe7GQ0SKt17bqJ7DXQEgiHz+bjvFNdXsboEis7pHRbuf+wmGjCyIa2fkK45yTd6FTaC42Treo
L8xayUkj6mDbEDG5OBqXIlcMhvEGjb9mgEvp8KoWt6h9+KgixNwtAShweQcVEeR8lJ37oO/Lhwjn
oj4BifiWhgmnLdYu1xMvC3G4qWNdql1ApLoKODuqfQn5yq7hWVVghYFFn/AydSXnZF3zSxbFnQ2E
rAFz+qcoQQpI8pJMuA21g6XqhzRtnLBYWWRfVjFRRx2L96C8PDSXQIoszHu++SAXqzIzYHtn0i00
kcqKXl35+9rhEtfMltFWHgEIhFSZES5e/eIeVlaFkoMfEwgXGvTZPkqWCYxhF1dczP08zI1x5hOX
VtbMKljHChsVZofiffi0SN5rn8IRniOJZxXRpceVSDg6b1jIr8705vNaJC6QoPdaFSCAW99b8NlD
UOUZIeC7BugImSR92wHitGoTHE+JwUWeArhfvlPrNAqfZCowdGSVQxQxiyNo+IjqCAU0cA1tgZqA
2lCxIRizjeQH2DDxnPeEY2OuHUgLDxokNlja+A1BidhA8pAkZwBpIE2+8QT3bmHj5kaN9BEfb2Em
froC7R2+FkftXFM6xZ9gCGVBMm1ULSDmMIRYtsTCUE1iNIjfSyxbkg7oEo1xs35cufFXktdYtufO
kdEUTocuBBEjuDVJ21wwBAQZZHFpg/ABmImPAyjeBE/OTJ7H5sDVJxWskkSwGioAebcRO0qv4CH1
3BMn/josFB0kp/AaEdehPMr+UX5Ek1fRxTtmftgkpBYPvHm1aKvRmiBq7nnmmjnSyTIM+waeKnu1
mHlQ4VLFxjQmbNNw/EaXCId8sCAyBK0d9arElQhCSnatR5gpv0Jcfc/0uzXxgvkrariaHZaKGq9s
TXy6iJP1ifbSfWaPeMxurSuqvDTW7kGnwa/pgZocE8/hVaMSz6trgkqB55UOszkgiNaGxIWd6y8y
rKDAWVIQJ6f9krmtNCMg1UG0Hh2/Rod5WjuTJ82La9mfbxM4/XhPuDrgX0VO6vfjq+zeJp+2Qzk5
AnXXukBAaq5ii7BrhOcTmMUcyAkczZcR9aOjZGY/fLWo/3t7IDya7eP97czYQgfEe+GhSd4Dd61c
vvZv5aUS2Z763e23HlUjIMDam/1OyMIgP4RibsPGR9jkM+6Cn9Jd7rFcD2zdC9VNLrTARwpfnfyO
CvgCS1n6/6ZJc8N6rTbD45UMqdjEX1BHhn5Y2c0CClRqhO/XNIkoK/MeHuueaxEB2S+BrrakUY1i
pkJbFm1Un4lekp/7jMrcwgBZ4r7nsJBwCD2rY71Ld3btzijifJrmh1momuDTrOdW0ojFULDv0VKT
qs9e1r1TzZuv2issDw8FxdGAftRVq0DbGufB/kS8pdtu1fjAEoAiL2hhxtnA8xMM1jpKOH91id7+
NhQVdzpmwRUu+phx5uBDsmNIFUFHGgVNqfoMc0XbuWv3oeboGsOeNjI1upmV6T2Vo1ljgeC2o1II
NaFY2YtLDc54nw3qlu9Z2cADXvsbJ45JRu8M1WmDGBUFtyYqvX5Nn1oafFaW7Q+L7HjEGN/9rpsI
9lmG1TgGHL6YYRRDmObaIlKWgvr8q4kAiGffydGR+TbH7df86aU4zDz1c6Z/bX71ABAjyfKJzzuR
2FDODjTdrAbRWmPpq/vjL1ZSe087V2xShXkrlXl7rTDox+5Z+rjdLDTx8kncG8803Wefv7kKim06
HqPQsPUrFXKrE5Vl1mlJoYbQzYyx2SUFC3TwrG1lkG6KXKl13I8xFUvcvwEf5j8YCuK8KZVzON7N
eYs1+XE5pATayMS8PNo9y5STJLqTVxufeTOyyC5WvlM4hTCGjXtJvKzzk8B7PNdtlLDcJ2TFf7gm
a5tj3Uw7mUSWB/JvJuoFwF7pRBoudXM1taagL1ib6mTKAGKxhcidHui0Qla/g0QgwG4BxLwxX9Si
3lE1s8ecuPD3RGiXTHzAY9UsyikAkpb+r6gaVu423nBAZCpoy0s0UEh7f86mMCJ8vLXcOrrOiSoZ
GhvpJAi/YaA+UYZeOHLD/Ry7KCmXPuod14zAqdJevGOlpA5TsyvwKGUp/gk+4kIrffVw6WiTs6A9
v2xzWaGbEpl4zisGcuwGOaUYq/7/tUJN59sch8AtymS1zv4yGusGXLry1xPnEneOknHAHVpZx3rD
CpOZate/uNEcwIwoLAfNs3EU9LGXdVtxTNiUFA+P0u6ALcWWS2aQN9WZE5HPATUDzh8hb1z0le81
5pPiga1p/4l0HuRn2IA//n2G1s9hxMc8xNzahMVGOa7+0IukENdHPffZeZ+DmQNsFG5F1cZX2SMq
ZyOV+tmNd06MsZj6Ny+zPgSUgyc4WKXmUvj+iiH3/S3ddr41iJHZzy9Lnsg1IFf1iswxyS9sqOtK
FDh6mApxCUTqbwr/upJ+mNJh8mXdLGaBfjaIJ634vw2cNn1M85FdeUj7fQSyRSjNRr8gUri6cdUz
mPibXaYL8Wxym0L+gtfKrkFW5j4/vlfVsDBJ/86AwlelRlqaFGd5H6qD5MuQqG3xH0oDedAMDATc
pRMGhQHvDA/evbY9zOG1unZwmzSLrAFJYEmOS++iXmX88MVqUTNyrP8E/rcdtLVJsuYTD6SEOXeM
je8xlrLqXModDfRz7K7HvIWLUYj1Ypvvo3B2gZSyX3LnTAOHP4CaPX4etwtji0kJoNZXNZfRWeks
Lj5ReMZtCcfsAGvfRf0RJAWNnR7XWJ21fBZbdNLf7kdeIYVWX06cJHr2qKd3PtGVTgIwuKz8CskR
HidK/B2M7sX9I6mCXdB+gh7P4b5lFAapck2e7pZb0ysxYE8tftEwSGYLJm0n0g3KGR23JFPemIEj
BWBgR2uyycoBrqIVpBLN8Re2vIfQ+C04ga2iF0dodkVRKZJJzroOWddSosJwfc/3tlql+ukfaOTi
OInVzAFfRM3M/ri9nnLEQZ/usgFr7gDV3gwMkRA+G3eFPpnHwWQF1bMoAwFIBu0hKkfwq+OmoyiB
uI4deismL6gea7msqqKFgKY0kO2YwhuaUz5HL5lw1vsdC7qZaDBhmObqEaKE6X3TbJ7ubb9EAaiY
QIYr19/DDrnTgOtJtwEmb+NlPpiP3Pv8aLPo/4LYsaBXl9ZXDgkC1uwZmpRKY4oNim/+E2Yyojtx
sPFAYPQHzS39WuiOzvwuXrOrYX+ElYdUWwHHoVZ/UZgPOaQDLRBYs8h7NOdjggIlp1f63mab40Ku
PamoRogb36mPQ+dzUjWrgHH9N3yY71d/UckmwTmJJK5JIrkMEy8CcCLbCSsw7arEKu/iKlPyV8aU
cqReOLjwnUrhrKOrvd1TXBMNnXvBFQ0SnhXPwo8Ix0/3pVguRC0l+POb4ejL6wyFp5Ydu5T24fOq
pSPAx5UmaKu9Lk3m6kaEIHVmVeu+X7gJTBqhenoxEnY4Hv07wCxFdW/XsUo7w0vz7zaAOeNo85xr
LRPL6zAhA+QdjANkMa3rnM8+QOLneT7oHoFYvvsMh1Y6RVOJqD3s5TVYjUxffp/kxPZhobqGhKvD
d0q2UzjLb875F0yHpNotOJHtYt3Kuzn7djYs3lPpdEYgHJ1+CsX5VSMUtZGCoNnWAueSKL/hwrT7
gqCcjChHBd0Smn4AnHvDLe6UduSoomFugLMfKMWy8CidTFdUo+epkOT6JOCbUmT7ryQe+GXgSbma
232DL9y6TCkKAW2iWVcvT6p14m2k5VdOMEoMQDbmwr6zDf8rIYYOqpdhVY8qCg4AYtG3V1Grj4cX
GKUXu4LMwFgvzJKw0I4HjdtDDQLKg26wpNOHFctKwN8gdNI9cQ3WmDmyXBMeMy54U092zQ887q7a
D6ZSKj6ADbL5X1XWsT6TxyN2hfOxJBQ2LJS2QqypKCig2YseVQfqOvYYL+f+yUI4CNThHaq6cVGf
dU1mqOUM8p6o+BwXEi/K5rfNrnytHT+qi5HdCGcVGFVrFNsW7qXtR/492jSppoIm03Q6Jgiq0g5u
B7B14yNhw8Xcp0QFsIOcODNCaO/W4f6T3twLgIvsJ9NwUR+So2zl/7N1bIL1S5XkOBrrt/Guu3ab
1qbClQan9xQeSjGclEn+xRSQTRUXJF9OwBuv8GWUcZyt6Ovz2AwYYTz8WwoTaxMUpb3JB0e46HBy
8iCTKE3Lv7cPQRy/OE5r38k8pTW39flt7czHC5ny8+BEroOhDfoq4VuJpRYFlOxudVf1+jm4efft
nZxkE+jB6wUoVjFpav/h82c4o83G4ofrEiknFaX+7botiWufqjYG17jH2VIOnP/49ZWF8sbd7u47
ZKSAXyWfLYDZVeIKsqryFzgCguhw6CV/pusWVQnRsyqDTBlY0U94aKxFImcGgJA8k/C0X0oK0w8o
iXAUvGvQOhbGtr0v5zbuPEAznWDpM6UvqeCDjEtM0ND35Z+O95jwNc3A2m2mIhB4R54ltV9MQyVK
gVbTm8tWrQ0zx7GWvd5SQt8mc4E86AP9tzFPxA35QDQpRmEYSGSTQxmqvrorkQmalVKJbm7chbVa
ecicrA5KZG6nt0z8Lw4SAHQ9X0XLdrkQidaRRgd4tFsEBhPzPJJqzIVZPdwMusWmzATDX51WayoR
Fd1rPkWo8cOU7Si7VT6lOBPdM7Iqr1xNqAuHYzkAUz5wztE0RCyFFpHdfgLdsEzQLdjnNvP8dm3q
kKYL/HhP+WIMOVD+ucSNCFpPNXw9T1eS3yXQVuxWg3NNgwTMSA4jGtLGAHl3+e8LlZGpeEEHNK3V
t/EbZPfhC6X7BRb4on/1z3tJS8NCugPusUNwTABm4S9AUOcK+4PYJk6G9qvLZAWNRoltry4BxavV
Vf++UaTxtumBlKo/XZMCqUAwsCpHt568MITSEBJow/aWrd4yRxRS68XfKgVUB0zjeSbfynacadtG
PjGS0+8YRAqkz7PDgyd/jjp36L/Du3V3ZnKgk949zvhX5ZQeWRtuiw6cQwkp3AM3yQpQT8JJAgkv
ySsUeLYqEZW19pEridKaXt7I8alVZG0MlFxEEvOLhJSr/y7SV7DJ72jdvsGFk0S7DckHX3hzcjHE
Ma3Tc5X7BIsfKiWi/FL75khXHBKZhEgKJVEDjIvStJkT8Nau4/Yl8Xa8mcnCmesP16e0yPr+i1LH
3EU7ZXkwJc4MgH8TvIU95IuQA8DebPa2zHqjrHxeZpknW5s8dmZtcJveGQXefRO5zrdRkZPHu+73
UPMFfRaDG8XicDkbRtD0T0ka7kCzio4MRmVBrDF9MPYO7dxQ0c3EYPMktmE6WH2OiZFRW+w851FU
MM3WNeXrdTHpljXytmsycSl83CVhaPVMH+EVn+QK7mqmJwaSyqh2Nv4ckJLeS1Y3HeGdwPp2D2jq
Re70WZbjaSKWBVhFT9PeBhVtGCaJxK75WCumVLlyqBx0ICUtnXZ3YL7Mk2Mt5pc/GKvJdz63Gr5S
QJwt1rOuEfu4FO6K9eiZ2ovD3xxh9wVaJ0REOR1J3djdtH4BIkFD4fPZuTLKs6IFmbKN/OI1RYjV
FuhLbH5MtjnByBNY+uQZx7PHl2PVR5Euu5Ysgb/OFwVtk+MVadfq76cFEsY1NqHlfFa7Ezv4Natj
Jj07LPctxUzDEMhNTGg/rxCASpzjVeTEW8EacUMLvP9Q05KE+NtPy982i75rHNWt8u3Jg02Do1v9
Pp/oYfSO6PTwiCzxlS4MkvY4WZKtYgaD/8omr/rRkHEAwWHdWss+RPzaAuGZYiFWkUFIDX11BRho
3U7gLjf8lEMt19vjHytD/NfxSCdEzZi6lrzRcpn59KdJkRkFAHap/TMj0MRF63j/Oe0Dd5osqeYI
hOaI5U6fNjY7BndZMXcsNx62lIQL/yAGa2309yOWvhV7Mcr3wFJeyhn9e2vajiqNIw31i/cgab25
VUzER/EGovQVhIGkOctcFpEaHdu3ceniAxhqLUMqYTlMdN4gB8DnG6bYjbrWGZRwLjespYMXmfRW
W4gtM6SMCr7FAtucFZtdD6dQyVMztHuBDP5Il6tTyjjkEKrhyu1wlmIAnNigTvb0pKKW7IoKMegp
66ve1oapzgx36/VHKxkgKg2HukUpE8hjviFtvwvuuHK3LvaxtQUPPNgZAKpuPR4wUyYexLzcFZz5
kotLa3KYl6Vt0NMR69XSjQMYdXM8c+pW9R8R/DOuVkuKB/D9b9IC2O0OUcEbkhssNckKAMX9dCj0
9Uha3JPpjZT9CAZjI69yMtFH+Ghg2lHQoxXFwhX4ba0gsaZKtSORkiuiDUPMgZqoaeqGaoV72FOj
3nOMDFrtbcanMb+86S47YeP/EXwf4WxEJyWGBP2EFigyr62X22rhobQvSEb2BppHlsj3hUuZ8et3
3tGPraAAOj2/KtFsaFnL5HzzdC4nKPmYSC+ImxuSWG/2c/zwP2izrIPoH7A8yNGxtsy8U/+0KQld
X/MY95JOC0xKZ68TQpiWlx/7HTcMq6vJZelaLaY79EUi9DFWHrBCfNXBfFglRZFOKTJqq/MvCIK9
VB8WN6oFTk4EujycX276TGWHJrO3i6nzHYg7FAPZtM25Z9+21of8V+XW5/BmLdirFWMrpyvtVCKB
dHPxVFcAvNdpfmf/qlB8qTteDz6Y4spe4DdopH8X3UEjEOX8uc1f2aq8ooM27beIvO9v5nvrea6Q
ZAZtyXRcGOZWRwanEhiPzIrGWBru1p+t9+vLcU6fdEm9Zj6u9IIsiS9OWqlLq28cihcXGuX/LrMW
Mf2NbmrXc/NCUtxxjQMcD5OtYML6lCbMzW2hSh1M7lAGsCzTcIMZwvkgI0hOPRetqVBG2eC1U9Os
g6c1Bdam2+VuzrCg+pHA/6C9XBurYnxggM7ToXM+pCBxqOPHg7pEpxKu1069X51JH9TSLRG4eZgv
0NtC/Hf9ja7N7X/HS3GUmvMAuMtfc9mOIzh5pYVw1frYWs/XvNd1rivzWIYkg0zG+EFLCvexwLb1
nEV7b8i3pISl3hQpmhQr8uPLmTBbubIgHbkmQPEm6zmzABDF3NqVkok5u37HGDcLb+/gdcXEARU8
grIvEiH7gQx0UUH2I5YDorgGr3wYZGc+0Gh2r0Ect+fVs/YDnXlJFPiPfHHdchksrXCnPdosqluD
LnG7JeolQQRZ+DCtv5PspCdN89LshVI7gG7+nI9nAKHaNzxzejGQjM92gWX2G4JgMAPngFj2Ggkq
jKpC1p86wqQd04UVjLn+WhkXHpOUvaU3poPIRbtE3K2PbDylOWX4giCP5p4hmJFKpIBf+xzQkAIx
BIZRLcdQltJQSfprhnDpI0AnXq9ozPGbVYXZAdvEFHHG/iY6gSsbFEQFIzwFDloCca5HPElAenPV
MAgGJEJjjA8BLUfHi0BaOSfb+dkjxMNwsdoJKVvWVtAtxO/4h+eF+K12j/XAlhkBYtJopfgY1U9L
iUpl0YZ7c5kQ+PdKgusaskdcgraosVlF1TAtrL75VQdloLVE6Mmrez8W8qDe+ad1x+5/c9kMh2mY
hhzkS4sq7+uYdMyVoyL/slhXdMeXUxDQbdq8TLnikcFy4+3bhDgZnG603Fqj+gaKoVgw3/ZMhKdH
FxKpoxYGBPAQiVz2st1yAFISHP4oIw6YNXJiE7UbIjrTCNlIxzq6RGSjOKATncIIgWs/eTCeFU8k
RU6NsbZI3yIZ8n0F+Ix1LrBA30nzlnGiCycbHYYD+EUaJRVNKhFTyrzwwVgP17P2kQ94IScMn87m
H4uIQOl3/QnYN+DG22kct6oo8DhCF5V9jAEd57tXXLHg4PtrSa/7B2wkMaBFc3W7HJA4uF04l9el
/0bty8BsNVmlNW/I1CuOjl0XrF4sZ5Db+9RlHq7RRpKqSdtacUjHbBmEAFPNIay62EQSAzwvX9ZV
lNdJh11mb5OIdQ2WnZSZbgTkg8529aiSpsanVncorH9IoSgBqAd1xB2JAfT4YcWwmEx3+p7BnW6b
SWDl2J8SrGbUwbbibknrr0UXx1QdxNpR1y4HcKG5mpJjd7437uA1K4euejM83F0zTNoCECfI1noF
37Aav92O31vnigG4jGgKTUSov3q4gM5LPYOEN9jpb+jmdj2U1KpOZSrKfF0Chw5SJ3UCMC+A/1QU
0g3no9EiBWk9RApbssZRIqaC+X9qwoz1l9GmpZwA7CAG16j7xzUx69I7fLexoYDers3oRJ3U7jmq
1cHARpBP9trZdcGjMD20JJc6J6BKGPc13X3QrUjvCmWMOl6Djk+m/ZSON7BgnCebyfJVF0eqPCQR
l8JPpYHlIrl0SSNliFp37H+hILcKZpE5azHai/uBXNOe8/25fZSNzc5JPAkwHcYUIg8bBdE1sYrx
9DyFpKdtAtsrWbAbMVEhhBvPBpBimtSveKj8q0Z3v2ofSXg4Nv1B9kGD5C8DCDWJOjWSwuoPrX5F
rRgyYc28eUOqIQQO1yk6W/fCuGdg1iOT85Y0E4RQtrpvX3aj7M8z1pg31paWlBkX9aeEGzddKqhf
BDUi1jm8WC1W/hwBQTPFU769H2ProbfZAuUHKkUG6cuKG59bsyP0dMRTBghvLFmx8J7gw1+ikVra
AmvlE2W6HNMLTynLHlvm61Uht2MzU6hW3OmNqhsBtQTuLBagKPIU/LiK/qPs4dti7PQVRPikyXhY
XjL+4xsXjmCCv+U3YchF3IrRwx213NZuc6IqDch4uH3A9P8LB4qzjbn0RfD+cOYOwXYh1Ub/FkyP
ufgkajWQpTDGLHYhQwwD0jk04Vc+wYSfXc++izP/sTJJPZ+oIcqnDka/1rvqOT8b4in53uupt/Ro
xwbD8/ojF8ooznzqxWgiVJm3p78vwyDGWiGvujJtC/1vof/JNre2lUSZdGEO4woprBgb71kcqY1o
AhArjlKTzNDGM+RF63LpdxhQAMeRLpMJtqVKraeviC+35NmZGUZfvCpO9bhAa3N0PmYTo0bDOdDv
XDYd1MwAzibuDqLjqHvaiRTKgnGlzW5u/7Qhzd6pKkpSdws21g/qVXFpZSyDiwLsTF6MQ5K8vwQb
bLL0WUtNwaLxW9atkA31qiFmlgMn2WiPGB54FJqnCxZ62KQdYEhd8YRcl2c3/89dBJ1QGZpAVqET
zq2v4BJLurHJzNe5Pj4RL7L8jmoyVPZqHhRqkJaN8Kcz6HsKfiXEoh7a27H4PBWl25I7eTfxx6uR
TEF9VEfsuS9lxauCBKzVvdmgNEBVZ3xZ9BiPWB5CmnjlePTuQ5z3IQZA/xdIA9G7YDkyAs4r1gbb
3ItYe+BnrI4vbZads86ZEJeHC/3k+38UhkI7tsBGXq++Kab5JSCw5uIlSa0TYDUUTkqOOwkdL79Q
Rpzm7OG/7hRgE/KVdY3Gzw1c+RxAtGG8px5C+gi+Kj8wqdDXhrA5NBMn7ntTRLngwHzYCfqKY5f5
CpyoYF8p0aPXDlXlfcEfgs+VsXYiR0T6tBtv6VJiHEN0XjFBTes6lwYhKW0DOzX02McFy5Tid3rv
zz/BRx4ieLUY/HvHOtsIZ1GFIRRVRM+rIGFFPDxRlAM6597JOwcYtEp9XUrV3l9RAZ9tB3j0lyRO
EBXMxDFlDlf+1ta45PyfzzVVLCApwXlp0j1p9HSwdbIa31eXNQd+V6kEDbgIRCs2Ds0HAZBCjkhp
rc4ps/E4afWPVaKbszJt/EID8/2AAOkAYnrH1oHg7XGzGAJpHhtFyemnbVKmMsjHImvLP+UVeRxN
mxP2lzWHPgaGkcvY1W1WFsNCoC2CS7kSCgzMAaonyVyjk/FC2tlm7dVsJN3DkKcoWr5nSab7Rd4n
c9z5alQ8PNYqWrDXxKLVHE7zRgJyDAEAhHC+KgboNKjjUy6ElviuXyZeVKzHpQoBxXgVtfmwRRII
Ld9fGJsu3KWOkErTBJUNPaho1hW6wgDdhq7Qb8KNfXh2IT3qHvp8J4SZs+eJ4hvuY2V6M89YPRVQ
UOlCY0NObvI2KnUs/yFh2nSEaZim3QtS/HDieczL6A+DG6XWiM0dnNnCCmZzfRpSgYBLOj7F1Znb
RaLG0ThGtNfUJDDLjPpGeG+f6ZEj2fx2qAHJ2KlEBDMZOVA+4jocRyp1q+wHtSAwN964d7I61dZV
keltasEAPnLpC3kiU9j69zjEzD8dBKUvI57lYliV5+AWvNmYl+BJHkiR7dpe8/7wmghZV3Scq0Kf
6B0bK9BxDHJV0uj+/NHrACkDddJkMldfDFTCCEmJSxru6cwgqI//Zs+iDJHtV+kjEYi61S55GiTZ
mKth6Kumeq8f0kGMo5hqomfaH4mbchB8vEuQAf5GwSce35y0TUgCHoczVrXfnqx/0dq9feYLs6gJ
026biDmGvs7vmYb5xgbb+0/eKB68pjQtGWQ8HxL8imZ71K3/cZnCeR8qwWekK+4qkt8vU84myjVd
07tdnPOS9TzfKGRRRTxnQwFb/vTcNBYxD2bRpY/cc8dWht2Mpub7TLR/vVWt7EOFPHKJh4NfMggw
Q3Ck9+uTnd2Kix0e0BqMuYqGxWI+iCpYj/2gc1ZEznSXcrQofsnJeuzaV0M9P0GRK+JcrxRrXIOX
nd55ff6MCa9wQ2nZzPYH+8YWCjG4BiTxCWkRqnWYVMz8fKCYRLBgnOjDJMV1dkfuHYX1/7xrcs/c
Aq8baheSz7S5M46MzIz5nce4QB2B5iyXIPbK7KTCTzZ0uj6pickAux7kEwWfrDLbVKsQA2FpFj8O
Z59yv30xQDWVbuTq26XcZZTHGlXtYLGe4r57qK/Ms+tzMy48fo9WIZUXZgPs7PZRSGZNfuA7DMYb
cjgVrn1/qWy94tTTurLE+oXGUpC5V+FoncNZ2pnOVyTkfpFrnM4uo34enxynAQto+uzdxqym7QLr
kdCkFQ9FlooqFiNshx4go3sN7AeWVFdo8klChU+WSDLpqsONL0Bpt+zsfWzvNFq0yz9LA2XTuu/A
pLQBYQzzVdkn4XQlSEjS8meJnLxmf44L/aVjeK0RG/iqhOgBGHPPXEj5q2NKc28/XM2IWTuuI81q
Hb5esqFikBvdBdJ0fAdiHARu6Px7MHbZk3IgQndULaYBsKPLY56Kpz3IjT3P5uFuFfxRicPd/sSl
X7aqLPcayWOEMdd9b1/6zaXUtRhCu5b6KOXNQLGTz5HwgkMczCnUwkjTSXlX0iQmFqoQjYMHU8Us
Y53RfUtcECL+0E+AVk8fQDNOSEHHjRkvVEaZFwgykqo/GufprfZiH1dG7GDhywVQwzQh1YnVvoZe
GEpbCensSrwJ08ASG7iGLyBYWemt7Q8XlRnLey0P1ZHIFfTKBEyVHz5oEoveVbQziYFkaSDzFOUy
+aYqlQV925QERm9lFeqCxqTEojqlZ34/rgqptPLHr7m9lVJi6foFLgpuQeiiSR6NpKUODW6dp0Jg
t7FPhqUGnz30KHGdLuODJbmGjMrEOxuz6ybQskgfpDZ2WgfcFWKJW+3whSXDlsnJKxbXhduqYpDE
JIvuhVV9nfPpqTydBcENS5u92MsuFMloTPxB834/MxNIvevcJncLbT9HT+CH+LR5sl2tfMrp3OGB
n9wGEhPG19wUPd417nMP50cf7DJcxXSvFUNWvYvXuK9D2oUAp4Mw3Cq/rYBVRrLdNFWUd4E4qmat
i2n8+tKAyaY8iDgSZfTBukBVt5d0oq2gNgMw/Zny/LLXQRw86MwVg+hkfg4V4iKn4dLFFSR+7rWc
Unq9T+zahD+2C2C+RcDGtmw0f2/u8dG+oNOm8NQysIOhowzZfyG2SKJUg5b0d6JcuWs2RMImqNpU
76W4XVPUKNQSi8rqDQCuWYurQcQeSeY1E/iqakbgU5fshrA6PA1YGLpvfBkIQPMyLwi0GS0eYae4
7dMSO6ScPKkIvsSuDW/2NiT8c5u4kM3AoeFDnVplS/SSQVj1Q4W09mdOdduCSfhEyU3hac7geE4F
YRpFUko7TiNHb3OUD7hsMeHeA96gDwuYhr120Bh7X8+HM15Oametl2Yl+CjMQeCi1/StZJbGaymH
JvKzP0bAbUcYbV0YQfXxpOmD7NXHI6qjIBjforLbyjUfAVmQjEo/uMLnafjMLU1Pjizr0NqEXGAV
20DmW2TSKiDrWtKdg2fGxYAF5BYUaYspi1YklgA04pTGir/HZb7wAI/F+82NLg7cCQ98XwO8Jd8m
Y93E/mczELMmgIXKJ+knhHx5PS125vpktjZpmJ1CybV6m+GTpqfETHRbtHby2Ho0iSaov9c4lYvF
63v/g0Wk/eYKAF4u5YziPrf2ABydZXqM/mMyFIBhM1wKKfEkTW6bwfPXXqaiac6Gxmz/W0Ez4AK0
5yldds2x0qYBlxLl7NHWDT3HhQtMxw0p0rriEILQIgNHkbcruL/6GXICD6XzUqjBj0BL/NlpSrtE
UXsZ0/+O+gdqsg1kzTQY1ONTCtaQgDBoyrht9e2LjjfqvG4mReIH4bhtMpBANGjPjSc9Jh7h9tCS
okY7H58e61TbDyx79DoGHFPA9cRJItpacZvX1NMKs3MfK/Sjy+914jhoHdsSG11tG/15NUErEKK4
TrJ0YL41HIUW7rYTOw/5+LTnGxnts34dJPoKFuM8DfBbQi6lTsa2OS9Z8ICYglgwH3LVIj6L93SW
fulLdK3R0t+eJu6XJoXyhO+7jFCHnpUlvDlegtt3K2ebPint2zfLf1tvrNOLa7bkDkKHSmOefTtw
UPoz3jFGZIV/V/rUhCLy9H6zn1xwZlXaMA2EDs7WHzUCYkZZDPSZR07c9uvXbvK0/cUvSUzj3YtZ
QSbwFCoB+/2kvceFRbtP3c2gjN+am3TrAGCdHHvNM6bE84nEefd2bZ047nSDmw5RfpAZXrYD1vgf
ZkLZp1hvCx7B2qozBuoyYxUJRDxIfAvn3jtRPpus5qTHl4pJgqdHH1QEx4zLI6e5k8mETj9OgrVE
vlOZpwFvqZIY8vqC7PnQsJP+2sFcdrxVGlJ47kRZdJkcvCAlJbji1NaXMEdqR9p1q+gI29qGRMK5
lm9Jb93pcb+wiAN/5A58rOqqNSiXB582WE8WvNUIYOkZw+oe5iGhNxUqc2ZoKY2SWa+pgJ4m3iNN
CuIYUzxtkFnytbYUDz2StBiAcdoYKPmH5K3s265mTnPdkeeM4IgjStpwa9KJxOFjexpzwu17EZXo
i0xYctijbFhq3Us9HQrUHLU4fIjvjA/DZYn9wBdfArpmuiaQYOqR6s1eos/FoXMri5xuJWEmsJro
o76FxYTm3ilHCon39Z78npECRUOUOY6xCXA2Tv060SWQHlka7mFZjxSLzAoe6a/aJubg0t+nAnnm
2dElczqraB2VxBIcOoNwvd6v8yCqx4lXLtHER/aaYpoA4UyeIDykXi6ujDVTbf4zcbD7rDs7hbMU
r6RMVHukkubB0uawUsYGOh9btelHtodgg/fADjf77YRRLKMbshuVE7XPj59PhfZxJUG15AGdzKTo
AOSW590phTwM41QV9dVf/uas1+fIbxCjPJZ76mccOlKPAZDUauuAoAmJnEW8g9eHUaili7Y8wQvt
z7E1HkxhK1vsC3jjYXMRahGSojuY+sm1P4ADLzPXVZFWk0/Bvy4ab3mFsCYcgJiEsAEvLwQoPF2g
Gihuc4YuRMXvjcQ5H5cYBqQ/OrApPetBS+5L/u4qvoIoeRtlmt7od+K0sZoOIMhcZwWbGwwOelG4
/tsDhSLShA5kEhletfZaeDfgFCz1woExZ++nmbnovfVFr+CBVQgB/4RTrK42gSzWcDkkU8Y4rHHY
sUPpHXz9B9bi/fiNOn2mLMhuOBXnU3JwOp646xmHR0XWgkM3p7sY8jP2nBQjUUown7TkhUpibEVr
kZZ2gP6Pjhi6ixWmIJvwpBsaiI6eOCM9jGkguYEbxz6a2ZAx4blRjLl8PN02qb+5CMhdbX6lrQfk
hYiYGWi2To56Nria+ZtxvP7H+kLyemLq9EiHDC+ICLJ7qixvqUxqV0HIOYPODuR7xO7W9jkKIABn
2MsHebhV3v9XFZk73vpG8RFwlEfFtk/C6fCNsuF3fwxUAcgx9AApKftluEXetiyRPiJoUD8OUJll
lpO/VdWL043Jf06nStfmJwhlttLF2QVfidouI6y/Wn2hHBEhhaMqZQpSyudoVJ975sE0qVx8Bbsu
IsG42fV1qs9O/g+dFezvUJj3X838ZceWo+5hMA0RZn0GOh6CDiFpMEtkahhAqJtBVoic5tBjU499
kA3qF13IGyOfBVX4CaEuBGlHoxcTRt9CiOkdgapozcDDCPCCSQl337WgvvnmktXZNdKtMWBeHFEr
Mjs7BcoSGQXQ7OULiXFNe2peVBi4XPRvpZ1XOGdKWhCHI1kI1JcLt8TmzYBEgH9SJg/P1EIL4AFP
7GAwaO8FuHAYrsmykkD3c2Xy1n7cLgwUW/y8l4l0svwA/L8BUwCe5RnY/+fjvZBABDP1xm1G/s/F
zmmhPSyKDQhf1y3p+kCaWLyozSZ3Nztwxog1kcYquKKB6ZqK2ECoIu1TfrCraRZpfHcWNkL+0pgK
BkPV3ee6+/eeWkkmY/hj3zkN3GgPIzp1E3LThOyPc0sdR1RYxgo3H9NauZOVFWAF4b10YZqa/ATQ
fj7OOfbKPdKvv9iNdh0RRAfK92qo1d1nrAOY6Vb3HHS0QKYYZ+1oN/jriWZzPkWzGVyAnA9DJYvC
OhxxKYBHNwp6PLEpIKCIdjFj5PQbIbvKrupIUmB7XBo10GFU3YBQE2nla69kLwT/YFkR9rDe5BTM
piA9pR+AxKAgyefzMe1md8jLNod0SPLojQQN5Mr9018oUf6BK1dT3jauvgZkNNjpcFveyKnmeLU6
Zfc9SaWsSuCGy5bOmspFRvznf9SfUnvN0jj1l0BfBKTGuQoyjQ4JlJ3OCv7FS9F/ktfgOcjoM1Un
cGXVIuGWTZHVZhjhmsgoYQyRuljCO8Ukqw8O0l3UFv6LmIrIqWSdyO/X2XKYbJxIiXVGFYMjn9ET
mWRZVcP1MzqcVo2QfmcxMUPGMRvvLwoz0n2pqzewN5yNqrwzjOdcyXquOz7qyIhxwojW3XKgSOmh
sbMgVM6EJR2q6L4Hw3hNVvNL5HmqrS9K+lSimA4viZBmpuW/K4lWSC5ypHEAHiX0Lf2jAy6xZ3+s
V1C9M+xmT2NbG5XSBPgJs8TYT1VeI/uwFmj7HXe4PrULAwvI8EBpR0xb+vL9UZpD2zt+0U2hkg/L
c4yN0I8cGQgn64tdB/0WxP38MD3/7K/Mi7pnnKMDcQUbn5mBU+MKc4YI4bc4pNu+u5Ap2TxDI1V8
RtbDCHfgHYw7RtU1d5h7sz2TQUplUGy02VKyaK7BASClQWihB5jM+NXnOuT5SfzYXEDX0Rxmq4Hc
Vfk7Bz7oPkIBl5bjXwURPiKWi6y3YG32SZq8gNx3Bu0i3Ma/Dpu7qWcnn5h+TeeQuL8RijXPNQGL
hD0ZPwAcKdSIcy8mvowiwqNKFq+MNWlc0CFdZS90juL8jjdCqRzMaxKSWwTaOWyMAmv/OEPRDrd8
M0I6m+7KWPbSrtg8W7gSeDb9gQV2JtHNDwLTQT9Z4WrBDWTisKBFKAiKOVRIRLg0Sp4ECTQdV/it
V+yTRcCSTuHqqnYYrsvPWR9GoiQ7hrcwqfqvZCyuzjm39356CPDunCnfz2t/TkH3VOxf3RwbLd4V
GDIw4J7p3br8MxBmwYbT283OlUlQLuF8gzGjiKiC64muG1A+WF/hvKzQ8NS6dZUgvtrMu/NWbu8S
5ZyBHfCRpshxzR1FwEUUxVCDPPOgq+Bu5bEdCbGxznn6RNbhocasrN7K1fg2jb/yhz1OAtimnGe4
8WizdaKgn/JVdtK98IpEI8gCaBw+1GIEpg9I7QyAs5ARLlvO0qBykqdpcF4YR/Xlkfj/PXc1apvn
YFTAOFreNxtOyJEfi+1iIkChgAhJvgwOzS6Zkh4A5uIIhfyOxdu6bRmgiGVmOKxAQDjBjzuzbfQA
6n40SonK9vxoNt04jptnYaUJvLoDW8iy+Lk2mq2IWsZdK5fXKQCUyHxhn93g1DjoaiE7EaNJTBjI
jIGXYh4R5GdVe/AlogQMZYxbAZkM3EjQqGt1bpnEBCkpLr7Tp1wA0kOg2Oux5gNVr/VOol5rjfaq
s7aOQx6JFsieBALaJwSouqPAWtfNdcVBB2s+gXaEqfo9OhPgdIREKODaKP1YsuHE00Fe0zpCJYGJ
RibmPcv+2tymyIh/u7quXqrXkivwRSfetHK1LikUy9PUMb7nhvosvSeXLT4epN72OsVp9cZ3l6oN
W2N6QRYx9PXixEkTKyQ1IB1YskcQbTxu60fz/kqhmaH1+nFLSGHXHQ+gmLVxPZzmLrtuJ+Im9QG+
SZvP3/4Y478z3zy5Fw+QzSUHR0OrImpPB3CmUXO2qjNmuYIFnbEus4Epop6k28gwKqxbn0vCSN4H
VR/wRipgzt88XLVPWlEig4Ne4uxSbLWwELSXgL+yMGkiH82K5cJLx3li1Zvymken/KbmQc46KKWa
YNG2NXpo6uVE+eTZIAvTl9cjtMy6P6CV1ZdfHSUc3OQpP3GCeaYRHhWpaDQFl9kr+tRWICwAaped
3RYISFLBgf0RkDHQHvdhBLlLXCEdw5l8vjcvY5/GeO/GmLI91T3gGlZZNIrdeHqSjx9qeYkLeiXl
19iAcVwvwKUBUMtYhxIFvw+tvx2PYcRN+Y7l0/BH7k+OW4RBTdvWWMYYF3u0yw/7yFf2JcHAe1Dq
q8b3WGqLOULr+AxFakEXCphcH2lUJeUePifDW0hXIG1afhNozJ0dvxMyR2BCgfqfmFTWivZBuYT0
+C8yNFYmwfsAMj9nRO/29AGWTSC5T0obERvRu21QKw35VHvccb4lbzzgCNU0bbCYdrLLPN5nL+fa
6bEMTF1v1lCItk+62Ew8HrW8vSS+qDe2XKNseE4Nk3IhkaXpgK2+SSpMp/4U0yVtf7oOKA0KX2zC
/fST2BoEfFL+OZHbcUh6DfZsxfZX81sdHWUgVWeSq2EYywbjrmB5vk7ihVs4Z2tMQ4mgncXxxJ2c
QKFSB0yxptKWJLoppPv6bwLrb4Iy/+qqww5yI+oW+7JpXWpW9JncVxU/Wz73gnc0iwZ/V/s60Fby
56aC2fkHtyEvLuQ3kTYyh1rBkOSJvS9dZ/QJPQcb+qOwHLQqSDe1Cr9YL4J9MF8EErEQD2EKCKHU
7ttJz8R6vOTQgKx/1I7Jo8BV2Kas73wUFDz6IOSvKQ8GW7k8XSN9j5GjFmjy6KtUmYMgplplAHHA
ncyeOeXxZwciu7LpfkVnUNRdYueXSizSH8y2q6ozlhu8G/ky+doP25n7uVrmFbG7aiIbdF84kEfO
toiWmfGKlbYm8tyNZnecXHjGhojU46IFyfKcXFEOxDstuCWL4HZPjHxvkKuNyjkj2EU3wCxm+eBp
Pr+mBRYFYXWeeFZuc6Y1+8UvEFDHN2oFb6YDgyUSVDmHClFLMzT9OR34Fi8gVM23cEed/EGLRGVF
371qD7Sc/G6p4jQmI98WojCokMjuhlXqjUzCivIpz0mpXiKt1eg43xgmGHIAcYULzhyRXnJs2/uS
Opy6kt/vGX5+DoWDcuE2cgmSYJbamriZLFZAX0hbmUnF8O9QT6fOYpup5uwuykOxXCAM6WS+XQIY
yOWfJqNcyPZNWEuciZXQ5wqEoYwqfk7CNv+w1kIr23bs50oWEL65MsML9qxG9uRTD8GD1PuxZdt4
kOWIW1oGY71HXb5EsCgPa8yyCo4t6TSb6Z7PWUNIWmHNFC+GCnUY0jSrTuUYXDN96YGUZhc6HgYk
0lbU1EMhJtQci4xim9CZbnn2VywVax/z/4DbfLRSR+qBx9CbJU6frVI2eEZ+kucfwJ08xcQ5ARMu
C+NvIJHRHHy98jfzpsxsP1XCsQPOOY5UFoNYx3y1TvmfgjS9tSxVmD3t7rkAPOtP1C5cbIJYBao2
Y4WjPUz8K6AjS8PIJoEcHY2dzQmfnGOmgXeCPx4RmIbFS+oHT25/rc0pgz2ozJOsEB+Ug4n9UYmM
r2Fy5w4rmmIPXPCcJhoGbPl/N8trF61u25if0vjwtBSdkXoSMVqT9Ltdpkb5mwCvfVOHIPRuGMd8
iFdmtfqSAciVF7xKp8dQkjWqfm6Q5vkCBH4me2L7shL+tf7MGOriTpzPEvY+js85vT9bTFGMIY5v
3RRco1GpXHwYKOEmd6KJAeMmM8yfUcof0d5Qd2lOQ61kvYwt2qupnr4EkiSQsSzgHJ3HkCWvJ3Q/
PthOghuz9hfsXJ2yEM3JCQfgsgjGTlVZRwMvXP/VCkoX6/6c9gvSPX8Brx0LoFu16c+k9dfJ4fv+
aBh2CN0Uph5qDX87gK7lA1kXQwPaqY+v0TIs9mTVBjPyHDq9ll6pAUD1PBF+HsnSCHZSbmRjno0s
qinMWBvozSGW9eFgVwZi9oOxUcQbTm17vBMLIjOy99E1i8aqwX6eCGTeSCf56VSboqmPIOiPKJcP
Ay470iSkf4MZmqU7pXpdKsFUXUfBOkq6gCe3KkUOXEpXbbMXomrFRN36v6PdQrW6wN1ueJe89lLP
jOp8cqBCQc688DLzD29EJcJIzkPK9ZwoqDiA2UGvHg62mYGWIdmSmVYnrn6JU1V/NNP0eL8wecND
NRsFY4SKR2kqzTeabWaocUvNyPGFyojQUawe4frqy8fDfHe3dzDakBXZz4nL3+2ltMMw6U+vrGPz
+0XQLgNR+JplTBOUC8lMFAXghAhKHHoUfabHuA3f7QU34k+7vdnhvcdG/vJMn/1e8bh8x7TSZU61
qAkynzmPGR1XjKqys3Bir4weNF9JFJKb33awbnpCpZB9uHAaMdU+Q9p16m9JC9F/3q7Yt25tMKYj
yL2lHonS1BQqxZ06kj2GPEZcl+HN0q0S9iT8NdGVULWoDBBYKAaqo59Xo7tUtaPReS5uxTp7cfaC
8fIjypNND3Ixt8hng5iKnRM1vM/JY0uYS84cwnTXKF/f9UBRy1P8RZGBqzYVmzmr+D2/p1cKY4Ug
Yyb8ENAmi3X1uPxnOFzKybvi+ocaxVWx8oUeUDBFmT0gC7YjC0cHrESry4WEMrzPK/VuOJp6Be7x
p1NOn70AUvw9Bqrq3KQVQ/1VeJP/8AkQ96Z1dGOeNaXZwyWeiOy9jwIqJPv2E4j0VnSamPPgae9Y
BK9cdMmJH2y3ncCwjydaKBmBHGD2QVuiUNC1Kwv1uZPbxNxGn1ZVAUtGphCYMVCRAe5JKHfLjG/d
+k+AUvRblB6/IkRSuaO/ijwc4ryQwIPhGfvio/ROIGUc6tJh16pFZNcPEbKDy0CfWGqLXlIM3ozu
hVnr9j4o6AnhGobLHNBEZg3pa3A3EAeXdY0oBjeYB3bEW2Qb546ZjLxYtJJ33hIgXa+PDI4P0o1o
Frn61zeIHKBTFjGUNF1s14Smm63/DCkWXNVQuc0dtXnWvsqRlJCbu/HP1vWsKbHdIkGe7u6QIdbm
w9FVVP+jCtxjGnWDcAD6KSPL9YD6sxgSrTxJ1F/8XVCX6bxtqEUkgNFHp2AMl4c8v+wIbB3HsDJC
jvXE/11IZhsNGCx864f7uNHN3tmxl9VEEa4WFsaufftUVY2M48BjNSYBZXTktif+T6PtfMZEnchf
Akpk5pRS/hgZuLBjpfwHlOLVzlJ1B6AQ/uz+7tM6GJROBP8+o/iDkSA51AI9a48+IwsnSE8BSy9A
xBgSQXFdsNgQvukRtVuzVYZta5itis9oC0Q+omF8Q4SMkMsa2+zVGcbxHcel7hnXZcCMM/HC9f/d
QI+IDiUy+7eMQNv/EyTGk50RHAaw167skPkQwSy+X4czvUX/HXjpl+Zsl7iPKHffe3YEM43azAk3
oMjlt7tvOsuZBQJj1Wl7G5wUyZSKONtriJIUi3kHsG+ihmPDkcb1DHjWmK/49y+8YMlIL6D0ecX5
vG8ALzjQJhATeHEyH19Fxc7RRf9I4NV7SoWVviP3Px/3JO3IOpNghOIL4LcEGjgMH9nhttwLGNJj
1hdGBz7bqKR/tihUQsJQQTgTqaywsjSjJSVLzo5MoVTrwXFGtg72QMPM18gjJ1HCW7dEnFxDyBhZ
bilVhZHZofN492UHgCQhHWxOxvBQiDi1TozZD8ltsP2MuCpMCwUYQzVsVropPo9ynWBBTiNTqj7d
7iXm46kctCH5aOa9v5SWSC9jVN+vBibmpK6/sHug24japYrdSZS+WzGXmy5xFBmlJnBSQRd3gkZm
piUeIjIDY5OaqV7C3fRFOuZnG6fTQVPBJlDNc+Zxd4nwoPpCJSjoAcFHOXy+a1IznoHY4jd9vcwP
amg+tnuAmJkRgClAv6540SxHARViZ04gc+OjdIjwOuIZOFnK2WYSrCGB0B+k9pgWxmnf6yXhV/z3
t55fdVSw1vS781Z07Cz9r8jOp9BUeMVLRaiC93FuWijaR4GV/Z2qGp5itWm5Qw+zjoHivCvef9S9
f1PJjaWvo/u0O8VorZG07X6rJOvTXZ5kqMlRX/QYhnhy5+mp5nLZnuhkr4ulejyxzg02W4IfwlEG
4aghXSgcfECPL2P32s4mzWz6UvO+RqIg7rynJCMv9YXDq7KwnTZIT1bZHLVKr3bdLuKgT5WY9e8+
QyXSvn8V5B/5KmE8ZSu8xqtce1WQcX05uBdz1LT24cF0Ox+g52gN5RV5lnKJtkk3l13BN6g+btw+
/UNvarxok8zR8BwLLuOX8l/9+uSV2/emSjLy44lf2T0ftwgeGHxAik4Lf2TSaKLXHTAvE8SvRx3f
E9mCRIY6mCp91+SanjJxjGzWBiw5jn2BzF9SrVNb9GtpU+ILzITevcz09eGIONkinXyT4jeeOTKH
6KuRuJJxW7Gir7zObkYbjAPV72z++VWRloNhCWqMFjoGKTVvj1ryD7/HlUa7yvsok3usHQC/gf39
4Xwd2lTMnMu8JDO7YJeTUIaPhtVt7gkxxue8e2nh8ZdJknASkKFzoN8wRVHdAlv2s7RvjcBPsd6H
6HD4HOv2L9bmTsrTYzzzrl5kakoO3apGY8FgthXJ6juunPAJqc0SejVRUC81DqroD3UBjcspjOkr
VXbBaNT2iYo1tga+rA6eSdHPDEe3TtKZRNFK3+SgwQzd7nQ9cpz/c8MW5Ny4WY1m6gA7lLh8iBpN
1CHxVj89cAtGpjXDM8fPJuNsSh2kbpmd0yOF7UrZ6EeK/2/7cwk3FkT0tAgdCnF8pjHD+OEqfYvE
GA88vrTkEyx6ncLmzdxGEDIKZT6G7jbigTuejnJ7++QngQOPGC056tR3SYXTt6HzwLJ4wUSlVceX
AOGW15MqjwrQDSMJyQuQyQOGhJxCIG34fBOGQ3c4DuEl3qlNZPB7h4Km3I+IZasKWB72R0PsBVcD
Bi6beajznSHfUMIQ5AqT+gwp41f4IdJy78TriYDaF9HzZp4JWL62ey6u/Wh1j4jd+egHOMYgKQui
pSPWNXf80zBy00L2ClXCvfnKeXoywRJzOJ/dX+5nWBDKJRRzAhyV3wWTftruxBX1rQ+z3QEoW1BG
wCpNnIYpgqW9RhSpV2vJDedTkDI00kn01fwOg7P1ZH0m7OnPTiNUeJ22yVgIKa/UWZ/7qWnhY3s0
84BRofpACVC5coRqddQvbHiZWVFyHpFZAAKKohz3R2LD3/vFW5c2SLzg4obKn381q8O16A5XGSBF
YAekjh1PhRKOJgnQGJQ9iAHmvGkoytVNhsdJf5Y5XyCHoSf23mZt3Vi4h1IQmFybu+nyt13/x25g
lVF/LtWfXgYuOBHMQwvkgDgmyu78t8eg+2Z5EYUPnM+QSmuycj4KAJx5E8JpeThrcVZ5YCb/JY1y
PwuPkQqFn81owMP7IjdIrGkFu8aRtCY+9EiFEYCZlA4YA7LcEe5GAAcg8SV7klkjkB/JVfYeiX9O
yDK4sqOccasSUu1muQeg6PO1rzdFD+efRjgyEK8qep8ot88f/bEJHZB/B49BwpMcdnUjX/OmRJqu
J9oHc4NmCnhwt3hFvBKs78ICyE77pjxs8Tsve3/mcfJhdzqAkKGkMWeMN//DkLlQolVcAjBYVwO2
O3xOvKUCOMQwxgIOV/sJ2yBtL7CXzvBg+6wakbypyunQV1F0ePA76YI4Z7gaFy2QYAQv/JB1qbTL
4B28CxYdzXu1cMSvykosgPngcIzHXekYiqpZadPKTlIEKEAHDLRSmPuj2Fqs6QWQwRXhcCCKuvqg
95SXJvSnCeJ3ZopjW1q/yIAe2Ma+q6m1XSzTYqzp7jysIn9jEjMihaOGg9N+BTHG4sLVZLcIi3JL
TtD7WM2JS6c5qDsxMIiL5WuLz4MsCdy2JMvKidceL3RBo7RbGjna4CnBgu2K1wVsM8bmcaYhcHkX
l40XUGK8j2I6MgDxCiVbi+RZECBLyh62820sgPvtAe/nLVqs1GUqUPHsKqfjAg598BeY+7zeQgVX
JsP2oqxCsmxM8oSQrXXLCOUslpMng0UXv+o41wKoIwFohg0Gc8PMoX7fVB2MF7QmeOyxNrlo9/IA
HjPaqpGPja2O+jasWm9fLnEnplR4/3BLz7CVjUC/qrrlM9dmyGxGNoPOV56FttWrYfs6cW/rrsJj
2/V3RUD6hc0ih1ZfkgLkL6g5MICAJOt7mOX7VKTfsEafR5M2RPyDASjq/jvP3NuCdbtpnp8Fnwb3
CnhTNwF6svENZGNjhqclTcMBwK5dmCPlOPJwiyWCkfhNKPR/7ttwYwvLYxxuA6H3eUV22WbLsxrc
5Ck9vFmpb7p1Udue1/XVixHHJaVfBj2CeVR+77i87ZKkWiQGTYECv6+SNW6Ne06dBDyxewdvjSpK
R2wR+4i7Dghv9Kf1rM5L4Ewep5IOA1lmmFha7aO4sX9tUiFwmkHjDwMPAv7hRkzLYIRIEHb5snUv
c49/TLbQEOFO9Z/udA5Ta3EncFUvXHwLcT1uqPtnwCNyUIljZ2qi59mB7N/CZc57ecgnEyxYM9fm
PApbnKTnG5rL+45qzMVfKDBS6LWlu2aGH2grNFsWY2hybeZTIuKHuSYF4MfNDccCsNvU04Ck6hR3
PgMIcDLrdmJ/P5uNpHc3f+j47Oyh1AiGrf+Aw90YqVnEpk7+YjULNSVPqXE+7oioPJ4lXWdnCzQN
CN5u8IcTLLMRGTHyE1ecSrJK3HsC1OcSfyLugYWTXY31O+H+RAcXKoUWhNGIPoqrphBWSTJ1bXPU
Bgc6CiKJVI/B7K1Mifa/qhCL2M3uietYTOjMjfJ14e+KhdGYqWvuS9oHVG+Vwpy5q5WGxg2VIbFD
q+7dN8bbf3gkr/5Wek3JUK7jYsoyhEkq1ud6peMbKYewRMEOaLqik43XTS5UOKBZyCW6cYOeYGf5
pSkg9pGRxts1XeEKiaGZ3lzXx/bQ2OVzI/GwQI1dWXZcZMaQ88YyyUw/TJKjWiX3Hput4GGrZLLa
AzUM2mayvg59vvRk3c4Od1NKjDmMqKFDv395Fz50juE0OG9ro3Zbg+OBbB4apDAWo1Q5hAMANiel
occ6A1toOyCIpvBdusscmyy8pTunncLq2EQZLpkgEvA6gCsFVw4x1CndaCfPzyHSTnPQB7l+P1oP
pZqGOocvbhHCYmR6CnC+v0fCj9FUj25euKj/BPnQfytU0vg4+62BrLIdwTqGMjJwiu0T9e2lczwy
IzzIVSR7OSHLSIHJVOKpHe2eoMCrNuu0KmcCdiFiKa5MwtBkMvHfSagYdbcgJW3a1Ex7VMvQ/zHP
Jww2cpqjO9BxJQqUfq+2rVK/SHVUoqFUdkthKQwAwgzeu08GLlCWiArG7pLdUqcBhSI/2g/cBdSL
/7Aq+L9lW/j8rKUz5d9rxHTkRRfeCWfFdWJIbnzbkV7EvP88WfKDnnTws42aGq/TVsc/t4NFSR9J
blkgIPtoGcYVJJnhRWBRuFbx1J9WhHf9UsQIPMP7ob6Ct9471UPXzOS6Dr4qM4khvPYtA17uQ7DC
wpmJayx36m8kLdz+0MTELPj722QelLxY4TJPBp0BV6tRoTH3frvjTefy3G4/+HYL/Z25JmKgVnVf
M7HTwMoMUtiogUYa0hpXPv3facjbEQL0F6XzTRDpUqKSVhYtZOtSclLMdGMscmkA3fyH2Sy0YOCK
VSSGUoTs3FqQGsS+NuPmxwf0pjbdDVwnzv8xoMgWVx820HpctRhzlqu2Tsf/Whn1LW3A+oeCAbri
qfOUmNmmNRU46Z/tYszkCG9a+8J2lMXnposwZJjDSj0GMJw8cjjym/IBzBjFEITBo/3zYReubQcN
MUSGqklZnRovs79En8eUOQk1CYCKoZGjPiYr3fvzZ0inGLwXPpI9bm921S/BbdTLAUMTgCi2cM5V
lQybfpaQdi0tJkSuDeMx9Y3LnoTQaaZCLRPNEGQ2VqKJ2ZTAXSimXHNTbJG44M+MqMhBrgCcLf28
ehtFBOasXDE3F0fRZJUT7GSBfrFSjPqgOUFR3WwElaiUhNQNSBa0eRolYoI7958TzQToWtmnjuoH
ZAyLOtfkrO7YTg2DTxsPHP3d2F1LugUmNKX9mVYH/Wh4FMnjw2of/UJMu21zHbQrINH03pryFjjA
hSEI/ofPOWzwGeNB+UkhxCPoZF9tdl2s6PFd0sbZpCRu8njmtpWcUOUARCKj6qpQK9pgo5k6KpY9
sdY7KrPLKtnxBNq/+F7X6C623jlQ7QT6zgU+zuCv3o5B3arub9bg8OZwRriYZhWbURiTRD/jPFvv
VclTuYMXVRXsO9F84nNkm93BI6shtVQt5ej3nWcZ/8/f/6/1PjMLfoBhbwdutiM6hBHyj2knSZQR
/Ajq4vN9N7k301+2xiVu9CYbZvwpzEvClbPad3EkXji+0ZPksIcgpqDCEUVBKrAqtyWTOsYaW3Nz
68k6UtCS00vX831/vQ+1cvFxoU71f0R2RSLfNtDLr2ccpEQOYFpulCZsCfvA7mOuwT/9fjhnZ+gS
6LPkQ5RKYxqO6sv4ERDAsGH7L4alm9mKeiB/Wq3EfD95iR/2wKA5aMRDt0SYqny/O8296Rc09zPQ
n5BT4NzijvC8yTRM/c/Nc2IEvouMp4NHI4y3f5aGDoz+Cc1v7UqaTMZ1B5hxMOK1cfGPLoSlnQ7H
Wk+r74JASCIFWA49xWKGKO1J6VCy1UE8u552asqYV9nMvo/M+DKtQ/H4vA5Fr/DIki3QYJ7/DGdO
C5BohOGc0oRHZvUBImcS+Q1SFHL+yiJw/8qNEOhF9V5NuCUhZok9cF0qdPM24jbCTlHwpPHxapde
zGv+2kEzgKMHmsefs2IPJ09a3qBP4bseTZgdnuQBiB5rYpHme6fwIHsvutTEtdrdO5FaH4Sv8b4U
mj7SNRkxnQ3nKZ+JFpx9bqAzLqZJI9AF/3Gy5BlL/6q1AIDaPWXVXGDugijY7og1XO6JXrvs9wqQ
zvjvHvOF8Qk/McMj/7yDSWbxDhkznb2X5RhUxfseC24d3KjqNjCXhUqoWUwuNUE0qxtWIRzGr6WY
vQ3RmfTTrNh6b5UHyZ9nW+k9yQdyP1gCr+Yty0uelO7SxrUXU5U1SxLSiEANiMs0waAQvuQc8O0A
k6RFVEh/deY8et/6Qj3INucjsjUyCq69MDy1uj1f774Ml4fSBwVmTOGWdH8vjE+PCJeCpXj1miJa
7/q+ABZoFgGmk2wTgGkE9MaSOtyLbCaeBUFkBDkEujfNsR3U5y4J9Aao6nT+DE7h9Hc7zy2L6V2p
kJXKudiBEOMTo+QrDax60OOtAG2mC33kQSdVrwco46oRun+Fnlg+0D9Vuq1EEYctqK1s+5FYxXGh
n6MUkMWvQD7o5I4qZcBUyUv4ULFwDW3X1le35wBsFpbP+0dXa9ru2SRq5cula887KZSN/Fuizzut
nJ0gsnwwFgfvrU5Vib3Vmjs0acKbyk5DvGWGz0w8sKL7IE5m9FOSGsArsB4HtH5g5hDBJ7Dp1+gx
D89kfvkx19UuLddUyKh7wlfCG7pDT+JdAqiGj3kbtBE6TT/YDZYLJJ9opsPdUhI2FZlZAVBp8JBK
fjSDirPnKf4mbwOqY7ykKjbI5Nk8CFWzm2cHekGxtQb7vCf1GA8TOt3c8b2I22u8N9JRCQD84R5F
5kByT8L9mNS1KxDX2YgyWHy77EZ21C5JlTubwvIfSgGJ/kwZ8ns45nVoXCML7jdPaQA96vem6TSL
hO51xFFYp2OtQk4x9ilhKPvGlqrVnm7l4hOw8qvDIEqUFbStaRckDqDYNQyD0q/fBec4sVxCsbJu
yZ0ZTUBtSZtC04TycYczjp8JbPlY65favpqcnUX9c+NLbf20erj3AEhYJ98tUZJ6j1Bmc9/+ahGi
3pRKvFaIA/WZfiy/J7xc2VM7u43kGyCZsG2dw1oyy6QPIalkLhbUsH82K1bkooMcoT1LWF1tJ+Ou
KZxq+XmkXlu/BJT5hDIaMSOK2AMHGI2FpcjT1m+V6qUFq9TD4mHL9NCQWAr6GPmr51xO0SvGTgQB
MRPHGQEy1oX+ZSAlM/+rNFcMrQhOiL2cH+d2NNQgzrNKXc4s2HzKe6okioh1iSyRjsIWs48+YJu8
j5FgEGOPiqgc6CXScKLnx6tcqHIs+E1s+WTN+P+L91dEzvpwep2FfvbO3RCDJLb6D16fCp+Mi7oK
oUGjhWztIv1YXjMe/yIz6aqrvgpTnPoCDAZrEZsBWN6yQeZo/kcxW9xk6cCcluLaB1hYFmkWh34U
PUHGwg65c0kB/NTSU3kjYR7/KD1zu9YFMa1CNKdtWOmQa5Mp7OQvHx9o/VApG0xRqX3JOc0XcSRu
Q4EbIm8EYW7bM2HExNKCrsP8DK/BDc990O9JSpLsVcKNoeIbW6e5GR5A9MH2fQiRMxcRVkPSTrCk
w+R/V9wPpzLs730szjy049mI4+d466PJwIEIOo68NFpJ9b2buOOu8JGk3byB71QGO9AmiD2xhCdm
426Qhj///K2NXw/Ux8BUh49ooCjliibTlzW4PW2DIT7UdcWfepMmk6lIFkHRvqiPVjreQ9Pt/lJP
y7IGsh8ETGtTXuWk/dBY9fne12CkkvJRtdSI5IDm+Ujd0UBasX8ZmjH+b4Hk6WAPmbFbCDu9O91E
7w3/3im6Yc/RQKxTIxnNs5HWlIHapeOAxtUNhpS9jZqx1fqQFJ8V57XyfajBT6Qk1IW74uLb6XWj
O3wgtL5D9B83zWxOdu5JrYDVUsN5dfCUFvl76g9r70IGVtgvDrrxfRRixmwU7V8/mlAbuST9X+QH
EvenHO8RJtp03HX9Qd3fIh1MS5KTd2r3X/5ghgCu0qV8g6lx932QdnQq3fprpPl43lQSQk/P6m3o
BO95IGqtAT50/OtC7TxJFUZeEVeRiYz0gqUPkAzZE2hL5Wz0Bduny11NnlIuol0DfVzoUUrVCJFy
d3OErY94+G7kzuqOthtZuhAWK9Q0IreSNyA2Szrsiwg7Qoi0df7iIHegprcP+aD7934uCTvqWD8a
5e088QLItbERRDCi+Mo3vpiEmYXZh+KvFo1B2flgvqzeUn/OvJvRFgEWa5vDVBl8HDZv5GbKFumC
IZ5tCqS11F9NSJgx0E5o2qCvVhS6pM1fIOTooUsHiga9DieX/bJlXzz3u87ncvqUWN/A56SpypFN
lsKrSX/7gT6zKPlTzHy/jL1urmBpt9XgYkM0UWn+XfY2kYGdx+4M52n9zAqwuVL7h/uebHz2if5A
gobQv8AeXZ7wgnKtqsGLXaQmkzZY+QF2q60wDBb1HysoOaTukva8WVmE81EHvh5fQLVWylNz9GQE
F6ncQtepU7yXyireet5iyIB+6lRzl+8GEJRYAhq7dMfFk166VSO66HdLfhif5WwL9c/n66Tq5s9O
akKeeVK/igUMtIjKSMfPwT8bhbHuHywLfbixpcHdJszTl10Mj8XOqXEEWLzzG5kkN6jgjqGsfMtr
CR3EASQvd3OjJoNtHK4Ig+lDCHlbxNAAgFU0yqfkpMq1LL+EE03UvPDWgYnOoPKZFbcZ/V9v0h9X
UgCfC7NlmZJxrR0Fv3ZV0rO5tXp+cqc5AUfNDnDSMjp/EFaGt4N/LbTyfH4MGzZ1LI87PLpBWQGw
jmbCJ8HMNqMUsH0xCoaPFUygySCjBZpYtNjtN+Cyp2q32uSZeiZ20bMpVS0AM8WDr2T+C3wk5Raw
QMP3awd12kyfU2dZJamSPJk7lXeeL2Xl6jr+ubRvwiUBUpFc5FnNbrbesTkNCPRUDMyO+fyQT05b
K2dWz6yZNHCqTm32ywdG7He/IzVHi2NLBpOaULWGVVFd5QT8m90KuMONhPgxyNwguPbI3xbaYajc
rO7o/wQ/ZOCdJGmk6IwWdmT4JUQNkF7OWdK2vlGBxCP8rtyHYQKrnfA0pf6cvUyoZZ6OSzmH93Zm
Hx5h1gjfPNTu72GYHZmsBc2+GxYYiT/rDu67zIPKdNv1/MVyM/DGxjPmLoOg5/U6Atyn0PndoSKg
onl1RE2xArSpI8broGXEwath85CE16Jk76pIBm5ski7Zyt8zVYhuuSas5lWrws6V6tCxcPXSJrIO
Gu3L45o+4bXGxl4fuRQwepTzDz7yahxHnkr08xVrtXFd/I5nyXHe12u8psR1ZTfRruPFcGnplcz/
yzH9sn0xCsf7i+9UaFKPeAqecFn3sWO8Ck6W1RkszvO1vrjfUZdAXRd50HowICLxIfM9SjgTzowu
INEAgIF8O9fqbqGvUHQvYA4Nc9In5qjIdx2th1adAl9CYwmPihmNs4zimiwAuJoRppUSWGO9+7rk
kHb2ALT2gBwppGY/wn+oQkPs36Jc5FDX5Z1Z+zvizVwA7qNDeQbg6beGKow1nombLJF6lKZtYOAM
5NJTywfUuHeFumdoR74x9m3sr9jGNYoI/C1UVJ+DrMtuwpAW3FCpqYiLkUSwJDo+eDyARKwB6lo+
OgolHoaQxulwentqtUP7mv/SbJ0QXTJYsJ5XTlJNxabE/OEJjUitraV3w4DPgm0j4ctFhN8BodyV
zqIxYSr5N5BRZzWfudm+74SMAVrJSpummxF3Kn1StKNxFDLeXRIC1kqBqDJeArXLoJ7g2Kk4sQOY
mxi1HK31GA9/sg0AOwbTH41vf63Rpv1RBJjP4/dFqnNIAjmQnQ3EMOoR5sxzTCptR61pkJ9+UaLj
CgaVziLf4DhM9d/hQpLwnXgNwBWBwqQ3+0oxb57/6xet1UzUwYbl/8UgZjV54KlNYp0SKOP7/LqX
VyVawjy7YRmJxQwYYxNQYLI1GJy3/QO5Q5g5Eu/3qlA1sP+aa+RiWe7t1UPqzlNC432HPFxsu8E3
I9L85bu/1Em0dZ87eW/NPfaZZvZKgWJE6hIZ5fNF81cmCul3+TL5oW8B5p/fenG6iveVLCyuaffD
iFdcNvZY8hBhEaXfQzOgbOphBbRLMOig8FNFfFUe2duRIxlvp2dVQLdPmv/bKTkkkNYXcp+V6/j+
5n4BU5dFHM/gi1AqUeaZEe7P01Iaktxh2h5lcYrdQra/PnSpsQ21F+5QhzsLYa+5yB9AaTbt38fL
zWL/ZDKPhw/oMGftIi5SynvXdHm55v8bz2HKQmk83NXnMJM/o3aXBdA/qzUuPYpQb4Tn3jqaJn79
joApM4TYDzY83VIt4fRCttPRh9wWu2dgmWmt8qc0d+og0yVuZ1YrDkk56CkC9Gqs97hX8vQ7VlsL
MHjSE+/hgfM84OXL2Y/t6P7AXjTTBgWVQUqzoWXWksjLSJDSheF8cYce+jV5xo5/xPQ8a9kDDeX7
cm08dm9xC2uBBoKPq9VctMtEnF6nLSTMBK4OMJai+hXix0wsTh0ZL1a5q+FkxI3BmjiDb5Fo2Y6e
ZOR4CdU0rU9yGszfiOXki3zBgjrKxpI4KHHAhA5tGUPUgl2bsiTfrUpqtn1h0AT+01gsp0AwTMRK
z+tYhUINn4/sqnZO0HuuEyOlZRK3jmS7ShInsErrUBxDoPzJiHykzCZO4Z0cOfeh4crQzp4//Bta
e3JWc+G4V0pazxpCksxViqiMzr1rbYDXrKdjqm5AwDdYO7sco5Dh/Ngcm2HLKMkZmj/L5irkT/Cj
ccKXGVl4eAuxAVpoLaXC7VoH9+oaQOG1enDKCUZZ70jxnafUN7Q0c3vqkbr6F+e7igz8MWphslo7
jfc35RzUSw91MBa2es7Xn+w8JFpKQB46MMkYAX+LC1AMDyO9nWtbq1BKm9nNRZMp74KfaKQE3/Br
w28BRjR23RMTUEj/OO/WHQ8bVAU40EeR7m+qu/2hOh/7CZY+uw6cFbTI5mCuhQVwqa/I+d/3RV1G
b4/UYcWi4r9zkYxWhFrERiaGX54rqRwYgnShRdHa4vss08U5cvhAd0lvFa6LGEn7ACE6hQADKwLG
09SdxpeV5cP7VnWvvA0VyMWDn+cZnaB760hYTiIZ1yVsZ2rhjRnMQv+4d/mq8ZQcu9WJV8P0S55R
GIxPylR0dtwxBLw2631jav62JmLoRbY1dqlRVa4dtEfcBRJx6LrRC58vrlQ6dBYwDMc5yNUcuBDz
jdMQVVF0N1ULc0rf9rk69w4k+ybSnuUrq+KqWJE/4oVvgoRQ+WwqDrKDEpQ0L6fnJvt3R4QDLkRp
eyUvdPotxWp+EdWY3FbN8GUrQVib1a1NhSnmo3HOGc2GFBB+xDmutaWkFqiWUQTdNfO3Y7J3KAdg
X9mLjVH44qoLZWZy0PdIOdQNCkFuSVo9BlU2TXoSNjUZRGdDOhdiR3cbt2bZQvUwQnz4NCDwWHcf
udQ40wq7gQkT9BmHMm+KY/DxebDCbNagiVidyWfxxD4mypgLKCshp9Hw5Hoi3YCYk93cX/3bi4ip
GbckepUfyVnQNkbDlb+4sg/IJPRHlOF4qRU/mUl1LNHMp2eMc8pqRGoe/nPE/3YeGdAjJGtYjv5c
5WuC8rolyLQJmpTKVxQ89n+JbqpvcYcmIPiuyQQTvFoO7acu5YDGphieEhwiX6C1u4Y49jFDdITP
2kD1AEjZXGEfvg35h1UaRhEGQPTZp/1aNA9vQ3F8EbrHlwvP03tlKtqwmGGEOly7oCA1PijqHA44
CMZ0gWNVI7TNr3eNxcWXZzYnRL133lfdHK7iJXcmVEr+es3nxywyzIc4J/3h78jS0EWi+fK4z4Yg
jT193KjO1u0UQoRVcwgqrzMsMCEm1/sz9QxetmhYpMfl79S9iz67mdrI4M4dodUxECu21oFS/Iyb
z8Cy0xbseGNRyVJqLU4gzGBhANuBZDuBPRJqbxkcIzyuAOHCqf0gqc16wLrETkAqWW6wNtFGLEv+
4YiMJCg4Q9mcLmlC9StWEpcp3NnGujDOV+kiy1El8wqe8nsCaYbr0KWI6g8ynBkGDpNHf7AwkHKo
i2WN93kwYdgLOEew0FJ6XnAcuTOGpP987HT9S+WN55U/pF0vL+9bdt0xuu3uEHcflguBG3PTScEr
n9n+4+YtDX8U30s2py/d8SFZikJNNi34fHVQZYsRDQKmsnQ7h3ErYdqWG+XnHxjd0Iohy0auBod4
Y9TB0VUNV4S3F20pKdLRCrgihWSR30mNgMFhkuaFlwuEsT3h+SyVWjByo7OOUS9nacqTS/FldG8x
qWv1nePozpIo6k5TCjVT9qIThU9+gGQ6sqS9avBOJubN0w9P2/D1cjR9iCWhetB6GkE3m8Fs400R
zPH7ymikwRNC5dhso98nrNZUq0dCFulfMrSaVnDqYZYokhNY9EBOyBRfWnMwBmEE+JHmLDpIXR/9
uxb3za8qPNuOswgyY3MkCOvukwPy2bVOj8Ix5HrtVh0XZ+bxTd9lDbVdy5wwB0c1M3q8pqSIKSfv
m8Rt/QPOZGv3/aX4EJzOEXH63Pojar5AAS+a2ez0Vy1kWzs0Ya6XdeLZfG/1AuW4Ddap5AhmYluB
UG9kM7e1zK1zH7SjcRNzS6wOdZyg4+8RRBmsiymriUpGkdCf+AmNyQRVNzNt5r95qFUpkdZm+97p
BVub6MOCU9TVM54uN6XW51RtvnQA7TdsWwSTWd4twI/6hz+4NIyhutuuv/uceJGi24bBDPKEVJ4/
hvhRd9KWkpTHPozug42G3+sUTm0Wu+QzRIPC36aRv71dsdVixKlMaHYxTAcDHNvLIH243yBgoOTB
9pFHHXFBHWs+/RgYA3zG5A+87B39JlpfQRSQ+yAVrHBxI43u/RCbx8kU1CVWevg6xtO6Y5oKP2jq
1O+Cr4ZGDRtrv5ig6nIW+z+dvxKzkfIkgFEd41N9P6jcjaCKWpmshvTZYuDpwdrw23R2F0LYZjak
czjQLuW4wI8VDNTl+9Et/3nCE+69c+iEgTm2OSBThRRvlNTl86M0XUQStSFiELsBH9DoWgEY3TSo
qbd34JPHZpvZe6gN55qcewtTlHwNEZxnu9490jMEjDUVjv899XF5k4oKKs5ZNU2pZzHKsQVuzaz/
IXOyF60KM2CUwF/73vXVbrDkv4h1wAF+POC9/qK+cyhBS+7vYEeiMpFs/NeblVA330wPGalpwSmM
2jvq2fEAmffW0KPC4NjULR4icTyoG3y5bmjdWf2qgz97dETMu7ZamOZ7naROQvmc9y5bmVVoXqfl
0HdjsoIoaO9tdayAVGYtDSE+RRdLEAhfFl2dx/apiCmd8NwfiQyW3/tIncxl2yWATuk9w8hnKO6I
/s4FIspw1CTwnRTRXhv6q9xymgPKbaFZq/mb7/Fi0I9PwC4eCvxp2Zb6EjvSndw/ibbx1mhf/eEw
EN+5jzoEQhlPIeyphVaFrWKZOxG0uJJ6wESH6BhZBmXFxDyf6i2IOQ+CkKKdPkuXGvucTFIJH/dP
z0pN5XZES1AR55tNnlHvWK8K25HMjd49CBn44lPS4kjTOOealxKgI6TGBCglT09vYyU5jrMSe1pY
vC3Uf+srbECpzh35d5VZTGmvN9sNX5NDkxFyHc5EaYRGoYNH9YofyB6P4eH9Nqh458Tp01Dhbgb/
G+iAKT0DCJJ1d+CsLKcRWjt/povaypt+e9wPx9+/QFKVUhfRu3Qdgv0eR5cqSPv6VwOG7lIn8R0+
dv/RMhcQpctwOhWP9b0POohS1v4x4JAjffs21repViNa6eR05kkTGMLS2VJF/AItT3X0RDWv/bbB
SgccoiN3AILneMq0XdghRT1a4J6/n1wfYFNwXKgJjKMqoUxBJIWO1UK4y9eW/aVZpK4KLltl3hLh
czKAruEmlzih8p/cDIVLJ50R983IWhMvnbKinabQCE60g5XTCO1vUE6MJP//J5kIE21ifvFK0JVN
+cXzCRnKbs1JIZOqTFaCdlNFxj3+1XszGjyjFD7sbVZJeZsKk3gwSAwfrTWnfx4Nxu8oE7l/tm/l
HgPMIpHj7ZFlVJ4jqqBkVnxE7uos2eUHYsRFas9sy4L1HS2jbtx9NYkUDUHyD9PwDsSYw6+3J3X1
a8z5FRY+CeZ8QpIAR7mfYoRp/HrXe3WG7hjHY4Rl0ZgAVq0qIg4pjDy1TJ5HxvQZnnvTRIlKK3Sa
oSsCpfOndwqhaYv0PUFB2ODy4qq68Givz/wkyI69V3jzt8AW5HToxHBAMFNQtB9zKnxslT79r2Qt
ijAlVFk/LmBO+dWqBtV5bcvkXJZhPL55pc3klYzv3tgIlPsNBrQFBaIjK9SOUmOuSv1GJHQH/5bg
BCL2MBvKNsJ7oV1Z4Xg7+yxrEaxlFeQLDIolI2swYjZNXrnnonneIvMJO/+/JRBA4iFNR5jfcbhV
FRVsitIqWIO3zrMwiDtzdGLGw+/yIFbVI88cUi7IcesqT4US6SybdKrLcr3peXnohDlEvLUhc4LC
pwnGeqD3SDds7bkrNuAE4nDbrVz6ZeR5DvsGEzDjGS7eCV9wgDQRVvq5jaXb4/S0wwq4rLN2Tta/
d2ysSM3ZAQU82POX3NhBKMNpTZ27Pe6OKo8q5Zeh6udAKLd5ubPeHyGh+GZ5PijJW5xecDg4nsL+
Vyr5yvv239T06AK902+i0LQma/zVe552vAhfFCl3p2dDjiI5YgQANtCf6dbQOf9OZlFDeCmyqEm1
nUC4xpYA0zLyvqLJq0RVQ4Kj2fc38NHEbMN7r1srZG1JugOBzFZ7P5oBC0oGt2H/4n92sfbNyJZV
p/BGTbvOBM7dyns4FHH3FUnUy0BylrEchmZimS56X82QYc5YJ5TB5TMcq3s82Mnaz2+V3+NuQRo7
9ogNgnDN4yN33BQ8ojRIk+nK/l0MD2fRanLNJ8IMTSerJtzp9/xCsBzpkBKJq+N66wJQPDM94oG1
uwkAfZt4F04bXaobqi/IpdruYizFPdH5kkyiFkT52b4f36hatPz8eJlbwvU30UFSgo+6WD/Z79h3
vqEF6TNtJZNWam0puoMm4vpecDvkpEx3qGTDyymo1JqW5Y4RHNGF9e6WpLVp1bi3LIwFGUcZj7Xp
enHP3ojc5qwkikU4My0OCeXYcsNjShU47wT+ur5wQZg0KP1W5uuQx9t19zBdObEq3Yn1dToxb/XZ
NcMGLejbba/53YmRY8bOgKVvGI8rlLtAmfbqww084naCpKhcSaBbl5yd1AUmKiwAK05RLoHEHUIx
JAYonud2KyeJ1aWD8NTGQP39a4fnMEdpV4kLsbhqox19uhOVtScTErsqtdrcrZodK+nCFfjsj4Xp
TykfJVtSsls23L984s//ezLNP0TkIY7TblQ/TSIymLL9/I2jio7Lvca5g/Bta10UV38aSCzcjXdl
XCU2ZfVgxGgChgjeKjx+SIl2IJTtSMqcYYggJ2NvwGhuD22HpqMWSSNeVgc1dl91au2z//PoYsar
uohVDWRxly5t8bfBh//PUFFt7zCXnH9QaMjbFonDwrwYTArNY/H/NupZHK9y1LUbG/b0lYkMihWh
jNppHN3mlUnR+MRtqO75CfSCTkHSGHCwJ+q3kXnd9/5ygLGJlNIFQaxMFgHXhII724aukBmshN/V
v+nA2Fj4BOS02ovPn9ClHUtYfm4latMd2K7pJ3mtQKjjY3opTP9X03/zjhxcvDRqqjmZEIVsdpwq
wjLU8wMYN56WfCQTb8+LljG3Gin9NEfItt2A7iqlgPPgAYNbgmWNe3gATQ2m7w5xD35TJbNBH9UE
wqhEgg3dsWbEIegDFi7ul4bLC7+GA4dWJuR+GcfGITOQS2j6Bp9uCEI2hcVroFRXSyp8bdxRlqv9
/HPGYVYmFaLbn6qJvZYMGG9fpUzksihbCJ4UymzVI+Dt9SKaeYcjhJouLycnRO4S7D9UOY8dITNI
I2Jfw98aUIfLArEsRblhwbrbPAGL6H8bIn/ehjTlEliczTJSCLCllLyYUvRauRefyU/closGMS9H
pbeEI5o7EcRz68pYtcDdR0rnhOElBqlJboWBrhrFzqXSCH20F355sCQotDXIBcH98ehs/zxVJqtm
cbWhDgaOpa8trs75sUWWG1BNvY7r8YF0T5pXzYPyA5XVVMNMBrmcU2Wr0OYzZjxJcS+pKn/XZbGo
n1luqJ8Ch1ZM4t9tCJhnpU48yWQwLWngUmb1tH0zV4ZwNiAFy5BPWxVX7+/0sNr5ssG9hjIhgXcb
7PnJuvPOz4TVsLh0/gVWxkYuZq5GSDxqsI3y54uhA5kQuUKk8vylFV4VFp/MkJgXPjP/wLCWm3zR
fTCuv1Cbim//9wHfGbsqTm2KoR8R/uRYm9W1qnu1leslcvPqP8u4A/6TbV6ikNjn2yM2tugTkyz6
GLsbXk7IeMoHjvFQ9JkHE2sqfMotF2n1ZvMufSVBj+s9EgMsfYIpDVmYy0tt6LB1hCuf4376c8ZZ
nBjOkGZrNKbUJy4yJfW228fKDrOfaWtia6BnyZKBFGohNMh4UF4q4k8U7NXrW98SCCo16LKl3F6w
sOi6GTGDrNZB11d/IRBp8UPlbY3j8qQeOG14pCeAbkc7zPPoST8q3YdlUx0rEocLcwmY0wG/zi1y
6IYXttzZ/7oa0fIXdzj73xB+OHtVnbeKihN3GHE52IQ6S9j12qIOC7hEm3VslO8z17uvAQoWid/A
aq+spAMO6e8YbGwKNQWRU2/f/2VJgsb5Iz4NsYDuXaAsapdBFiAOI4U68Sth32p1TJ2S4oOt3VwG
OZBqU/ULkLXWkimqsu7mPCuxyuueAqt6vZCcKXU0OWNmcqMuu/KM0rETu19X3UzxIpKFdb8LLHJH
ngP0smBccITU8kNGmn4ktpzvFLUqui2t3lFiAgdPiPN7xGJEMwvd0XYwjzwxwc+X1c4q2N6nrnYE
adKa6zxKwSgIrceFq+Q2VHSqEJhEZkCJj3rSXI3J0HLyKZ56dsda0tUuKyusCXqohWzb1+wnWivt
vs9ez8qwlOY37kwlmc50dErgj8L3Bn5+tKYgBpnuWfEPLu8ltjYgCYAaegrirYco1AGWC2S68/4U
Nj4VqUpvvAtET+217e0pXekleYxx6QywdFFpREogbo1y/DVtfTWSiSiUfsygDCvlxkLsLdYVv6H0
Wlm277OtYNIQxdfEp+86lqSdk6lWbGbxftsriMe1kfEUQfzRSRtOUIH4/yJip7MxEJtYgD4nNNRg
Z4J6Rg3kQ2keyN4WY+ggLp5wEX9xgliopGCFnmLkPDAdwSmYAvACGSC5O2Ei0e5XvRZjt7E8Av9a
cVe1CVacBSoj7KBMwir0WM+x0Gkw+9fWsRfidNQ5wT+2k50k0L49AImaPhVy4IBIOnw3CXhEzmHk
earSOiWkB5toEev9gYMwNacfbPbgEy33OStjqzJzXWL0A1cBfq/lq70OpynqAT/iBMvRll1/iZFI
lhAyqmnd35A71/g16ERn5Flq4qwnfethjHC12Z/MXg9oGZFa8w7dsGTcF4N6IM65/nKwnZSlI8s5
zy8TDopycYm8IPX1ULbhmAdSdODpHiTVyY1lZUKpA0cXCya6BsdzHMgAsRLrZP1Kl6t/MQUBXymL
rc3FrMtZsCHCu8wTeTBeCoz9VGqZQm/60oO32TjqImgnQm9fm1F+cEdkBpVl5H+EciSSUtZFHjkf
0OJVOnuvdzELwCacWV3vkusbSiYCxEpX8Lv5U9Pq5I3I/xh+63O/Bc+qPA2LMUTqSFIAGD0EzInV
7EQ1ozucmkChqixLfJOBd+H2MVWkYmamBM8B+ioffozLCkELZp75ppShLPKPuWeklXB+mkAyuH9u
ALaq8QjV7oNikgKyDAoZFWtKQP1gNtv903w47XA6naeaiNYeMlWDoC5SYL+rsE5/RADuhJjSXIuW
UMSsQQrqQQs0RXKZomKw05ma5AdSa/mI/yas9nt07X57J7oqZLAoDcGbMx2hPxh1krgYDpPqWch0
t99Co2buYGEYIaw8yX4PoGHCVlfQppxCDR77CjgMQh0cjUAgYz/vjeXjSf9xQEAYvzsy4nWx8JdW
e60AuYMipWapq1zmberOXrl5XeHvsnBHDtLoI4Znd98g0yxa6r1r3I5CtcLQREp7/rJzixUxt8Y+
XWCu8AOMNP8OvYyL3riM1tClwPD2GyRZD0RaZrBzpdPD7XegR+/uPT92sjYXl87iLdhxTb7n33Nb
xuWTU+M6rOU9thqV4mMYCcCmEIiSjKneyGShZ/N7fbzXaSHpueMc18EgykbnLs180ssa6Lw1+0Rh
GQMcyuyTuEVuejsQMcqDRhVfIUCEx53d1pby5Rte/aEcgMUDKb73x6u1yQBElMdfJHEAAswGwAnU
URD+nI0XqbvKcekqKopWVLEctE4IK5cTqCk5J5q/Bl6AY+YEIIf2YanLzD+JkUHoizkbn36HHoHT
5MloKZReY+7lLkN+jZnG9d53pAafdzZg4SwWqtN5805b2iyea546FiSliUxJBR3n72Kx8b5+qXlJ
QnCd0k32LxzkKJ1irQ7CUadU6Tcw21ltwe/M5a0R1ODC9krthp8n0r9gX1fEeHdcqUIoZayEHnT7
2MEg2ZnHIF34jQ5IJw2GSCSN5jov42Y5BWJYl6dmWBaPWy6zH8E1GSGCIhBuBse66FSDGXj9cIIh
nogD0aAP+hXU3Ke8HhS1Yon9OGz5nKIQ3sF9s+HfbiAHuW3YntXyJoMW3jjcV6KXoHABfvELWiqi
XcG5IZwHEAzPJ0ww5an0tgmZ+vQ0J2mx7IRBfinz3xa9IEIvqwq5e6dBhHyeU1A6rFJXbWlYkgpz
K4zl4Sb8jscjxhJUFOpZLe1YCDkTZ1H4ALPfThnwG6zNaO0jO1Ylmutv6Zy+4Gm1qAXmCIJlqo9R
Z0nP5l6EEFY5Wc1UfJJ/gLFZDZj4Y14Fm/QzW0RUkn4TbUbTmN0O5MHhXdlkVbWWh7x+unGblsEC
ps+CdaRlbJG0NvOmLPrG8AGjGYiIiXHNaK4UVFXXS2OMu1FEkGH5bjtElGLMvjfpfGbEfNfvkHGg
qtiWWPLoBDai7I9OGwpcjBgMHdUzPguDJtnfUzrrBGUB4iXvEPRr209y28O2V+Qryli5QP9LCjgZ
Yd51Bw5VIDxlZ0WKuUfaFhgsZQ3UvUhy4afXTu1Hf8LsPhyRXtVnfiZypbANcTfDKjypW3lfOLd8
DBj20RRZOIf1o9GTm0u0y7QirkRvKbtGW0bTJ5JWvyYCP2cRdkyFW3QlrR+3WOVBhm6fh8TtJZjL
jEenhVHRWV+68P483Cy6iG+zsv9XPApqtr6l+M26tthXTBh+de182iH4Fq31mRdI0LsOKixWVios
BK1y0EWff0qdut7nbKLTMLQXtZEJdwWKMSRha2rOKLGUI/ucRMLKDrci5zQr6TzSZdkk6pbXbsJD
U7ZzyYz15sMTHseEhwpyyxAIHcuSIMRRwAuxn9FIOAQgTcpWawjpDgpbE7MKTnoLVLzmJYZTXaBp
vEd0KpwUiauZvN/jO8ASWsvMON2ANco9BYdi+AsYSmQL/mI7s0ji51cPZ9wYWgSrFtmnER5Ivk5F
dZjWJ6O2vW8NDJ8G9GGJTMbgmTpGV8WWpFY8hAAAQI3B8AiAwg1Bk9aUTSW3Rsu6aCbdQIr1BeWQ
+itdnHqMzq1er1XKtHcZqOt+aiiP6MZRB9i+uoS8HVCpUiFLFhTCHM8UMtYnM9AMZZ9NVZ4H3qDD
K5XDmo3lgZ79Bu1zFcRejltx41XS849eX74ivTOWN71xwwcn0Zs2Yg51nI8fVI1n0ck7Oy+qx7vI
WW146EOxqL23xkixoNTdRSqzyNCvTll427boChKfuQDPmV7GajXZMnIc6AUZfUdAT8eG+NLZgENB
pbd0kl43cxd+hXP1SOczRAgEqcMTWBaL/LfB/HMtdDYbheSvbiqiOmSSvqo1pLyu9uASWkQDhKwP
99XsJg//qvPEYwrGfDeQSbOc62wwcQG2EhKWdRTAphhj32j+8sl0jlugf6AvpeiDZ+gCsoZNY1oC
4NmaCBk6dndyJHrY6T2yhpMQ8HZKepwiKP2wZKx9FfzUIJd4uWy9AuiDWqUVouyfd2mXTQpqL4ag
U3xY1eFBS+xFW2W484nnMlPGUK3FmIQhckXqC0LcnimpcU9P5S61ttTQEnPw5Xjfaz3yZmkAwqf4
/2KFsRlhmY9/tQiodUGp4ZXsH93GBhMiwu6l1tXD0dJg+j+zS+Hnl/fPmEsL9AKBdoEHX9E4sxGb
dFC9brYch0sEwt3LGDSat4YddUHsJjB2EzTwpZUEQ4Gu7s+HZZH43u299M45D0UW0SAF5PgreMtD
Q+Fzmqoqykpeu3ciWelvxcPS+42yfWx7sNnmvfOnYVnr1gokT3FKi8s5wyYLjJpF2hjHjvxLWawz
sWa+2xNeHfYfoTlUKBk9ak89zR4+BgjpwkTjxDxFkML3kWNS2Vgbph/twz3UOAWulfqQ9nSj+8F9
Hgi1T/7DEEqk8pS/H/O3gwW7LGJpZTigazS66Uz/hT4/dRYVy2FGj9FVfcUXneRp1PbMuUVvBXN/
F0kTck880ZyrQiEA5CiJiaA+rGmDvZ3PRtueZBgi9Y0jF6HsHeT3ELi0czW10ZWwINAN2r/wd78Q
Zhs0FWSrtCXbgrw7FDo3MgbSYeqvI7GnYobryc1/MQ0WhElDWKLeZQZqtOjj/iO+a3wnK1qdtY4M
5EZCrGURys8gmE8YyrBS5CTNPbQtMqviwxJt0iK6TUfUjRv3CiS+Q0xnPA7QfNUXIfvYvL/90Vhf
yTKyH5TZm/T7PNECvuZQLI2BU1JgIOQsJNHnJLvLAq7dEl2DKGriG/Zk9QDXJM7Pm3KMFzPAnFkj
k3vmo5uHYDavRo3OvMiuBWivtUKFvo7v3iHP07DqPI2w/Nvg61wOsVgHKMpW1NjLFrev3R1EaXrG
bnLgKqfP20Oak1A/SBKJAYF9wAwGX8VbjQ2Y8esvYwfLGD/68W0TDHhgHy+74al/98ttptHqUoZ0
cHKi2M6OFJ+386D96DM+XX0P2tEG/HkBUD3mS/YW4Gb48kypjmYEEK+PKkaz1OlWsRjVTp/ZE6WP
2dhpZbe6Uq6tz45VczGg5wn2T47kH9nyEFmHgGscwKj7WfmdQwluaKUtG2HyxoBNsbI6h0o0HuYp
IHO6TackpFgtNKsIzycxhhS8EA29+e/YsnbdouaRsLI2y68mfNujgaONtfQoOZsQSVt1SMZ36q5H
eytfBH64BZoRqQ/MwZ8wrmKOZLhNUtMZAPQt9zEMCIENMjUPQYOhnlEAzmS4pCtwBXeDUFeukt2P
s8Sg1vLGZmmPDg6JRPq1t9I7bR+LrGCr/soKtFPOZnyumNFAXB55YgplUZT+NwNJcSSWr+BprkfU
UPlxbV3CzvvukRvAFxBVH1N9xqKSAisvA9NCbZzxiPA0mbz5zuzKyA2zNyXsmYt91PPYGLEL/9Sb
HFZxB1fhj8SB/vfA8TC6S2hk2LAvJTp1cGUcs1xUICeNaSkhmvg0vfyf8oyJYhkObUcO3aJdcy1Q
0qzkIcz37aWBL8IA8PqRXtSj4wPdLfDvPPQt0KjUxQyHIyTpywHclHpiEafRGs+hHIQ/2QAj+bvC
GmIVniRh8gKCOUNTaFjZLAFfGkwgn5fe4HyxCCSPI+GXVmY9vAZoASW9A+p8FfiVt4UTLaFTUEBZ
Lr5qYINLxW6IpgFeyzG8WA2XLw8wRm1K2sn4Shp/ZCEBWvyRdCZAN53c8bMczoJ/ssblpPaAUxdm
Wg93Tgq6Toqcyo4bmuAr0UHfXbB4XoN0aiEWZyODNxRGd71c2+R67/W+fSUpDueXsnITdne9uK54
NyjDYBoJnzBFaYZ5POHC0+oP8mgMti63J0XxPvYat7ExcdNKnZFxYBbEEWz3FYmJJvvogWX8YMMg
e2fPqz8dlo1VvhWa8RmJ+QpMthQnX4I3hI8uLc0B937LxPnTSCgA2G10+YtMYVgBgUagu0Is/nJo
QpWXiAQb5yesLuAZI5NP13cfyUWUu/NNkAmGvz52rhxdt0eciR0h0k7H3D+jhc4JFEE2GTKbF1zn
Dh0utyOBhDigU+zIwhindLEG3PctJEvebzOdwRfl9iux6x/QD+jujgsJM+7hAsmUuHV556oM0HkP
D9YAyw24/pLT42F/sJYsKf9TOdL4hIze75YDnyX3uocMgtH8PIDmXipmL9IBlhdtrwmxq2idhj3B
8OmX75VsIrN59hkyrXzXAOjxNjlRwnpcuPFoPNn/tK4BoCC6IP2iVbNaVL1F7xN36S5RLTNPdKSA
rR39xRh/8OiIDH9YZpmnPeiEnXA/meiG4KyfNanAx9V5zOXP9PQnlbHqFhAydtsiPa7YsaRSNzCq
+8nZQ/2D/jxSZSs4+M1XsoGkRGh2uM2LmVOKUUs/+tOVJ/ANq8+NvfOcn0zaW2TdS/YrEdB9LVxb
YccxDu1eQWCLvEH40wIDk45VAgs8J7G+rIABAJ4ggFS/ULWqEcBQzKzvJwj3V+DLWefu0QHVE+2F
WZ1gMWCQ2L+kQTn5Q5nfR9L2gYSwJ1lTsthux7QUaTzCjwURRpvIXU3NOBTUCijtitqNYxKC2wT2
p5gUoXGMfcAOEjKdCkLw3IFxwck7rVVZFtrjUdgOjAlL+l6qA8EdzhqG/6cEqfliHVuL6IwGjmrn
5GV7vFzHsvXif2fEXYqYGGv+eDyQn0oOZ0dd6R6dtb0j40lerf6y1toMcPNGasOhDY2OT/Lmwojy
HYq3eLrcAs3p0UBHRY+z070tSo1Ks/I2OVQnhM749quLQ4xzoh10J9F207qYOLMhM+AyQ0M0ymgG
B9ckS8uoQgNKuVimJe7H6rMR6jvDB0uPvLzPREC7nNsIxMYt7+ohW8t7D7kIEOvyguCkyJitiQjX
i8igSLLhykpP2jGaPky64kmCxGDRgZSl311Gd86Ndo8QANTp1aKP8WVCbgDdmxR1WixxmwHfrUkE
/b3Y4iGU8n65OgTkB2XkcornhDJotAQg4SysHmJJ0OgOk3QlBjoHetl0yb+D51jCbzJvEDO6cn2t
AuYkA+WdIzqPFOzJlEyNaHoxcKet6Ek5bZVq6u2r2aMsLiWUCQ+klH9eDWieQfNe/XhWT259HIe5
yYyQ9DmIp7psf0Ar3moER+4NcWpxyEg5ySodqzkM/oq0RDVK4UdPg14OE9/lYBFLumR9uj9byR4k
55Nn0I2r4lKNCVDgYnyB+IbUX8AEcwhHgsdwJwZWwUDN3oiQJ1Plvq5c/0/7Qy4w+FctaiCvgQrc
Xhu9XlWI8hruBurZlH6Noto4KZaF5XQQPySvxCArWTF935OCmIajlHnGN8/077nS26lXGeNOqK0x
pKv9jDDbvvLDKOo2q92IleT97x3vZVgDZohs6klZMG7qimrK47nALwkFZifsDdsxH7mkMtlo6V+6
yC6x3NZTPaQkSrbIvLSdkUhRkmU5TafHQY4o88yhdVTb2xI885nB8rmoh9qv3ibMljviznnqZddS
x2Iw+XY8qQ85pI+3ixvyQHqKS96J8LpHJEexsfk+jChIP/q0+py5V1WHVJMC7aiakDfaDbi3a37o
NxBGV90StMaGv3I34v5b5czPhRhOIiLVZZhcdYnuVDFH8wgHB6kcUkfdlfyr+GEvQLDA+FlCF6js
HHtpEnVU3SR2eMhMf/bBClgOdsNOY09PGDNcdjgb77gYAoSvSt0NN2fNekLrkmSPBHlt1FoYcjBs
9mqlncEa0pgzpdfPSA4qe2hTphEZP7si2DtMdElw7sIrAUMKkyOU9uJH6rshQj6dtFr/IEau8egX
9yWCop7V3GxxPiF7yZCT3FJROQCiJR61cUPr74oLGoD3NGBN87SzRul42JCCc3nLePdAirlqhVAk
40Um9E4eruxDdTWPVuUZpHAVzwFwSYCUOoBZ/DFNrw1m0e1zmkUDMwc1OvfV1LsEjPAJvvD6vX1F
Qy14sj8bgqvr4wtps/V5wT4nlU9VFNCge+HOvQKl6N0mdFu4yY/fxBgIAVUrB9U6EVwyhMgUPgy0
VJT62+fFTbPpOcLgx7cjxSY7hRleKXgPfkrvnE1Io/787jQE4GHAYPP50C8zHW9mseav/Z2V7Hn7
9HGO9ESYnT6YRakgIcKi69maaaGqe9xp/L2m6BWhEO3SiMsGj5xCxV68vMIo6Bw+3Wv3o+IdvihZ
WIA2EyV6lFvDmAau9zgaItN5WlA3Ycz3k1mmixS+GI8zpWPFHINGJjwpOJusIxD8F/gDspWEqTlA
cF/lNRf+FQ/aEswElRvVvTwmNyhMjBD5i5xHIp7FnfwvAnooCR1ZIjZGKu9xNovB3hE8JNSZ/Ejt
rXJTkk1Xffnaim/aQ1ZVIa1oG9qIz5/Ze/78x4bwWVXmrqQtoazBJwUagtGqGutilfru6Bz3njgf
2cqWbtj1pii3w/cjrb6YOzRWmsDoWQD6KC8JShQqdF6pJdAwtspZVuscL+X7J2M9dofXajNrBLzQ
ZshN9UrnaXxdyg1R98exggXzzHW12XUYvL7a8Y9TNBRfxZtGFdbWh7jfKHtqs9BSPzY56icQJuLs
IsQQkcyaqdM04W8rS5PZuOjKyMA23A2AtHXRwAcbm/82OdI831AbVJs/fqtO7Jx/MBEuGFvX0DM4
H8uKfGLxukv0d14H+pHtkTBY7qM/AU99f3XI1xh0NLvVt/NuCnFmsmPoA0rYlBq4455Q+oOdjmvK
AvJh3+l/hQoCYoxz/rQxHrhoOSB6E5ryE+Tj4jjZAQQfhPeS0YW76bqpRfIGzebzOmVnaPBWRv49
lwP7uA7ylOF3T9nWWDJGvBL+uZaDEDeNZO5HMj4AVOtLYA6VCGmSy3egAjT71ulpRntr9+mhTxaw
XMW4FPJGAShHuCjftROyZ135RMQS7gQwIOeV6mov5EBDUhKfNnMhYYyfmul2cmB13kOoHLvd3tVE
LL2jXrr+YLQ+sRcn2nsYEMhdrm1VudD8sp5RN9YmB7ls5gWvoOKnBgpMO6f+sqac6VZnJ1Xjby1X
m63lquE9Yj6aD0VYMdEGxoLODQp4zjBA4slZEa2Wv+1Z4rbGytT2Ls8yQ90zdNc8QbkIFFHBXckw
v9FWWZAHWr8VCFyZQ4e4wyx7ojPlAfWhhSO9sI+Fwo2YgaGQOtMEWqqXXG1a0+7oA78icUdzLsHa
c/aluWlhIoqNBtBBMHaY0yB7FZZcEABr//lqrnIyH9K88OZVLzO8+1CtneI11XO7jMJTI/s6v/wz
O1QSxFGdVGluJ7LPryLJjE5WNmTGIupXgp6lYIw0slvYgcoc29oo9G7G1YKKme4DvTPRhL3Ce8hP
EtLghun7T9RMgIPCbrqpvbanj6bvKyByTOYWLsb5kkZvZfG5hXzTdTt83CixfKsgVcSCM054MdII
ruehwBbEUV0NzwzOKQJ3GvwpBLrprVfPoFPN7zmtOM6AkTxG/F50rU4yfRDAHDbhp06/665TkYnP
tazYc5ObFF4X2qKNZqEQAu0XzepDgG7nGXwBNw7fUEFtuQLUrNfFpE8szhtjHRQ/kzDh6s1oeL2X
XoiStFtAGp2flr2qIEu/HRBmI5CYD9Z5FchNatqHSQeYNFNLZN36NhiBZoXn2hr7GjaHdDzauBaF
FsMsrmmiIc/odO4X/cDCQuwIaZAOtqoEaVgRsddx396kofmONIn7m4z5RqLUxC8ssnc8jcB3xqW3
bHE+YpSqVo/M7jrEWJo1HWUxWRZDldDPR+EqginFZGJfsZ9F8lMldrwfQPs6xKh4Sm4aPtEoIcLo
rO3xqIjjejzzNOvvxCsOCslgCZXYcQI7i79QD/4X2x8RypVze53ap+rdt9QRS1KLPllh4hv23/j/
F7Fa4L6FafR/R5S3lL2vehfP4DOAnH44wYer0+mmTfBi1/BRZC7XJ5Z3qYrjwI7CD9VKE158MLhd
FaMPFvpFW7J5AkccdkcrLuv+/F6xa6TVVliOHTc4KiFzuceWljHSsy/AMyYE5FQ4puQWzOecXQ/f
JyAOi3V/ikjzbxRrI76wI0yR2mZzoDkpHTdDTU3HIcf0zBzLuecOh57KsJInUCoNKSw9klmPP0m/
kDst7PN0KUXHMKce0Cgp92yXoHV6aQ0DL+3XA5NIz/jjEvbjgOovCV4AV5scnoCDMa3foRhPRUMI
7C/KuEWaCAQvMb83Ua/QJ0RzCmrGNUqCAiB1kEEpmZG/jVwt69VGTxKspgn2FfPp2goDiTU+UA/7
4JAhL+lgA/PyrLrCyoybIgM8a1iAbfkjq47oOu/le44Y3Zs9/bTrMTjpBFKElraEUK4+rqPQIuKx
cX0zeR/W7eY0moCDVPPs56bpbuSVssUtpEfXH9TlJBBPTWyq0WbvZ3NAuCAL63tC6BQ66D6KVddh
Q5Y7oQ0FTxRhfQ8PK+wJBS1JR/9Q7KHK6PnLZ0z2fLcmNXJy+P3Xcz+EgQrAm+l8sIn9Gn+0frHQ
ZF28JAnZfPteHvtVN3kNl+E1QgOYd6XZnb2d9Jghcq6+4TD0AGiMCX/qaCaRIoIr4qywR7YVM0J9
sjSBk3vEIYOxiJ4uM/Vah9R9WJ/eELto/Qmr8mkLPMhRo4GOwuE1RoPe61dVtwq4gDJIEIgo9lmt
xI0SH5wBxaS8fwZJM2RwjeEZklxwK+1RlR/XlYp8U3saMUQh/VajTRAeLRQJgbn9o+qf7OotvtTT
I5ZTR/K4Q0D91Ws7mL7NXrE3FUv+xInGdXSzljajHCN//Uq15DgOmBOWR2c+OblI1nMeagVMbxy6
w+8n4CHzTgBWUp81x7utlFFCIBx3klT7/F7GywQRQdDIXxUH/KdrBHGe/kL/nKnpXpokvlM2j/PV
qCc9t6Ztcssf5h50FWbxQrqM67yCNoHUFRagNjTKBvkGZT6FcqrKZSPbsba556vKvTL9ipkR+G3R
yqHeYqp2Phokg8GkA/CvhGkz0zfuOblTqoVG0p8SDSD5S40269FSCbxaDbkj4o/jwU5TeN1CtK2v
ottrZNaBpKDrfqpYN29mFmf439N1EPRyzu/Yyuv5jUFnpDPW0fhCn+z2e53R+u15P2e7XplFnsOM
DxsaJbq1PrJ6+r8jEqLHlGf1ptPtw0JI6DDdg3hSYMCLZn+QhvYES6Mveh3ttHHqYw6Wi32MPUEe
9EbdLmZQuj9MSAJs45kf9KLKIexR2l6pPuBvgQTvrPfCxVkHRwZR34qktN8qPn9o0UONeUfbi+I+
iIXl61hs8Eip20rCXaALKtUpmXNfivPFFc7nJnCBYnPhXdjFLW5qGBgtYhKGRlUCkr4eR8nHf+Y3
Os644R23hFLrLsCsgDTMfB+eCF8J9vnVonPwhkELjZ3+gCnk9FraYGtnkzrVdJ9zinYf0Q7Na6YT
iRpTzR3yX7QbunqCtn8qdo7shkZge9vlRbqrIe+JfBpLjlrkh6dZxpkG6308z4pDfiXWmM1GbZD8
2vfpqflxcCvCVaGrrgWyxTix48JsfzTPMrrG3LscxyLCVPlYatIz11g14u8XrS0j1SKhZqZyuqdM
RR5Lw+YYZwNlaTIjSQBbIojuZM9FOTdTLc/CLVACiIsAw8ovNYlW4F1XSVQhmuWQIytv2+p0eoKn
VOK7ZUrCrN32YqufKPbmuwRZ8h78ygI96A2kA+AlLIZUD21kTCup8j4nyW75FQSsdGkZ16IpS1BT
pDM3bqlfEskNY3B1zeSwOAIvMRO/GOvw+jgxjfOw2ULT9xmeI84rmyhICF/5EAgXUlMIoocfxKWS
UrhAon4PLa6KsY0VVbfv1Pdy8Xea3AA4BEdExiio7yZxQ4MGwl0TdDQee/xvRVh9BSIQ1TL4Skdl
0uVYmFHgNi5tCTIYfe9EjVVGsct0Ot0x8u1Gg8yMXOG9AYOy5eHTRazUP7Yyzv/L5abnVVMaouQG
AymVAxqQdIZbIJRV0SxakDLfQsnXjMze5Vv9zA7YYpqz9Ax+3H7rDhCmSd/5GaGpZCJP66xSZe+a
RYmFyfOAiXnT4P7HgBwQAhedbTpNdP2AQZYNY5E4B9VjRsRb9XDVjMGYwkziC6YI4EoIK9lHtTGJ
4EhgYM/JJs91IQ1PNUFU72g2VsRdO3UHvqy5kaOvkITVIrlydFzdaWz3v0sBnAIkDMPoLAVYZTAO
/8strJEF+5zDh/2QlMWWUFXZ94xG+mZ22clEKevWbEmECEW8p9bdpLEVzWpIe66ghTwIJp9Iu8fN
YCnT/6ykEIPlXtnlqR5Qj1ry11rahT3YK5C+a3/KNbf2Y/6wgIIBwevimvFnj9MTWnkDJQwJch/4
6AWO1dfsBze2GN20J3ILWZWkJnlEd62bE9gf7DihgObJH0KbKXuTjGbInP1mxdmzzUxQXNdA7KOY
bsLZaHPvaYfyZwTDEGIkJFMEiYoSz6Vj6fBwTlC08tHFDAFOu0O1YyGtDNKR4MrSgCTzKLNRjKRX
4nf/aFco9CDefRMCqdH5NecwBJex/mpDxv/Z4Znaosb351aTfLbkFL+JjzsqrJfo2NVb3EjQ8pTa
38vfHJKKZpv8+hkrmj1N3K0Qdsq+9NK+RBgKk8X2c/+3e6i0zqgqgajPLr7FflCHpHFA89P9iljY
3IV6XA2pTYXVa4AK4OKuhtrjgqhqDhVvxvad/ZugV4m8AK2uhELcG2onOXh7BoslCZm5q6d/aQqA
H/JteJOYkhF87M3A84hb93mYufKpfA56/U4usNKcXPjkIl1/t8PAWf7tDWRwKpK+J2LFu7H91XiK
bwk3zBp62GvINPBeErOGv9pUZR8XykdonMiA7SXAqywILcAm0dZisTjLGI0No7pt875HvvPDHwFS
UVm6QWg3GMziTDKPYnF+Kk03aNgHuMiuLF8xZPUkb5M/O3hmcBNc/eO0Yzxmhity8b7yDtpPZjHV
DeiZPZ7bYmGL1j4AKGiuI5ClMgr62t7QENojS8qyiujFcfuZcMy+ak1/Ns4ZLXsKS7wvW3FzEwae
b/vOMfkCRpFQwFIiwZP89K0+oySN9XeP5ybqHMWbw2YaT0dgyYnfn+r01fH2NeT84cAIdoHdYn/k
YNMHJhMy9q/lF4FAkWagqhlLGPx79tliBzpTrnXQRjI2tsGvuRd6g5Yv+5O4mTSaOaAsy+IXBTSk
FKWncLJCX1Uw3XAfbQocw2ZtPy3yaKo90QUf4QJeswkMeUwJPdsv1H94q4QcDUmuqpm7XBajxzfb
KRg777g6xXQrvlZnhJAJ0E/YmBwcoq7r4zx2JkK6YRW7BBpeuGiXpw+S0MlbzquaWLM+uKqQ8ZEB
uz6NnArlE896x1Rp7dkV0CyyhTRSMy8ZfDwnJScKyCpNjRnQqdX9FrykMcQ0qmbJZibkY9G3rbi9
inqN7idYZD1xyqpEyw65Ada2F+VoTcg9TyZlm1eHM/i0Sq2Oepua28kQJYpDD8xCo+CFzZtqdtq9
oZQ+lDqAgo63Zz3swPi2GLQhihvSDAKJNM5ChBQtXZAr5cQ/AIHZAd1IriubQ17oZF6p0/Y+et2S
AF87LcI2BRZBoL8wwWtNfZ1qBIczAPKODYkXf4cBgfiSrY2Ts/KBWvVTWa8KASTtXRkhVBMsJb82
VXU2QeZFzsNK3SZax8LBCjXyRHO/QqOrGcypnvwnd/Y/vVkrZAOcPunAl8FLryO3GqC48wyA5PLN
tbRkPEj9gQ1UvAPnPt2iw15AILnAjgUQ1Y8LcN1xZhgIJFL75qAlmNiuUfkEWx8o7I6dK320ruAv
NoynRehxbOw2SIDIA84MzcmHEjJEr04inGSbI9RszgsT3s101UU/6wgYnbmBuBDxjCk/S/IB20/v
iVCWV3J2Y+ChPIzGm09UiziwVPYxxrf2M0fn8d7IwJZAU6VmfPhRvL/RWZoC2XJn3YQl2z1KGpOS
cBQz+FOzhU0UqxNiQIvKh+Rfvm5+zzO0cyxabJ+DzBlfZ622eNMWxW3lDQPt8XOGg8kvaJMNbG85
wcnECjIquWw3JwsSa3CTwzov9EdqM92s5eQF1WnKBCSC0TUHwzPKvmKbkC4P5HCecix8XyU5Re9i
b7BxJ7Y4GBcPmzF/Ltx7ayHR1NmkJH0gX9/TdCX2toNUfiqgtnMMHzVssjQovWaa90JgAfiMfS2P
/QbK0FMxVc1gOKgAMHSaI0DLzYfgbk1lxUKgFXluSj1Zw5WdukZn8KAOthNn9MiFn3TLGjjDM2Em
YY1+j6McZabyPmnY4TWiDAoWm9BXPCb988SgydWLugHwb4yQqlrKLrJ9geG+al4iE/uQKK8Jnoiq
YL8jzdkp9TLXANTf5+Xhq86fLKVClCnuc/UuskoyLvXPYF32rEYiD1mk9EY0W9dOAuBij7OcN1Dl
rrj4u8CxMMAGhqOCR8k33ThBYTjn2mF4kWgROpPUPPn84XQ4Xc/dVRsv+/o2TVkTHdo1EH7TMZyY
bGBF02Nkg22wuw1O6QSze3UcSh+ZbXI1zGgTGAbpW81jUD5baAcgG7f3oNocAX8F01inja8+y+dM
VU90FV6nTPhc64FjO5WqMe0ejMqiL+gabTekqIB8H+gfj7ROfLz2CzbFse3pgZ1pk+FvfSRgJ2EC
qC22H+dcQyrpmVG4VfDMuuRMmDUxCVDylSH0692yyYNrIW8QdbIWSTG+NOwUJeyg/XQWAaZWLOsO
kVt7vdZvPpXxbaUzYSVNmm70u4eS1gUQmsvJU6Du2ndS6sfHQ7lhIpAaEPubWMu3q9ZFi7yYRHyU
6zo6zNmh2afVi0z9hKiZ+v3BicttuHnzut+gSMgXjMHiKZLQhaK92so2BHsGyGboKgKDYew6r5CY
VNfo5BIbCY3gUYXkINLxaER/JpTUXrKgMZVQZxrXiV1frIglSkB1XHfjcRdZbBlX3DIY2hPY9hab
ip1s+7OUGiwayPcgKxZMXwuEFotF2qkHoBRsW28HK+bQqnopE4FACl+YiBvFOinbS3dyLewftBb+
oiusMqRfbWb0SMOxGTdKRZOPV83ckvUPLzOlUBcw7irxjwYcqyXCB/clsgEfOgG4yanv8mDOy7A9
Mwm4PL8Qz5o8JRIsYnlleLSCPZLYkpWbKApu37PpqNUxWzxq0zxtVUdAqPfSKBiV7OZunxNA9SQb
xrAFUwb4q+dwXkV32tuzk6VCokekk7Z8ajBsEZOEhID3Yry++Fk2e1UFG/wGVpj8jXiWT1SKShWE
tgP7aSyiY3By+OLI498TAjyIMJTHBWik8x6VctI+96VLeFdb113O54QC+KlTpjRf9V+0MdJ3grsc
xRK4fj0i/GPT40tMly9b6COrXx8qSBuGjSr9N/QQhK+qu/uuUso3UA/Mo+LPM1O0fO/prHkoLOQB
yRoTR9ohS9MFI3vRkDAP40e2XBcuebK7Ze/5xrJVipDbvcRJT2NErBXkpg7cCvcL31GXp0vULci6
itip40RWJFMFP4yudgVQq36SoSo64nPuh2+ExZGOLXleqT3Dyea67EEzkgVr45L+oTvtGirSEfDd
ps0pcv51ujUn1NJPrtLbuh+aFaPNVIzJfALg3csGzptsFZ+r5Qq6w/QwFRtVmm4bYwmMIjtuTWB6
7ppUNTYAVOkjd4wZEwzAF0qxCmk4ctRSglW0oVO1krJ9nRlSi9OWedKuC2Lfr1t1Geu3FFZpyLQT
7oDNZaV0LTNXUhNW/b6IZq1vm2TVYBkOHV5DhxWYzZAi+iqx8DX+vYOKNRTL0omxZBL3kt3QGGOI
XGqWVps9kgSPqw+n+NOEsGU33XfQcI98uFlLcfKKICBEUqlSbgkZMeMIi/h8PnueFLGrp3HQ283t
EnFFIjrqnyNUYQAz9zqJGrSVrl569PLCynocJ99hekrNnw6ylr9pKs1bh4LzXHthy8yIOetTGCsh
nrZTXKDhN/lauF9T9j8QRIoOwuUW/H9Q1+k0BTNGglzsAJ77Rez9ynObGWZVB3L4hvspWEJ/NUh9
cz3imrZGdTn0gPfON0PNQqVm0la7H8FtglVqtwnVmDkS3ja9JpIDz76qUsAso7U7BiqW1EQx6XUn
PDtxW2Bkf2/ZlXcEi+g4MsbCTLmHAJa9iXu7YPiQx5jlVbvMG7tulmzbPmEcizt66q4ytirZhCm4
ogcUWjD5Z9TAZlvvYBHff/tXrhdWdDbsRbe1upH+0LfdX4Q7IgnDiPn1Ae6BcUPj/Oz4eu0dFJcQ
2vWoI+AQOAbsX+zUJQPQO2dq780aDHg0u6LyoqB9xPT7eAixWHrByPzhzmIbuEDOIa15orcVev+4
sw3PnvObYAVhQzb5YEVo2GF3gQDR2gfM8ci5BtvlTLykE9B6sQEAN9vlGeWXhqNpUk10EVaKSnYm
jaCv7rggKmVzbgrxuWqIXCjdV6bXXWDSslxI/i77ls6RijsPoh77oIJ8CHePLHCRNpSQQw+12x4d
9RB3mxrokqKHadYFrvmi1jHBCOCRmoiJGLhRRimw5ZLA9Tw+h5y7hiL3NrNP4tph39eg1sEydbk5
LtQPpWBu+ZmbpT+aSL4s/fLY7RxNsE/hAQgzfphLEmUGaflH/clo8fsp3uvSd7brgSJ6IlwE7Cxs
cL3/2pMT5veCQZTy/Zz8Ju+RnKtokR3hvwgM7WxLBYB42wnEca6Hc055XTEBJUga58hCJxfnw7GT
qM1bBxqEGxMWGbPP5a2ZC3zVeaHex1U1PxowGDO8KWodbFFBJlOuOBg3s/HCzakRqZ8ubOhh+Fv9
f04byB9lHv91/S2pb+K6zcvJvxgp/Ep0TDWBQcNt39TONnmEhYSKlvWDHbR+31blcErTjQJ2/dBo
Bdni/SOTUSEJXwQxs8LAQLcVgsbRuHSZld0Y7IfnaroMQ+WXwBCuGz7gQxpFlUBL4OWkFW2MIRkK
yziINEazVXr5wbAHrRpM5O9FX0txU1BfoL0FdIBToPrvk/LsRSVrr/cPaEjoWhtsBPOMBTiOM2VF
W4BNyuw+XvJ3Rf9qlUI7TUL7JkmkWytIpFBJMBaLeyG7DOYuek1agSjIJz7IHxWsiuHh2H2qy++L
aCaFVj0Lm6gRCLFjAwdA+Vh55Vx5+hz6ZGmEej09jsLlVVtvaG87FMHpQwPVMSXHsd0qnz3q47lH
undDGbZ24siycLdfDX8ZqvqHy5c7Lg2sF5aMamL9pQ+5TXBYWH6PuH8MkBOaCNphiQ+P9/B6QzGw
JvEu0PQa0P6UuU9zkvJi55YvAGfMj4xG9lXJb2JXFvi5u6E+PRBQ0733LWymJkvt8tQyEKQ8qfz0
kbZ7iTDBJtc26IS7/pvGNV9iYPNIQ3Tl2lDveWpjWsuBoMq5AwduAcXny/spOrb6MRfMT3N4T9RB
e82xTUvI0bPh+jnKZ/yKSDbYR4z/ZujE7XnLO8+/CX6VEf+UBsKULITPnTdBkdSzd/mbZL62rEDC
8TGfJHxjCoSeF0v9iZoBq19Xmu1mbdXi27CZWtkbyhjhoZf16EQ6QeJvmP9GrPQCncE0Ji7HHarS
Tf40H/pLOkDa+DH7iwFdZLaD1BPcgPjJ19EY4Q7lzjzJwlAqmQ9WDbf/boBXIu2V1ZKE0J946nx8
LUuZXyO0qFIc4i+upnZHBIFQrcTiEeZ3x9/TiLsGnxt8PX4QQRXKxDlTLNKfUMz7uAcPlIFKO79x
ssipEKVRfFxnIWKp/gnQRqlhKBeSZgQO3Cy1IpwkDng+th0+VaIA1ghbM/R9huNSAE4LolpCP7xe
B/ywmFmjZG+AczmJwKZ68oawWN1FvBqZusLSD+JaXR0+ZJbZvwTwEjqP7bbliZfmyZCFMc2obsAt
DjMt4L1dFv2RQx0eOm1PvV7gJg/Kny54SE4pFhRr9Y8O2LNF0eTQZHyKLCOkedqlOm5aXrDvOQ2t
NgBcSJIhJLOmYwf6m2q1vXdcw328mUQ9XcRFSqtdo0ePyMUVInBwA6WlpA8txB6TrqJpP/VFDNKo
lViwsoqrO3qetCz1/bPZ1p9EmVS2ZM+8CetloCgYeyZjXrxMFqNvdoWv2rAEi9gqAADDl4JY9fit
nxYao2gO7i+n8TbikCJxllbd2MLpS8AsnYmdZDsfRGWmQEbwK8Z0lWKSyUARbQC3ImZ+h9xQWBxa
cUqnZHXTna9Vv1hprzA+//tojyiMknikD6+GVESepsmmeraYPVmumuQjhgpkrItY9TMU5Xyb6eUd
A+i/z1xmWhur1fXR39v2/rJyToo1uzcM6B1Ni6Vks0UNzKpKa28WmZNgW18Ix9ovney9aWlBRuRH
k22IgztijqIHNvIE+I5ljmNnISdV6+4csh5c0cL2dREL7M2qqyVM+uP+dgB7b4Q1SRmdVnELxSDs
kLxoJ6W14EKS6wcx70e3nPrkMnXMeOJLDzY60RBJwwQDZ2Ca0DnQBI61diRhA9AbGCdp6tGIPdhr
bkY+b6/mZXXJm7gwfmR+sGQMTzQLaW4dUaI2kis2jdBVAVq1w5ndGF+8s1U6NiYA3dEkaRGCG1uh
owpIhIJrr3tYVW3ODu/9MZDAc10xu0Hd2m3DIqpDKB+h5/CyJCvw/irrJLd07poDZtDeGnkylaku
TvCIdJJ37h7gabCRa4Ww1erEo89LIHWRCQvg0Fn0uogUIOpF16Z26sDnmlENGAsfpq15ssishWz+
tkKOzhVEqR9GINOu4Rc//19eumIPEVY/xSXF5v4SdrZz9JPFKtG8lZc4WwHX/nMK0vT1aA2VCYbD
SdgyHzsESZqkI8ZOVCbFKA1Ws0kYq10EmoC5PDlB3z+04xTNNRVvSdyrjLVouTGbGDGpn1ycuKQ+
/Nze+ccQPaXJk3Nb8P6mUpb1OAORqT3RQ7ecXID4ZmHCr8aWZY5HxHRXuvnPegWkwdwdSclxxKEU
KUo7GEUDr7Zx/XoxH3HavZPXjdEdiu0Z04gnYyaEkzdO0dzntMtAJwh1A00MHc2F8+DXPnbtbu4j
ybziH4x1sj2FXhP6obMtbWX8jnY/f0Yba32UuhJ1g/kon+k4CKJ9q+73xr6FYBU6RvKjre4tisYZ
u3KtwFP2ACIiaWkSfi4ILA3c9h1U81dx9oSn2dYJ6uaFllB0A2JBJ+1sycbdLJ8qHJsE4AQ6Ngj7
WfTvL1aJ1Y8hqGAqkCrOCkYVq+VpbiFOVzdqaUHN3tHn8vLODXSrRBmvmzACNbICMsnlx4YqgvxV
Zc6TIxBqae0PRmIPH6u0Ve4bCmxfal7rLvWf2xWuskesKh9QZcJIsoQhxXAS2B7DTRig5LnHQHzc
cQrGSLyn+ssVxrxS05WOXCY1KgH+iH1MMHgkK96piDgcugLRB6WrVM8tCG2HU7a/AyVirwIAWJlD
dKn+Pq7KgBcpwWvbSUn2q+EkrrinwQs0l3euzFNDZpbPQzWxGRpUOD77+oUxIO99bZS7g0HUMQdw
z8yvNS7WegvMkjhmJHvmbXSrzBeV6tG3v+IfYSLL4LBFRKF/6m4J3VjHfUXrrn7LFAqcRd0rbNkA
sVDdJaX/a/V4eiHO7pukHGlMxbb4q7dGY2dov4tqtgU/AAEDgmuitWMuAEUtOAdyjLvXbKsPO2Fg
qb5A6CTemXYVql+FRViw2Wu78Cee45L+dTajyqmKEHccYL84TK3eJLHVl/4YRbHU6Lp4fh3gGcn8
a+MhYZOYziLkQdCskTfLCjq7tsp/AC8zehWjgBBYqkt44DCuGi93B+WwcJwtJlLthR69ILCuEVtw
a18umzbjOMUeSlRd4rJpad1XOWW0e6PVDPRFv9v+NcvpOfglFvPH9mTkoyuBEL4+XP8TTq+v3jlX
lY7BZ+fChbDYqJBM8fLG+9KNnmiawigIyz73WKlv1RPVapmV5xpZwNYnQmHIkqJxXNVAcVRErHWx
nnwYCU8qLZkbDS6EINGmdNTtR7JqFHfT+uGldWcuHzQ8yssV6dXqTDQ5Pcrk5otU0NW++MWYaH5X
y4kCznxzjDQelmEJw0Ra2Or85ZO+gP0daETbWnf3F6Vlb35zgqOyoW0/xXxgxRu8tXPrgpJRKtVS
9cWJGzHYkPeyFP46bu6hJsF2rTfJz0oSSvRdLtfk0AwsCx0iiIogZMwaIJG9ifZFqmFopehLLxIA
PqFV2jN+R36qNF3iY/E0h1hY6dDJ2uqJHuJ6jf4RpHzXcKHGiAIQh4TRJWNrdv/QtpIAW6uyX3uQ
4vImJPYzF7+bLS9m4ye2YKFaJEkNi6xPoiYJrQn/NUcaZsvU8BCEEPRkqzpxk1DYUBPh1xwCNJb6
lyyxktApCxR+Nqn4I2s86cVLrRIXBYJ3zbG94nHW8asURwyTmUlzOyXGgT1re/+u2Bj7QXNUkBhf
+MYhU/78XgUcN4p3Nd3KMpFIkaZDgTnfIs/UlkQl7kaGM5r0wIH6v2Z1MmqOMAQLfUMjRNAsGSP/
71K1G3GbqxHaIE7GU01PZUYyJ3h6RGDNMEYVJa42KzaCopPZD45+5sZ97YSsWB/C6FWuL7ePUhyw
vSEfD9zEJXQjjlIIGfPfCkWosmNMOAhj3fDpg2vkLfTf8a8YRZKjR1yEXIsEMk4qKm6N7JeehqLO
Ahg95OrYo31HJQE2cblVHQUxpXZ/6sWfZu9b2eiPdsHCZaRqEYIiBY8MR92OtkPRhFsid9xHf322
g+RQ6a4uaIaEazngAh9CCBG5ioQRrAREY+6liDfWXZoPTd9H2gnShwVn8rV9MZk14TEodxQQBiWn
J4xWUM2EXEQTROXmqMSyg1bHAz3mLJ9EhxPgFirQYjLWkiORil6OA7vkpqmmCUu1J/yalXFeeHy1
tVDRTrOPx61PiRiZSKl52M1ZBuNKmDL9J2ciak+HcNf/8VIBVlIJKNuDSeS5H8jXSj9xemL3JtQh
b9SmaYEB9Ya99p9jkUyYSiW6+8OExPMRzX5PuGnGqsYYLPdGCC+WmhrPsZfpIElpQxYKKmvhgmHu
CuedTKg0y2pMagsMYU09pTC5BcoGviuG7c2/AHxU6S3sPvDLNyDXloOfDbwx5aTDBH3ZP9fmUkay
VNo0ZKUypJ4pEcHwW45v45CPEGf8xaPJV2UETR7iHiIT/MhQhpa8BhgXWEwM2Kbgh1AY/9Amp6q7
R82yOx9jNalKMh/nzoMy1AEVIo7/ugQcwncI7SdBndp27QI8n++Vm3V6LZkGyMo7IZNDZkQ7ba9c
UlAUOQY4tN4p5MqP+JS8cO1RGLd1hVLATs+oXEFTAGg/aXoE1Fuoy9abn75d8lOx7kl2SokQeylJ
tY14J8Q0OOBbaUI8NGvtrWcBEfGEp6NxlTutdvAiII92vPORzn7r1Fo0rEjXipnTndiIb6xVrrkG
cT7epxU28AwyQklwO7Lwl8IGgj3akrLZDkA1pP6s9QBQZtLSKNgWTv290rW3CpaCuABCzyUrvOqo
ozCtfwye2MlJ9AsNwRf3/NMN/gDPKtoBUJGtO3BjEKrl/QDrEOObRdsbixrb3h6vmOGK1t4fL0Kl
7zvdmf3FDBmNVYyCSDxwziFX8pI3J0eBhA2IssEv5xGz/UOp+quuvfdTqGNt+haI3x52en2vpnQI
dgfun/IPrBTBeAODNSe+D9uQW0Lkxjn7OXFaD6hcDY/4LGMGpPhk1HMa+7DBQEx93Wr070dRdRPt
pB2BcUQp7uHu1wjJ8in6Xu3lvK+Djib+B7KaWB3G9LWiKABK21k/o4FzgtF4/KtcTbqanx2ovjk+
QAw9RkZRWtUpA6JZ9AQIF0Z7UiYKrrKM+BLZ4oNN4F3xlu2PFgirxJgmRe5tA9ED1O1GCm09us5r
3K702oDn1VyQJjyLjdNMPs2zYJ0rCMpWrg3bZXkQTgCXnYOCdGGEt8YYLt4DgroGKgjoboaI6bk0
HRBSKDZa5KJD/eGSanP/o+/5hFhwZA8M5INl0eyZpbZbKZl7TsXprfFMKe+8zf7CU8rAlGqrtEyf
ngQqDZMQtp/WCVemsB9aFSyWb9cXKX0vDMLZfqVQ9y7ictxBrFsKw872FLs/VbxoopDoljgO610o
VOAjKgV8uIoGyHf/uE62C5HQPOdrvv7qJl1K2KbvgETtlYyg48GtNDLJwWGLOyGmIrLtWL3hk7bD
uF+BowLKLOqPmgTJMi0bfM4aOGt4EfDocSztacpi6G+qUuJX6ARroW1194OGZvF+7Tkt8e/hJWnD
Z7MDHKyAkKh+Vp3+/eayK8Tax7JqYu/559Gwv7W5hC3k8FvvXBS9sWQZiQuZ4L9VhKkcXlXg10s+
0E5RE+nAQboC4RrT/OM7pyK87B03eB/DHtP0YcEV3gcATqQJ690ef1Ra1tw08fSvzvcYSHKvVAmr
o2CfNkERR/Ko6OlGjI6odmYK9aqoF1L6GwJambfw8tCJbSPgYmhWPyOJb3JoiSrQyyJrlK3T5vyq
DH9fsZTG/jiuzil3yNIuup04I1crSlKCDPXrqAT5xYt3TdL06AsRz+jdw0Q01xtoiWjUPC2JGhDA
jHfcecQ0pY0VNsyxmeQ+k822RVTPvLq4lGlQ6/V+PZbih0JK7zzqsFM/G0T/BDgiRCbPvwoYbvz5
Km1ibpo//ARfyKbxSL1QwLo4VEKZu/pHSiuI/OqPTZcPoWiEcNjit5ZmFvELo7qY6GKJ+BtAIYF8
ZTPKiSYTw/4a8BRrL09X7b7/2d/siKhgEcwVWfCcdIsZuhHazJ0oPdbaiMmZgKdHYj4EV6MSirzr
FySbkHHlbO2BhJExLYmZlhfzbfQJMCSbSbzpJppDKf95t8P9InVGZHvwOsMDnklanGPHkBZB9wE4
jPRDXm0cqSA3RNL7edrOFFjVHOga5O14+lvb/9RUlDcPFhB854NEnELKSe3C2mIGVWMui9Gyg09M
NNSAAMmrouPxRX0+Mplm+JFgNO9wyUfmqoNyN0Wfx7cBomS8nrIhAkb/0MB+hLaOK0V41ubjPQbN
iplOuiEedUo1YjjfYftTOvm2Xqv9e1NKkyvCBYfWdDpqNVsVN3zkm9QT9AmrmzVbY1AztxUnxjIA
pVT2SdOrWKlCA5k+IpCwKetG07oyl5hkT9JtB5PvoJ7AavPYfBSPbMlAwGOKPv1AzhYQ3Z69yVY4
wQ/QVduJpsnibsM3A0mct4GFVtMEOD43DS0zYOI/Va99Dmm0oMBKUvSJ7AJIoiV7XV4/htTyfFas
SZfPZ0ASHmytkrSQKYdHuK9k0+b4lyI43KFKy6rRO6haVG2AQmm7+FJWegK4gVI1KIAmasGBeGJf
lF4h9pwUqzP5pcI8M6M89WHw3Kh8BC5d6uSEhzZdwG9/BjXAsJLnya5HUXYg975au6aoI8WsZ9v8
L/6XyY7yookd+u1SNsPORFwJZ5oBX89+xsRPHxQmMFoMeyKZWRlHdrcptOruwgUt4tCaNo+HdJMZ
bimhCbER926yuBu/CqaP9QSpJjtZ9E9JSDNgSOFWkl4aWKpOEci6QNTmG24DQR3ADm7irQ9c5czW
kSUdlSbSc7aydUWHglAzRZ1J0O/ABYdH9ezxWNyuRV4knUeZSWClud8VjfUJalpOUzRkFuJkbz6H
n2yKiR1mkq9MWpgDbRQP0jtARPmjpfk3MapRjhNIKeGnqHm303QV0jI3lCO9Iy7PqNCuOGfT4/c9
02EI04H4oa2C8XyKVNjdcx8xyTYbPSlQy50rM12VdvS+wUhEjY6l2oDDCO5cgvAZ/yF44aBdQX9p
tTKW0OXD+CPjtBkJbTEc1sPXNNn7vf0PaQ2fiWzn/GhDHyNirdiOPXZSuUccjCf9VWfMvF/Cp1Us
jbFw7rjIwfWiKiXK+tnfyGwHlwMBHmjhsaLfHNaTRTgswn9hU2p2YBCupKe6l7xg/tJUHyAlx2ht
lZ/sPO96vPPenfrBLZ5e18H5GkIaDDJYwKB1vBaIKcUFb00AeKuLogBPZIT75m4+XbxnRROdt/dF
e9JJyvgWvMOHUewM2Wvt62y7F+Hplei3s0VaAuX10vqB43hq9FQ4gT0SuJ1Wdz6XdzhCKVgM4cyY
QbzhZsqhgwIUJEKepW9dNR20dnXLdoxTmv3V+9cQpcJVnrITMnJ3yGgleleYqCwFXm8IVlQfEYFy
T+zHGvDawuXCJet+VbOUapUcR35468ulFmU8QOpRbQ8hf2CUg4smvlhxiZjkIZecX5l5YtzMn4tV
7Up9umwKvRpObHVb4Ukh5D8uX3grFsxPYIepmJA4PmqGmQixCB4Tu/sGuqCweF1U9DxZNGShznZm
giVNXEQ93wztYsJI53bZSyecWmvwsX5b36bKXi/y4xqaNmPYcF7rnEa6oUjblS3Jzs1BTh7t27Pi
F/MGoKA04yVdwAbhSbtaSaPGrspbgQlrj/93rRsTX4giTScZakOiPjJaZwhx8rzvzlIUy2FOOWUw
FK0P0LkuviUyzNjO4L16a2WUreWZ3Tv2K0GXcMp9wq5ph3vO/qQRO8LxSZNDsHQvVUrBBXjRHEdC
UyEVnMDTmR9IQIU7hSYxPwHTn3rxOUYchMMkmrO7nIl0ZiSrTCF2+IlklB74oJpZFj/pPMynwlXc
Xm3J86AraTUMx27kjZcx+vx6tcud3mQ5hVNb13mqgBj/cKg9KJ0EF642bI5K9MwmqebG3DDhFQI/
VVqc4FiAK888h+S2+9i3ybZMdDZd+yd++v3Xj4CDD808tqE7OQLvJIuYtp0pM4YTAKHhCZKaJuRQ
hzicKLQw+g5sadZprqH1f+/uWhMwERdD8rYZB4kvhOVO2KC8AhyLlGEbuBsV2N6W2NE+1emcowgW
/kqlSOPV2VFQFhbLO6BGu3KFLLvrOj4YWvDrK297g/pq+w4eecGdNkDm3CAjKcrbBqroo8MYWy1z
tL2UkFis9Os1JA6Gb2Zv6qd0wQVFl9u/Ku2hENQ5vCYJB1w2O0hdTGznoe97YM61eM/0SWad3NWd
yIRofMQ76P7+1ARTR7N5d9WIpWABYc83VYeyWNsfxOfB/7nZG3kga/vUdQc8mt5TToywrxLNr/Yl
SrfWOkj2nR2ZcCpqHKyUbrhh2vPctyTMOdVS3kAzCIIr4zimp5tbgupL0mfNSUsNQq4EbjDPMxQZ
2Pac0lACGv1sEVK9zxCR/d2l2MImDwrQh7FiLuP+d3QTfVIbqBw7nVMb7RLm/yJcOTNTFHNgKEEh
Nru5Ghgq+4+BBf6fFXL+c2CcXIHYcMufY6cAUwetrYy3APXBlcx4y0OhsrvUsNoUVGZqMa9MGU1w
maNcWiD/H5zJrD2t1hRwOVYItPFqybhYMhUz3TwRXnuVKOk17s9O+weUGgR+9MBieqW5PNh2KOe8
kipVo8/gRWbQRy+lFhuW0Q9dTRLSuB1W9rSJ3lELKWlD3d+QgWlDvBguo13TY76oJcqnCnxsv+4o
g0+MpolZ+x1eGrYFDPyyXUy/Ka7N/8J2jAhJmVoHFrZ2lsVM1FkqIHhaCeaGjPTflsfjaCPX6EJu
c5ZMGTzv9UAeWKI9fNhUocyJ1Yn9lHuiJtG8TJJ17eZTUmDlzYwacuA9f390ja0xhJvCOxZ0LL0P
ch0O02YUtX1OtxVri1vRqyZoRveacXeE84cXHWqSQfVlY1qa+6MqOAOd4hl7138QxTTqyO9VMq8E
+uRgbgmruBn67wzOJENcKuiQnl/jIaD+55GyWxWVWP0eyCtrYkARsSdm7JHdNdeeOndGbds4yA2I
B09/FRqxtfvPaN6yeEaetGuhmMq+O5g/gM//eBKjk9CcIHtWDAiaIwFb2Ktl9Kjj41Aq9yMuNXu0
RGYYQuGrMteUmVCP2a+9FDpenYJIolrtSiBUfGMwHndJgW6gIRtFyD5wPb8iG3F06OgC6zBGVm5M
1gjsR6AeWrOGoe3kwDgbzSicZmCZ8lfQgsKTHG4QaGB7HHIlYogKoYlk27ZpViX1pZojZppKN4+X
gjx5E8FbQaOhdhhHVg9pSbZPFgl/1YLYEqT0jmHKwoG/MiOkoJHj5AxLOg5LM1HSMDPSAWLEC9nA
g7C2UY03r4bfjsUTzcHx5PFdnCHmrGcYenmjl5Y1E6oZUh0/VlHaiBHgLm3dG0P9mD8So56Q8poB
FOSSUlfBRbBOb8pZkP5TZ47eJbQTl/1MV98jJ0mfay7gCQErKYX/8G9cIzi13DXBHBpKv7Yg3FuY
XzglIRVRN7RFc274j6v65/vTLCgl21Nb1YHi5lA+LBfUM7Ot3IYXkBu//34PSrNQLbU7jx2C/p3S
Cel3psUSYVkaHNWKMCu11abQzcxzyfFpCqVPS1O9YmKGaJ/T+/a6GMDdUNOffqOn3MU7Q3uAKofI
cEdQuXwnuM/1xIQ985ejTh53flbpm2sztWxvAZyMtIhbSfBQNcFv9O32QQ6zh1aHv9HLuc4nizNU
LoDv3y+KfGS8MRki94KLiHg0qSAf/7iQkLMu23x1J0y2XGbTmaQUc2PW+yILCSciVH4O+S2rdpu4
GHGBMIHE8vTGyX6rioeLrc1RJFCf0fqDwjQE4zdiigoTdiSVjuoHrXmIaFJlc5jSdSJlPazfDJGX
cLDLa1GFmswdbMIhIymA4QI9bd1kYPM0FAAcl9IzoDlXNvMKIeD1mVx2zBGdzdSLeUzvJNqQvbVI
3No4+Kn0/XIhCHRTCQG88zmcpdtQCtpU2yAyE3AkBXMET//L8XEzgOleszfROKcjG8NbJdDPzOxX
kcnHSBR/iKtDK8eOwSwwzJLX2MVEX2+klPb0rqAYIbDdnzPI6rtw4CCgw2qHe4W0ocARnLmGFWwJ
ltLvsDAvOOpqrxse75iZH838d8Ao/4ZPk6vVo/vlSCTee+XAycpAQ96bPfUXi0gms/1mrpdrMPRt
LstGnK9q9+EK/sPNlOcYs6AlBq4aufqdzbhrzDc6GbWBg/QpwVEE6D37xklPc8QoG2MlhhGyUGdg
RlIzwR0Drvnkpug884VCtn969C2JKcX9p1FNZSjO5rtThpaGDQ13OyvPCU425CmN3xQZt4jAwzbp
S+H9Kze8+5QTm/0j3kqO4U7+aTpYA5Dt5c32qela0J+4zlsFdsywlH4YeBjvNGMIYamxo22wKPzh
LEbiP9UPxLBQMz96NGcRgAMM8+cS3D7JfI+CTW3yQG8xRJ90hJfM4+WVaLOFEjavp32EwEujkK7c
oiOW0C4beY9JyW3vPx3GiKoHHEDOROZqR8JrMEEdI4g7W/7PkZ2ViKSj+Xc8gZN5dDzNEkO4rwPM
Pkh5YngbI3mchYDM4cElJkYCKN01SmaHqy++SYJgDXtPRWNH9WbNJb4MeeWuxYNpfhcPC+hsOSIF
bjHYepURKz26Ou6oP+X2OAU33AVQ1HOCayTxDBv5CUERJ2bUr9mLs4jXbEHVnhusWJweUBuYWxYR
pWYY6eV3HpRQhAPRTNvy/7SpGFBiSSfNF4f+DWM1WSu/bC9qDaiCMKIVSTvV4B4P96Bcb3l0HSgK
0TtB+KvduwXFrid5oIdz5fZ+EgdH3IJRy92NBL0ugTjLkNlQYJ01T5Ay3OYRbi+8dq+Fgb1ZOAxV
FisowIV+TXOA7XvErNnpSFSDI8etRi2LNuNsPyHol7TOI0wBh3rQfYLc2KUgfj7C64PLNvoGGAkX
8dJJSkAltirDT2w+WR3nL5yX8v4xxstP57tEasY6GQalzKrQp7SJPzy/H3tXZkOLRdr/PaufuXOQ
Vyn4uVbOurhX4FKdQrF/Oyoj+bpoE/dBFBPWYeB74RDYrbXmU0q9tbysS4OV4MRO6XXzaAEemncT
jXv1ZbcctiCgpS4XYyTL5suLjPpFaoOrLSSkJ+7mAZdL2+fBTelDAPbUnUCI8pDsO3rDJnsft6Q4
c+Ltn97kuP2oOgukNx58UO3O4M4r5T22Ud4mkFNk6vRTzld2gXsP9neQmnlMd8A0RFoKEmxylx/a
DKB6Rmou4FN2X1jwoyI79ZvupssR7OLbS4eHnEgeNSbG7daAifeurf5TAwcjl0OqRzDgwL8zmZnu
4zyrIr7t9hKkkQi1sDLpwk/L2fl2BAiILXV5RdUnbtfUEH6wIPEV5M/CULIiDMjz+BoCm9M+8S/w
BI0BNAHA2orZPa9KnWlWFU/SposZTvBxBDR9pIBb/mS8cln9UZ59yt6QAidjayI9LlrLBJTwVlwX
y/IBPb5abWCzAih9mTFRn8QVUP5CI8DapWDoYJx0tEJmBlVaQ1pfjnV8Q2p3BzQ/Q/EHvstosQ/Z
4YwdHkm8hMW7m8IdEe7ra8KGKvUgpgvWS5YMYkd8pGh61kP7UpiWj7kZeOkt7MmXIgwah+FuSYBq
oxZD9x3bTrHSTvt2mDXcYGcqnNojukmxv6Mbsw+g4yzJlLCnQZwMojUWgB/EySCU+F83RU96n2o6
ynFxY0lKMldu4USFBA9zPUqJwag1wdnvLi3V+vdAq++vaNugt4GRuwfIw0Wz5Kj8lKbJUvp5noP/
ZNpIe/NRlkMbD31Fw4ViVPtfJu8cPhLHgrhVcdyaFXDGkOm9y3ObmJxaEQlKGsLcC2EoMLs/zB06
DGlKSP9t5GtuulWpblMT4htnOOzWvtmpyvrIVffW1he1w2IGJz2WbJIGrYQa3191CykkznWZhvZL
LC/8Qfwm58LvLAKOjlmfWqgJOW1KHsMOrEi1q59zUv58pf5/dyBVuFsuDkMfN8Ha6f9fS1KukO3S
PL/6NqlwzsKjet0izmWlBvkL4NOnAe/+0uc0VYLKK29vbPsCdv/YG7c0SELZBejLBBLoS2e6gs4W
LjIabxUZrPomTUIlUJoVvgzCp4LEgAZnDvGOKPNQzGiEsbv6esDZWNcSlXUoFdBk9xBMRY4EDb8i
+kzdDCgWvgOJ9eCD6n2pq6R94VA3yzAv/4fY6KLvp/EJErZss+d1VHyPM8Hzy4RCFBGIq9ikwtNv
K9yOCNXsKWZO4ox0jMkee6WtWUlPkGTv1XT2uJVcDKhSNyDzBmOozVFNU2HL7yjrUYpGRH2GlPdZ
3tmSiJZmu4oQVh7Y9BVbRH1lFzdUT5HdtFazFh19QkWwsWjcEPXgZ3/HKbmqKZ6WkjIMURHtHDjD
M/3eG+K4QBLKQk5GCkxsQm+1jHDJSQgUBSxTNHFbGtzZTzdK2D9bi3ruFqaOCbwax/mojSI+sM6k
EFjak71jMo9yV0ZPao8NOYjElD7wS8q0q5miIFpyRBm5wf63G9kxlWR9fg4sykS8xBcUYF1jFjTb
4zSWkMOI46daxZybjdr2LA8eRJQOn2D1K0e9gr2zL91VByoB6pbGziZmRa0htPUrlC/Ug0vGEi0u
5SJrTrVKg8V26K+R+hOsLn4BqkGGfYLOH6Y72WFgEDkNXHshtoTAjLGhSoqnzV2byFnCQAd7ZYKI
MmgVlleRLgjIy67ao+taR5uPoGU9oh0fElyFVn44+rCSue6wRNTMUh5boOe6NYnx5j/5pLeIfu5p
/aoZt2u+Hn/sRm7PdNzw2QeSSvZhPWiqtVCZ42aJKbwRwbViNkxiR5fy00OD8hHTLxffkZqMSdFQ
+p0tZVqGDNtu436o4kccZgwWw0yZY9cf+/GkvtTEU9iaGV14n32W9IsiTcHMvtxvcpmd7MbE8d5M
nSYvjkqJLDOWCWiydEVjvVIVpz3XXr187IqHsM/v5qggv0IhA3ulCMzjKba3ElTFXyXVtcjdV8eC
3B/ntj/N5YhzrtD84ajjMaIaI7ynRo1wYta2wnYEhuzxcOD1SXkF1Tad6gh9XKUyQrPtShGvTWYI
ydtxAZTj5jINGGU+Zg+5gg5E32u5u9v5UaQQzWC8LeZhnBYWZo9SoP/Ne229DVOkFPUovtB7A9bb
xc38t7Td82G0M/zwF15YhWPmDidZ/yMcuWQOiTyu1SWrBNa5KsPghKsnv8oO6QJ9CVZMm7BAzJYz
7JBEJOjKD0LEc0MuFjrejiUFGGSkkrDyRX/RR5fMM1k0R6YpQZ74HMR4cVTqRgEBkfkveVZTSdNd
Kg0c5NDUC4J+x/IKU/Q+RWoaL5KIVf0wjLdUxNZlE1shX10Njrgl8qXvMYZ5UYS7D16OHC8thJ23
md/GfdbWSxKnppso6uCqrl+SoZvM9CK4sdIEoCLLie94q4bYdq89B7EI68OfuZtVPEOHsU5hC2WV
/yEciwtQzOJK86tdVSTAOHZUSEkshJs+xAPj82m/G26vJ1y3HDpAu/ZWAftI0B1zNrmPjiRspPEG
f5eh9wFl4EQMfQgZbt5k/PJ8lbgC8AwIOvIVH4LNqA9irDzqvtXedsUufDxcM1CcESPiDRprBrGB
a03DMwNLCFF58eKtY8u8NeSUD0PwugGXwEViwa9ldYynonQJJSFDK7s8g0zUkeCUumwzzo+bkIr2
Xca0Ouf1QTaBCGsxh2q5zy4lVoWrkxu7iNFeeY9HdcxJi+2YD3l45th4H5XxwE8Fjy3DZbbR37vG
0wj6/iYrUJVGfVnBzJizJrurbdQS6uhMJjXtTQ9CP5hKto1fK0Dwi9CcdDJBsNZteRxDwkBB3S9G
Q6dBmD5jrYip4sRiC1FUQvQowSqxGRD2RO7hftJLhoJyKYuCludJsROwbnBt2aFYPAlCzMDmGqxn
bLlYUM3LtSjaUx6Yg9bReWJOZRlcxJ1SWYnhVdgyuNYLTU3fSvopj0o79mkRF/oMGdEhrda3uGpQ
kxh0NEtwsJxyte9kf9nKb20xynQndfNvAq39e2HqS6flZ7fnvilTIo0t3PxpusWocLSFTtBCJqED
bAA+UVxlevLhgmIjk8H5PheEXifnanR6c9tFFb5QkGmS4NsWuaLySiSxOFUDxTKXbeoIhMrwGdnD
E/fQCQ0p5SWOO04dTZLGx8c++X/3m8c01USUBVrjkLCEBFfP900HJYu5g5yvXtx9aNQ8Ski00vGy
2pEgbJHcJp/AXn6E1N/x76uwjThlYd317+lsNzJCZVxzndUhJ7xgEMOlMdbCDmD21skCcCQYVaqS
kHgXDnOTaAKg41klSPQ0/eGSEzTDjzwJTVSukvei56TodB0G2UacJ6UutKTWV2FMpfFLWKSlYmB5
tXneH6bmc67DBnsdqU05fSToz+FKvJB3t9xLNJ6T7oanSp9RQaPBPS+qTR3h8JLdHGtR44fz092p
sugqZ6xSxN6VFRcRpjdloLIW+JGF6CWPDOaawl7ptZQxMLp7PkKWinV7i2L9qyqTqboCK0k3WzRu
18IYaOw1RjaukY+fazHimw36obbLsLjYVVF9kW0fjRsQzozL9vPWzZZTYEC9URIGOea97I1JcL2y
iQLBVmd0p/f+TRGWul3U+5m82JDGMpLVn52OGP0W3ocGqRRGxPJtwM1+bxlWSP7mbHxmPa4m24U3
kXnbrQ/9gpCvzRk++FqyU8KkKvb7xmFybnMDYEn/s6K2KpfakC9q0NZJATQWJdqGr5aNnf5LODpU
vQiSIDmhWL6Bd3QUAjImowqEbMPZy0aqkjhCaqTkO9NahLylXASWtX719bYwLZMR7E8BjLWBFnNy
mmYNFe5L+H1QusjEVEIBNDGugFRtSqQyJk50O7VdDtjLic7tnBUA1THmUsmx1PMXhpe4jTU3qOuT
tJBOj5VHK76CVW7t78rf9EUsFbBP6MSiCz2FcuLcpvXwi7AXVETBzHpj46E4XXUR0Af+gDc7tcEp
ga9JllMcl7JmQD2iVrXZ2S0phgvROxOVp7p9CRX7212QE9l15iCs4CqmIm77aJnKn6kq7w7Sr4CZ
JAAtRXqsOancxr5zm/EC1ojvVdm01YJ/6/knYl6K1S+NsAiCB2l4CyVKLpnoSuvY6XGWC8uGYPEV
5tp8RCJNvcbgFsyYy4slpJby9e+qfXMgTE4wAfSmtxnZTCILsVvKR0Trq5ZN/CfceyksWKmHuMZJ
TA7kjh+NH2mizq23Z25UA0L0JOt+6PvvxMFS2SnKw5F/sFegW+AlE0Jbn0SDo0nV0Vbk3HvA9K13
Gyy80TjmvoZWNFAJ3AjC63ki+BEK3GRlY7gqvZ9QJ0SO3ExL2Za3UdCboPGCrCVMNdtxWJu5yt4L
ElnV8ahd0Oj5WHOKqqK4e+Tv9Q6RNzkE4wbNJUBSBDyponE7fNxSVcuun9hpDovGTW92oi7sQ6kl
LSwWgAt7/1AfJ1IRc9tJXlKBN6fDdr0amlWYbuSthEtbZaqoSrpFavhrfwO0QkcC31A1ZTmUq+KL
5CaNa8EBp0wGHNKjlzG1D4yVX7ovr1vCTFiN+FRm2K/lAibJUKxjgoXIEtKdb8Uom8UykHohu834
92sygLLPA77lpcXJtdo5RyrNHra5cuv85s7BclUf4Cxq6rPJqNdbe0FfHJky0aic9tMceApBM8dK
jtA5d1vTCPfNzBUJosU576EIjWLopiuDGiQfP80k/dKWbw3j3s0jZ5EvOMyQ3P84FJgJz56liCz1
D6Y1E572QmWgEXy1TY1DOaC6Myq3SiRVYchwvgR2RRDJMJs2gY9B0JLXMDgQiVjo5SKWCR6XrgQI
D55PSxba3rFdrizeiEoMT1cajOk3SsKINiNhUQyl6hIE3Lwyv8s+1FOk0unwqdu79+Y7pedM+orZ
burmB3OJoC8YdPcyoOij/0Pm7DHRTtTu9RojonAXVRz/EVb4mDdNNekgtFy9/1sUJoJqaeMk2lk9
ZW/MZMeuqkhtwkc2FLPajDiB9DzTSGi6nbc5ZV83BK/HyNecKg2qUYnWXyJPFNJ9VnZu4hM+Pove
XkeT+aoIdqnoFu+bzYP82DUdaGYG5ba0kblheErLWjj/INZnW1Qtbm2wzUly8G3g2jmMn1Y3faY1
WORKUdb50z2nFAjfTdkLxofiivBqIpbXNBbuFq6gWX39gvHH8rFnw4v3FJR+ynpXQv+08Rsnb0PU
640Y0v+s35VYotX9RFYGoC8IQTYK0GWpI9ROzexOYV3fAoEjODldOCIDuWavjVE9GFapEaL1xv/m
yC83izngvHc/VgbJgbL9oWwnET9lxX60rOy6g1BnBBgD3rX0349PfHNyKNeWp0zcqlmGXssxLP7n
HoKsjzAJXiNEWhc6la05kJPzhYYPD7nADjq71AJY/5p5hitJgx5subjpo6XYhobrvlIkoPehntbU
iv/Ad0h3ccL70JNhjSoRjDYpKPd2HdnXzvozfaOtYi98riP53bvne7OKJ4ykVPdbYNPmPKgn93NR
d/kkmW8xuZE35I7sqDtadH6HHsDbxJuBtx3xarS5SZ71+DxsO2+RtSUslovd893/qJ0JbwI7iNx3
v+WtdDsyras0ct/68bRx201m88M8CuoIp+LaP1Bk2vL6QOaq2jumclKPhQMxwSBZWOtOa/74cnZO
GXtHcbj449C5OvltbETdwFfvQHDg52+IZhLsUYZ9FUCOp/hUPeldfg+EKqEa8lHpYCgxuZx/MuUf
OTCaRJyNIeTQrExspbndY6HZZpOLJZNUXSL/0KUV0SEeSy6rIkWU/B5WC4AfG9ToaZbG8dU8Q4Ej
o6zAzfXtwCPkbL+a1AFwZBVQCBdiNIPDcOerydlKahEmOkf+fW+Ov5OXWTdAsFN0zeI7HbSe45SH
AK05mgCsZOUPJkMcE1F0P+om+phPJ7r4d9JrKPWuvm0cRa1cRwv02iXwpDNUsHE0/XcSVQQ2/JoT
rCbDww+zoNC+XZxPZ4wp0owFQS6fDVDC+lIVWvH70wpFf//jadRLpgu8MAJTKGQZUpDYTPcqlqER
DTRJ0FC5Dz0JcRR9KWZ9GNSMkl1h7jtXlExPO6PeuALn5m6mL+Yq4iW4wKMdvCVjsA8VJ/kkPaC2
l6IyiC3J9350nk6tqBNNhhrujbSz4Sq4ndMGnqueV8NPh0XZpxANPRPrxoV6PNFTm8cNJM+qgFWI
J83BC6TNoftJvNPMWQunHtKlXXfBfeoaXMI/F1PrwioyxUorr6aJl4aDjFZaEFQDHd9I8+2JsGeZ
lTBvJN94VgwngqTSqEXwUOOTecSfJGG4CCXdeHeykSlD9pT7/ohYDYVZhO4f58HPvj0eULdOwVbe
7UzZD9lGIrvX0J6x1ixhSuun68QjRQTPgRx9B5mELgOnflTI5yXP+XtETcvluRv7OqT/MD8wGuUo
YVbhPkgzIsHGUrIXj6FE++OyZ5zo+24vxv0fLj++51xTITDhQwSWrqUHq4mT8jWr2+3KQIDt0PuN
nzwTHZV52MgrzQ35yTviTFAptMwgn3KhnOtCr8Ng7AqXVr+LcZ3BdIP9UzVlAO0rdKJzCRI+ArAS
2ie03f+PxdCcHUvQv05CRT9YH2CMxvRSuOjLnappfnTic5ZyHmMQB+LyMzTh/paXTpmly3tTsbhT
7zleY5krFL9nRf+fCa37I9pNwKGysTj6B8fCpUWXE6/hp4EWp365HyNHm9sJvZAEV/wzCs8WDy7p
VmrWRgtLS5lNDnXPs/rHDbUW/5UnAUwSF+ItnaHVwjMMweFA6Bm0esjwUS7FLCVcutH85pGvW+fA
M88T4b38H38IreZxM3GPNR3mRjtzT/QbvHl6uMVufUUZ9Arm89f6ZVNidzxaWAyYyufkvXsVfqb/
llfkUcAabOWLCKtcQbLDDsSER5nLXSLx+I/OhU2Qav4QdVdZ5jCT9CLzocrpyS1wR/OedNcmp27E
5kHTWR35c6YHNhQfzbmpFCP56qSMTPr6QSpiuDyw3umyUsk0VLSKtMWZhrCXAINupF94y53Dlvnx
QMuNmKPpV2cMe4rLKFYSkFe0imQsG0J1T3IE3lqMKfB220S30U9tJOMMpgEBBEIC4uEchXjnhP68
VzwS33RnrZ+9E9ClXB0Ziu0j2Q2e1l8FcOZZ7SsRQATbqILvsY0SyLBr3rCAZ2hlzkDbpZ3niwOH
72jcRaEKfio4XvieslGvfv0bD3SHV8+O5RdkNieiBg30U65XH8r42iecRYeMYAau+UBYJ00eaZGq
FYRS3QeteXyeyGQDqCWtzpepVsGTuou7Dj5UwCVSfEfjdEB9TONKNgp04rUJVl4cym7HYeHrU9Zr
9Ya7f2knhctcMLiaB0iggth0lHDrkJcATNc83M96h1lbn0o849JzABk3XcQmC3wtUV0Cw9L7RAi3
UYVGsiTCy7PL29Ls8aY0SkaHFELsNTtm283uOKaGsRy4nUC/xuDetBEFvQZCDndBWoYF0NB0wNPx
73mFGNA585vDLStiGmtz5n6pvylgeHoUhwAdk+/B6Q1EpWkA1JRHjnhqhMaMFYybQfn/kVkZW+w7
lNezpsXkfFG+sOpStokvc6CunEoImnJ+AJ7HANlb4xvItoAwRIKKCnNLezvOCZjEokv2fd/8IjfN
sAcYPZhW+V/4lBrJIzbnh/UzgfjJNoMm7i7U/cVDGT81j8ni4Gb6hjFsEwqR2txVkLB+ELenCZsE
RFjIcGZTCWKl752pz2io6KdvksT2/SWdD3pr1GuvPG92fa6VTJ4mseaMve8oiclc5pG+1o7chAmf
Ci1cdnPecI2OeTISJsV0qo5V40TGlnjtD4Xy3Xxh8Cv6xmdhMVtUC+iNWOv4OjSOxRdqm5jm3/YW
IpsVUPd8xcjZgIEvV1ZNMLif6fPMV9kVqPhyJSguSbFUpBgSk3CLGIBjEcYvuH8C97zx4Pmtk+t8
/26RViln2R7Q63l+benU7KwcMWpCcx/C1vNajPFT5c/3rUxcZBzwaEIYDfcToqLLwQcT8gLlmYOI
LRkQN2kv4BVhcYxYnkb7hkOFYeKNwMePP0uLV4AhMK7sr5k07XN1R0nQIq36wYjJKoMrO5eMH08Q
2whewX/zVs7nVoWKy8rmgmRlZ8E1YLNuG9tzlwlhAU5+ehk/z6AG7u34BSauuE37MSdQvv/oDOPT
oGBxBw2WazIkGiEn8WYitWGTwiHTrxoBAyxo7GztYs/BA8q6KI3cyZ3oDXyOO2wl7fbb4bP/RRWh
u7SU2NeZuJBAmVIH8ymQxVynQf7hNz4XZamXl3aKAd5nahLRg6++vozXPBlM/v79gV0E1XiUdlP0
5suHHbMAxfwXg11j81g44qxe/d76FZy+e0RjVbZUZQMDSxX+H9zxTYY4LM/rRXC0oI64C+Gpo+QH
mY5jAwtVsSBdPrlGJ/ONY3SVkdyDBcO4ySbxayr4otzIO8Y9zlgEOopc2BjDJ5mqMEn/FJ15OgTL
rcWrY0PBvnOIFdI09BTodMCQtFsRhh3N1AiNvHQg7/uKhEOGKYzI+JHt0su6dJlfuP+PcwZGG0nb
H/7nwLZJtKeSMqVShkrLmjLCO9nf8HifdHAIWbrX+eJTj6VQ32yyRjVgnTs1SC4R88sowh1WlwvO
uwW/V/DJRHytDkCAf5fQvqhecwyzVLG4b3QrcszNcAGYF+EZlnrbC3327fvZt+EkIvvkymkUddaI
YRvtw+vWY3ChEZ6kwKMjH0TjeYZ9BsiqMUKDzbGWiqjbEFXAZ71QumOUpVrnB2b5NqAjlq7GFK7e
cqYoFjy1ka4uJLhIh/K0JMn4FTCaWU7368Q5yhb47b+xrklF97XlFmOWNXpSHTEiVc3h2Q3bCzat
QuxPTblgQx4DDlcb0tcfNWsyg5foIUH3E07uODrtAZRlW/rleNjtJwAy88enPNbpVHYXY581A9Sm
z7sDWlCzfjUrs1BBtBq8Zvj+Z9aSnM2pAbGtikipk8w5JNN4Pj+O+IWrwCpqyeWvP0PoGDhE/GJh
WsU/6AkUZj0rIFD5FXGrV4DtU8ilvUgQ4LKXU1jokHlvL7xEmdmwe2gcQQaStelxyjlY81L4sujD
JMyZ+NvlXEChhWFBIirV5lqRRecOjyzx69KyP3E0PPAP5QgSh8fE+FGlwaQlimlK7Fx/OHQazEKE
Z1G+WEq1UlbaWErzBEJCZmYpAxPbO1oeiOj2pj1WUvaI5d1slnx/AZi8wCiW/IeBTWmwsx235CHK
GdLhlp/NSgplx4s+R5hy1K5W9WFyIyO2NwydY7JvlvHfuzHUYxKoXfiphJWN0kj82FF9vfM1l1fR
PtcF9lintF+qwCb1qU7tSssklSDjLlYb8r1aMzp7K9r1/KJnVivuUyEutP6kY4970bVOS5Rr0HKJ
Dcg/pa2ej8N83OBaPR4qOabsfHYYrmAeHe6qV0H00PfyyVlYyO2otka6CAv96dWZr/in/FNN3WVi
jrwPJKQYKHSwhIkDf2W/NI2dvt0Ix7bAE4Yz80jHeQFL/pXe0T75K9osRqIfS9t7wts9yNCaC1Ei
8Vz9qHDDJfWb5WpuKNQOQ0rgDN/rwnDNVs8rBmYvLd4LCjwqwAuMAOGu2ao0/DEiggLczRnXSQHM
usAuV/bVPWy1bHObVUSmdPi+wjfKi5OahtnseWJFWXi5Y8AOmpwZlg2f0OI8JBWszED2VvbpPuZG
5Oiw+CjPvGjyd7eFQ9+hMXvbJW1erKz6oGgarjzr/Dapf8rudFo/8UVKxC0kSBFDaj0nHVulVQKT
zakPqugkoQOFoIuvBpTIvMi4+qvLG8L8yXTKWe1R4/r/bnwzeofDMTjtqwyqbaAQL/8RzbEMuM0w
nexCAZh3lyeLB4IgMzyTVMRl9J8ly0EAJ3aNc9nUepC1VS5xNoBMdBYzmBHUxzAuC1Gq5cwIM7KU
FCYWNDIrneMglPNH6RICsE2oEHd3tpbI5en9p3WuJEYKUddbBA479VsEEv+1leduVi+gEVpCzvnx
M25PiN6Otam7cp2Rf4Gcthlx12oz0qhVu+HJWR5qLTse/8O2BtfSj42Cek9M9R9gDXQbdBaLC4dp
JcNl7UbWkgPlRr/FkOlGWVOvos/dwu/6P8q2mINTkfyAv/MCgaePsL1+Nwl2fylFEBukwCkLIpYv
1qjEmYqyXNPkiCw0q52xfyNtGATm2O/UCX8Km1NGTfcH5VWtnpfiQIMBJl2/W968CSiVo9FRmnrv
asuyiuXSIoYkTxhPRTH5ZqXUxsUvM77qI/CdukJMCkdGJTQsrnm7qbwa6CfEcOyJvYxxWJZblSV+
5A70pq74QDTn9BPCg2TMihamByEoJTwFW44bQ54xWEAYeyrd77ctvux9aOMZGZOqLSAegArRtjx/
JrEvcmSPuPu1f8lroiyIbybf2rWBf5nAmbI1IjgxTzC7wDXh2V4dpLR9OsyBWL6joDaTtcqtGaK4
vj55EdvXmf30GBgsFDuVdxeoTuhCpXRzPZC0/uhrYVj718S9UAMWwzNqOfcrL84JUjkPKEP3s+OT
c+dp5T9ebP6BaXWQD6uAWA/3dvdXXHm339ifmUiCcExNmRIGfTa1xo0J6Sa81MqRGopAR9WCSWYt
jTA5nQg3h0FsbV+B8me/NqyD5lDwP/RcKBO9qxQ6wrvUADlmkKfBMy8o0isf+bFKcGfbfXnYAmpX
geTjuGuoy7P7xKTAKkw7cLMx1K0J7dSQgcUwFy2cAo2/3abFn7tQT6Npnszh7HeHDqHn6Z9g1VV6
AJQ6z0K8dNDdS33PIkUn6Xoyq7ihq5PrhSk7npo687ZJs/bkmxqex+hPvYO0SfryspRdUKHCnFZN
kLWXNCOuRegRhf1TUNO+11oweM1JI1I91nVX+wobnoZhYc2AdSTFsRha+jAxs5YicwEOG5DwaYUE
2R5mjvK9uzfK1j0ocVvcrePEnpYUJbe0H1BSF0rit106QumnOvkGZl271icfCA2pADBiL4VbV1Jw
z4kv2ikCmI0QzVqySQxz3b1/YAhCQHPR9lhrHG/v4iU0GxAGVAJZ1z8BbpkkEkDsHuxw6qvHfkch
lwLTMqPnORnSc13I9Z7OtxKXV/qWFv42WLCPXN6LzrSdrxzkjJIPFxtPiyXbMsL1Ml/DNG9WgOdT
o5hdpQCH+Tipf6zGoE03wPYEFaRZkp/vZdglswf246i5GKezHi4BM49QWA95Ux6Oq58B/qU450aE
aaJfH0qdj2C6xz2K+KY1Bwc+/SoXgglsHcX97hPw8jPLfswENTliymCgF42S2uid/4GjhK+wArsS
9JldjVWaX/+WYyvTH91j3yW+2D/nw+Ywf0C0kaxWfEdJx3V6HExNppOdkHUoYF4CLXPtvVtr2Ros
fORw5JzqgU0Dfqf2vABHelrUbQ988kfZSEshFpV1mU9Y8gSWjRxyoAFJrBpXbfqpBeyyXGXPdf2P
zA4vG7LXUc8b1AThHZ2WmH3K2SKvPQVfHPD3Dcj5KLcYsnpcZweHm5+Nv8SWjad63iCa0hUHBpms
Er1F5rCMK38RsP87YpZ3PEwBhCrcyuXrkfDZPcrc/xkoqREiOi9FDxkpix22lHtSnam516ZzqEKU
+PCACSkNc+QcPhprkct4Gw/8L27yZZI4Bfw7nMgJJTMHsyPq/T/Y2mX6YSbeK2MExmyOhu6LQqVm
FlK75AV58eE5To3MqyMAnJuNohzlF6Q/yPTmAt6Wn6D2RKuayYZ6g9a/g9X5A3lxDqbnCHH4Gllm
d7l9OxIytaANIRUCghdgGKHk5mp2tcoawDtZxX0UjGBMUD2ekfBHsWymNUYT0uubYoYCn2SOaYDW
ktdCJuG7zcv6z52cQC3Y34Qy9tGmE3ZTpQgJInEb6dV186Vss1Q04CcR6NK2aCRwjIRllhzRbnnL
1f+8iV1nF7CJyHwQ6A/vvW2oFrpixNR7ibjRwnZpWR0xSLy4K3uLxWTI318RWTp0EKsUFYqPJQg+
vqXrqtkYgz1UBRd0n0CPf49VGbmdIlpBf+AwPscOLMOaxABRaZwWb/WYoE7USfT4MV/OtT3HfmPD
ATwk142/oj9zb1YsltbvJu8b6jZEDgNOpvBzulwqgpyT7xS4cq2XY1TghGud+zAdRmvBwpLMRTm1
8t/cK5bXtnLUOov+RmlHP7g30eAZ1PxsU1Jtr6FzJRNbNHUwOMtDIqjAoZnLLYnR8b4XFo0eVET2
5Q+bMTI4cihDNJhc9Ek7d3iNWfgleeIokm1deuNP6TumvZeafKpvS4xHCbgFe3S4HOn/1LBPAqTe
eYKZe/9bMF59zMNfSaWtqU0EHMRBKVXJRLPwhux3BFvfIYjfk3eFW3CqDeL43+pWAzqsY66vDyuh
SkGvRq9qHbq3yoL5Cs6y/HYSxW0h5YqotEseKjrvuTu4gVWKvWjuqCnjp0NYSv/QA+oXI50GeKJd
7c9x9Wr6pQjm8AlJROagekMaOrpNInsoviPDImq0C0WRjfxf5Xe7tdcmo2+uP+BbbgLCGwm8EPLc
CIKQ6/GK0GA/BX5gxlxs9Oupw79JlHtKPNltj3h/j6y3UItOSAHkci/AGyfjK9bWrQU6pyLEeXyi
p5veUt+bcJsFOH5O03ex1oP7ln5ggagCUq2NbreshD1259FgFUKQm+gwUP9utHBstkIL4JcUp4DW
VxvtbHSFibMPAUtGf81HaAWqrNTz7HPqGwjcGDDBIWBFoX0ybQ/4W4sva+ygZnqDHtAhOgHZ6caj
NjFz6GVZVBQUfKfpbqRLNiYaVeW8nHvljc3Ahfgd3iU37EP1VpU40iI81DF4C7zZdu/LIA4oaSWV
KJiwkbH/Ggk0b4t5268UuBD7fxUJkPAGOTLRFsa0bJS9SdBDJ81i4HqYjqFj/a/TFwkZvYng4CRc
bjOtrIqBKJHhd8lEMAicMRrTEJeiLQnSmixC0FP+qapp5yoE2v+9FtHCKg1PcPWQLQRo/QzbPNvt
YWdp5qAbGBgZ88hMIVacBt+ZYd4lezI+lJ8cciZdo8adpCUXyktNJKGORvQeOg/sxemIjPbp5tx7
Xdd/3I1GwA4ZESOeLZL5Mi4j4rtoYWHU0wERITxgQ3GOfOkv0R2/uPaoZgEQaFJUrm46slnCR7no
HdaMC0ZV6Ey7sNm5X08VaiOHavdsbz9qrOHdkPBQIGFk7Fxg/m+9omx6ozeBHcV9+sgdx/uU/OPv
tNyV+/UdDjOnu+ZkNA5s5cC+aE3MRbRxrbFKrYsWDrCL5gVJiMTPh4L5kuIjPK8IIJeewFTigdwS
Ryk9M9WnZIm4FbHL0nWYGSQ3+94X6MAEZ/VkAxgVTpLURdlXg8tjIwJPPOrRn5JSIYoaT/3IQ3bf
/X7ZIUpXs7SaRv3NViywmf+XqWsHpQm2mcN0pErYEyb4yOmkkwZu2XDlBPg6MIHA8z/T6D2bSLMf
Bebt+EP3UzFA93h6xyiGm0WB8/8lz1Y9Lx6cbku5/YbBLT8DaApn28tzBl00x6JjwPru8j8zU8BU
e8XLc3DEf8tDg57lMcw+WSQxB3Owg5nuzpE39sTolmvzX2DciVGQ0NwPmIvDefZ6SfhnyarzbFca
HUUIG6WmSN1o76Wp7oObEicVye8wLSi/TtZWxPcBz7wbFuhOKarpONN9/UzMvcsyu0uTnVSiEy5R
8ZXr/IMOhrU/+6/3iQnbCAlTl9o21B5FNFiKtngl4d/UmV4Fi4tinjq9LyF0G2pgAGpjXeYlslV/
+6kcegVIBzdCjXcYULhMwjH+jtAwg4JgF/KgdHhTCMGs4PK5eg5+v6tzPOslz7kB42bSc+5BxZf3
WceKw55LkR4dV76OkPBhDF/nV8pS/q9/tpC8fI+zU4n/Y3e5WB4PF/1bnjYJc6RyKSPpF0Ml0yGb
GJQSMCmJ8eEHyTmxLtT6WTieIAJao2fhFtE5fNiEDcqxjqdFWFTLBbIfYSSls4lORPnRVk6eiL02
VpKoDNv0iLBglsN716t7NNWtQEfywxrhvKlyLJ9LYfmVcQT7vQwDFFw9OsShJ5zoTWI/urAEzQH+
pIWqa0DWrZpmXmWERpWsT4/GNb5/SWE5jE/fBhWgGAYWG1mYUjgxQPU1R1jpeBqEmAXw1v6X6UqI
JzPLamK7uw3yogBvCJbyQuVbJ/CtuN8kPNdjt+zcRlFyU64ZtgI8nsBkWYK2iYtH31kKOhJPZ7Ek
zaXdldM14J1RcI8TUlc8MyVtTrZVFIsjMvTnGeW00mfgvugTexrCkwsXPjgY50xFuIj0FndA0Wv0
jlY5dFPW79JU1yDHkvwkgWXtkjPCP87lF61VF8ysucBCnTweeOV+kHNMlG/N/9ZLU/IYsP+2az24
JYER4VCn55IvrYmnTP2V5Q1DTvHyZp4a5amCdeI59NpVwpTP6DXklujy1VIWoXacXcqMXpO/Tk7H
yMnfchSN2UU9skT4Z1TimmMdsP1O/LzclWTjPCrqkoaC5sMeJylNJVVQcga2xDr9O+nO/itrkLsD
SjckWUhf6eTTxTfeujxvVw0WnMysNwSj5pLiTIj8Q4/NDyac+XejEfCufUE9NYQQQnnzBRmUg30a
P5Bb0jd8WFgSTxADr4u9K07R3rT9OBmnGHcFyWCgSkkt+e5Qse4J4JQdNfR1u2bDIn/KMcyNBkvY
Xcu9a8lsUz62/VpGf+P5KVmKSa0fvU2zQnGnLylgVVMLYyfVO8SNqPWdKDcEnMABbdz7YXZk8309
gJ0KVB5RiPrJlD0IC6F39k37Iby3A9VwLIUAGkc2SAFbCakq3VzgLoUfpn6h33mDC5JMfXgQa5fp
f91uLIwwjXOMkdFZiAa2ZgPPCCwgEQdnQK0MvA2H4ZsHe6RUFkD6dUT87RqycSZX7ty3pQaPtvdF
jqn2XFoKxEthHTp3My/eEJJ/9RKKfD3ltdPC7lITMEoJ94dc0q8xPdYNST5zLhmFSpX24wVm9ofI
L6P1YP11EfRn7Od5I49s95NrQJ5raPRA+6AN+plsDW2vuRJMbvKkmrojGYiIdu5g4v9dHWLgsn7m
5q7+ul6M7t+149NkF77NB5ArvSsHVzj9P1UTJjOMmNLt/bGfyuWIiuvICjv29zffti5ZgH8IEjXo
H+tg3nKfC1HdOXo36mbhZpU7yNNRtxCnabwVaLkWAe0vuXWMTBDnIPKWITNdmvWohd24T1WHu5vb
U8z+KDcWvfYo7qbOSC8WqPnC97rMdrAChJ3dMOEQLvtc2uzEl3oapRNw85Dg52+8oFwT48yLNDRp
kXUCeax/RKnLSaDj05ZEixH+48yr0Lfy5NkIgWdNOrIzrMZ/2FQbyanNwDjlI0JtQlXiLumCVVj+
Fd+BCLADPKAB+SCcQK5USdajeN+TKaqGNhqFUh3BDbtKytaBAd4dMfWj3uohR77TVJG1kZxFQwcz
rAKS/1F65Uhlx43gMEwRNcVKoTXAPsdLC9OBcDbIeDgXgV7bCW3ms58qqeVQeK141gvSoVdjXXGF
D2F74dSlb1u76FWYEpvOtA5m/ba5PcB7WApxDiIWuYVB+mNqPekEyQsbO+cWqsiiPc2F6vihc4on
RJKahceSUAofIkFVz2uzW6L62MfDhDdlk5n6ZpHRFn6WlfNiOuBvhN2UhTQB0tfkG0fzzdWKzsae
jUPKWvixosDPsgDi9p16sAkpoZjypW/AaYenHHaG7eG0XNq4pLW51zOdIu9rn49tQHbpmfAA0I0P
5982kmLgTfaQWXOubCV2HY4KTtWuEDms5rtsstNf0NnlRMAAL07O9gmPmLaZGdcvt67PlZbXzVoO
f5BmctVlRSbZ+PZIMSZQttMLL8sES+Gm3oKqQle06cciFJCRraUtOENA+sUJMUD879jwyhDEnicv
rzFNVsIcAPvWqDhJASNPDvnfFuSaKMKHBjBzJmtqR1P1DFYyw40p9g6ABiZlVE9V8wg9sBDc/6u7
2w3kqoBfvg369hyPoNqsc3wpbbDbz/gXI+b21vbAdNwbj8rUh7WDOnoZbwqfz8dsehK2Q3lVBg3v
oIy6MfF+Waa8ApmxObuNxbYX3n4IuQF5QqksWuhyUR+WAY11xrqBVX1M3Z5A7P6uTzAfiGU3fR8m
5n4maf99tg2y/XX6byQvblCodxq5dahCRMzmSsxPh+z//IwiHIScrvT40CbfYzoyURydE+wzY5HE
VW5l6+BXols2kinOSSTauPZAjjeg8C63ZQEpatyOdEco+TcAM3NbNUogjOwC72hVLE0L/Yh5NRRB
mFNCM/xFUXyRJfNmXuTC98pUTWrbSqjJtaYHe0N+lQu3PItSNrFY8AHUV0zyT0TawpnRFTudQm6i
D4HpcrOltQsZowxOiy5D5MEU8BKzGbQIcdjZB2UxNZJ4XHLab1/fAdihaHMV4WroggmVLq7z7Abl
V7PBmW2TrjfemoTY3cpvT3YWfSzpjS9xcIBeg4qzqmUxR3C9Jq2f4FsgZen9VZFaO/FbKoUUewAz
aK5Q1OmdnPo35jgf28Ut0vsfPQ0o55Be6bED0qhVSgjYnWkpxuAb+QQHR4v6jq8PT9dkp86hvwsl
LHtH1j/hQhjLSN49dljsDygUwIG/DFfE8SdfL51nMYs78FgbyC9ipIbl7trFO5kH1IqyuwiMIpIi
FvYTl1wFn5p5e58BYFEjczjeyzZDByLwsZDitgR22JjCRTeiA1WHbfy5OKGsQ9H6lp+ROzhdCUVZ
l11fVIbEtiPDszju/mv7/sQvXQI/Q6IowZ3enZ8E2YzXDHK8wLY1ZtSXtA4eLb7hdzbvqBN6yBkm
Smhxt0QUV7nFobMq6Zi+u0y9jxGGZcZZGLVdzcoy+dypW8gD4EDTwJ+xo9J4b5L28wFg375IE23S
PjXNoFfXU3krcK68pvZhsoYkJ8YyIYADlfuI1dD/fRtOuRvoGkKcM59HCyk9aQRd09q5uY775gr8
RFO9tSgD7A+O3eVFxTPqOZNCZK4aW08/rXaH6SzTAtdYfyZyVyy8wluBPzgovEkH7UM779x5fRA3
1vH46U5J+0HlVf31BCAUyjDjSrHbZq5FBukCHH7clCnHpMKIpkgAZTg8FA5Ked1F10HtbVR4Ps0E
EDePaoqVCTEl8yKZlJPdybo73Y8H3NBTdOyehJmHeMDjIgb794zmq52K1umgHjjfWvCSkWvkfBfp
BqkYa5Y5OCroW/fRyP240ueLfnw/4Br8czFypDgVBdh5uwAMSUsr4qonoK7jv0Z7YRPgxFfdsjtS
hIsoWSvJZUG5eQVrDt05mubvXvUbds46yBdrATCG18BWiDchRGbScSgq3A1pg/8wsfnW3YP1nscq
s+Nb1xomINda6vzV66b0XL8utboqkjUJLk/86vC89N544G0kYH7qFTLm2EjzwoJhrD5e98gnUawe
7q+P8xvLdT8lEMFp0YkeRgUh/TTfh3lXKLODDv8+c4gYb2r5ERI44nKC7eklnqTsJ9/1XGuETX7Q
0LQ/a00pR0/GW6X9hnCgPYSORNAiGlpPWniZKbCsyPLrz86NzFUrcfI9scmbygYf6YudNo0qqlf3
qqiSmVmJNcqFXnyBV6p4pPH3BxkhIj88oAg0teIee6sWqh1HnpjOnicPTYkhrins97yjQxtRubus
jDZkEn2qC47ExLfsKtjp+POaNcyJ4bze6NpzUChloEgyLBCt8rNRWkVHtZeKVmOXUVAhTdG+XuiZ
3WwC8FKt1I+sRmdkg0VdzJk9hENbKKbu1fVjDKp5c+XK5ciIr3Qv34bSnKzFKLWMpgGODy5FcqBR
EeSAUzqfMRBvWaoxODjKWIDy8apaSyilvxGPQAUfyGs5Oic5pXK28EPtnAeHcxjxTvIVpE9MUGeN
bjGeY3e4XChY7ndvAz9ga/huOHA4u3qkfth2qSEBFjs2xdMIBWLu+BkT/p4cZsQbGTsdXZdxZt6c
wTR+QARp0DqgFP/vLnpYL0xaVxk+dsdE1XVtyK5V67QGvyRzhOUGy5MxDxU4mpz4mGvmI+tH2r22
sUpD0tywtoxb1VvAlbgDWK0xdedYDZB4pzo7Y1lN21bY1JBoOR+2Ow1pfs8VzZJ5VAwguWrkPqjC
1wn4ojhE4lmeLrMTo8hjeXm0HUzv/gtxnSMzubjFo6IorE1fK+68SEwTU4eX32qYVFERGjwkhZrZ
RJb+Y5Tw+rFo4dx0sodw2LUPbcfQ4/T0ychdwnK3Hj2mMeZYcs/iI1AyzQHbfN0Go5oyeKYyzRjS
qvdrwd24evg55saW26yRJQiR99gIJHu4FOQKVIYsl+xoEBBZhPNzXNkzY2t2AR31FC0HIIzS6TpU
AYQjBbnHjDPIQ5kEn7SjNTpbEd/+y7RyXj1Uwao2Z7fLf7SaZE2hwsOyAxcH+2CUujHFdd/V7H+8
xuDZH5WAS5d4TAnPwfSPTGza9LbEiT9sZ1rILcFSTtWyclS8xiCQya9jxelYUx7yWas5m93Tv/Yp
o3TVuCwHuKYqVg2ihXWKMH6UZBv5tIzWptIHtLJPd9qmX37kjW7XxXZ+MS318AJYEbHQ65P+N5a0
b2wTeZYxgMStOUo/nrkajgO5K7lAwTYRZR6y1QLohn2v8ih/wcQ9s4ec7D9Ev8lw6xdKUskcoHin
V9c1M+D5CeEF9ALi6JtKTJ7kzRvNv4ceTM8wrXzx7Q5I2Hdn9iQYECKZjXDofOfisIXHKobBYiS7
KCTPzLoNxUcTkUseTtjex0HmC/nsFJDsPtTeBTObcToldOLs/yb5nwfu8tzhJbfpeL1PBmpOJZPd
PlRMyNAaFLMvbI0UfKPIZnwgrABwIHw9Q5t2BmuAUAhtMHZO24e+yQ2wS57NX0CjlB4o3yJieAbb
OanyS5BQaTuwt26JZPyXACfvkpt/GIZxxcd03/fHv0HTHOaHiwQhhHvK0BhnLkGAPjL0zSQ17PJu
sRCF+4RWWY4Qp1vWKGRzOdwHP8LGNi35iV2sfpwr3b/ixBa6R9Ro1oLoNelJbWHXFX9cBZrJ7YgT
a33qrYBHPVFYjXI55HSoXXIWwJYLZILY4Qh622BRs/Zh29d+ljRzMg4Z69OMaOzTAPmS7nSJZhVg
oykO9ObTEO2rDe2fHMsRfwwSLiO/pAXRl8m7gwhUmJZGFlM7/l7r7E9MVdGZXoEz56iT2N3bewys
8IOVidBa8cKXHxeReLb2DIlh0PgAjcwk9TWGs/EnIBf/Sqm5MvqC9+3ZvThyOLAzioVf2fVhb9iu
C4c6SNcWm28phMXWN/V/FNKYXOCj9QxCz8VcBsdtWq27WfRe9TS80aGauU2+ZdmBd+1G/2k0fqyG
rAbqXu1QICsnAfOkPl6VPB5cBtUFIJBVn7j7t3ZAcywmXaUxB9WhdzeJDfbpRQOLCJqBOpgh27bn
K9gUe8rdaQ1KVCQhGIXlky6f0EyvaKREIaTwKVkRGDIwDiL10aHTTnQsW/Qa7NdZA2S0ruFSr4Bs
Ca/iLFPk/vYb39XJ++LS6S74t98FznUghaqjN1Oi9OqZcAZM0byGxW6QSYX1q/epiDsHsablrFMn
ssDmuR1y/ODc0caZ08y/4gvYiidh2jYaf/BinRZnJ2uYGabojIEi5WxSN4pcuDfKPLSAs4ueQx1r
n6hS2NyePA7ER/eg/qHajBtRG3pPZIrNpdGSTxZm41rUtiZamI7aGQyAFA+sk4mvPftdxBUBk+GU
GOOHsHwQNEMPiM578LXqx5kQngercBYS6dS06eUWI4pyVzAYsXMKcmmQBgWRPuborzHPq5vBSIhY
rUp446QCEqwV89/erCFlpPS2ecTR1CRQf1x0JPbClf5vjDGyVfAh+WSaJCQqB6mwkNrXVSiHkvdH
jxMUsLbuFMZm5j8jmNDAlE2BJmNau4cZt+K/U1oimhdIT70+TWrUqs1hyMYytVExSz8gAHBGpN8i
vA9uFsp/4zEDhx58/M4xcImUSHdJgu2NfoP+38ji9coFzMIZIkWAz6mm5bQPTbM9vJUOFmTFYGoY
mV0R22K3XmsnV6YL5nl++As9cejjDzyJn2tYub86AUw71kwjfAa8Q88x666e0sdVdSPzCuYDW3fp
u5q2uMOHY3X/FqwcXa10oyVu+eofy5NPLtoOiyJcQGLqzfd9I5bE9bgQelX6LWMLn2lGZ5x7KS9q
56LvdIYfQEGoI90MnR9L4L/+EErKttfTTO9vFVvol+k38eijFmuOg4K7R9Ci46KcvpEHxy6pKBBd
HMzSoLip4Udf3tLUD3WiwuUtTSOccH5gD/pxMNjKTAo5xLF9j1EwQqtRg427Ga88mWKIjUV9vDij
vUfoMg29ESQa4G7R26WHOofrsmywzduaKA/vAYGvAhWkHU3vqBCBGgdcrjAv9XEX2uGa7tLiUbsU
dJP3MJrjzq5O6yaNOtt4O4XEgO5Xd/1DiXnhuKdFET8pbSA6LCJ8cIz5x2ZLFWAbJ55Zw0zy4Cso
0J900rD5IG3zA5g3avw2QIf8fljgwkt+yWeufU09t9E7UEHXrsZWrUzYkhhLfYfl3U5Zx7JxDJBU
j/HLPpX+CsnTZwVKrJTCxif/n2Bgops83xNLFRAL8LsKO14IenUb7/WyGxo8hu3JPTy9YubcygUY
7wi5Xsf8h6bgLks8QUSnf9q8M7u4I9jCV9r6ivNFy8u8icI/7c/nUg5s/VN709iVk0g7Oo/SaobZ
ds7HnUSphwo4h9pDQgHzxxaiD5WN+r6pyOMec+uJNrc688X0t9EJt4M6M1P7LerYhKYHSZhX/FfQ
13vTxgaMMNWGDLL3QsQmNTJqW5kCmnvo13zWgL42L2Ju+VA2OQ4QrQHbGgN1v3a4NmWNNBdHu1m+
cVBVUoOefWRwjzy5JodncXWmBPVMI6gIvGbXkE4qUZ+i+SaCt9Z2wcwFX6GovB8zSn5aCpc2KQEm
kAfh2TEkOb7oyTI1HJySGKPN/OVGoR+9FJZSyfnwpmTd3NMpwNbou900olk/UCXQdlG/K5vRnsOR
2e1FYBvPHdrVi1QL0nyr472/D+4APafCj0ap9vW5fAwNdGdhmBeJVmJj9nUeHsE57Ye8juANbN3L
UY+PzS2Ty4GDvKjAMw0Lr25Zt76pOeOeACvwrssXw797VwdN81QHxVwFIC83Xt0L3YUuaAg02r5l
EXJduWT7+g5lGuIWqhyyCUsCoP2sDOGYdl/IzdbnxEbcC0H44e2Aw5bNDYLOl6jCKP0+44sJhnLr
zr3Jh43b71qqRjGx4b6apZrtaPuM8MoLgaF206vw1oP8iF5ZmP1K7rvUiX4VRGaTWPe916lvHjf/
vsUo7ZUjyZizyQIYeNL502tx3j2XFPCzZQKYIJoMIz02EVDqI6+WWRMxzFnkvdwWZwqR3uKPNgP1
UDX3y5OqR9KK0Kp1YEEbv6sD/ZSq/RBwvNkMjmRBCPh6peTQprLkSRehxUdiMYJBcs7q+EOsbT2C
4VWF4/Zx9aRKCBn1IcYkNbVgONGq2tYIJr4sG4GQ0YWPBtMQRniPAqN6umhP7VZIAxwgbHwn7a/e
QacRWoeReUcr7baLqcft7RjyISkNisNuBSlpy4eN4vwMpOdc+yj9/5rMl6iDLV4KXhyJdBtQKDDG
PznNErOpGXQ7OvOZgwKRMNCHx7uEP2lagOBtaci9Fq6n+zP8OgvNaphTgfMwbl597iQ8mUQry3Pv
Zmklu5QSEVCjrd7xpazXwWSkqJ/s62+Hj2MkPRdXVvdHXprJPsGae4TRwdwuYovvPk41XXYOWCvj
fU1D13jjnpEUQ/MRmBvjsOCc6GX8voahdFGQUMoIFoGT5OPn1RD9O0SlQ8wf6kaH4qMJWkA3/8B5
+5zH+zJeEUMgQM3EYwKhxmWyHbnXGHzJZjgxElUg73p4gkDF9FJYDf2QS9o1No0wL3eFB6vm3swX
Sdi91aR1J/gsUiifo+DJ+Mi8aJnKpC05crYgaflBgg4hWw/eiLpFm+sJrStY2xzyitG5aL0XGh2D
wqKQfenwSXrtOSGdeRTKduZ+2n840a++bgQie3r5uvVfVroltNrJGO69HQco5yI0zrn1VmRz+jAz
xrxGvs3ExtGER52vqu0ToSsVeArdBChIlDCx5hycm8+yGYkfBSA+JSH9lZO/PHM2SkSCLuxC+c1b
Whd4gJITyE7FqVu6zw6Aix0UopjqFlvEf1yRS+UeMxbbQ/iSM5AhOnIoitbM1Yb/dW/xn3NGlW7Q
eQ33VPSbHduirfUQuoekg6UPKfDMYvo3jFOP9IsdUZ8yzTojCCMDHUYHEcKgYxgVtwPxIum2LHB5
erxisAHFumFJBa0XHJL4TV4LcTzeN/ZtPhNc0VTqn29Pbzd2OQhX3EDD2BrXLWLHQ2KKN3vRvFWW
VOV3nK32W06d1MVzcSmvsLSZErSj17BIA0Fi280maOyW7N6MkI1W40VnWLH6qy914IPS+lX1MWaD
p93aeN7yJv6s8/ms+N6K85cRIueCN2JzT8XNQUhwjUK/61FdH4SjoQEYj/DQXKHCRH4mh1XfEUKT
Vhxx56G+ktGPa9YiNUFgDdrJQgWISfguBE4rI8+/s2Zr/8pp6yIai4Fqf25nDHGeaz11MG2vFKoC
U39JV351Z5To8Aap4Ed8I3Qq2AeUgpZmfNId+A3MUzXuEOCB0KJL1CwfDXWnCMtf+znNBlO+19O3
LhOC64Y47Q0bcM57SOj12xxdB7IFLy5HiC3t8WkQX/W6zYW6pZ1OsQApJKSLhzC08I2aaqOZRffQ
MjBb+IW8hgkPoLdp6zuh9hypqxfSFUabQxs5BcQwp9rQzRBkSNjpae/N1yv3BgeB/f8T5/Sos2pM
smRQ2WnqjpMw4dEYaKfaAPv0HFWatVl1eK6KdeaBrT3EA35E7nVIQj/4n+hvNIfLxjhFTPBHgiSW
t0PPf2f9B5X46CrZyyJNSxb0HIIEM9j8tGh8SakD7yKvnfymIHsLrXrkXxtumaXL+4PNFl5J3FTh
/Ppd2iXSyDcq3f5JiYcXvyOqhc40JJ+o6fEk4TsUxF7HNV9ruNBciFgAnQnfVCfCoYBWKWjrk+Vc
TgHHphPWd8ZKHyLGPDfMubFuJgiljYgXl9cleKyZWL00XwgJGxo/c+1XD5db+qKza4EBJBgDSzNE
z5TWWsI/bI6hFI8fqbedRAk+ywN7OklD1DtUjkuF4mbBZMK3p0zLupyrnYw4V5gNk1jbqebMUIst
hNJXDwljB/Ym+yc6D+/t8lsuYn9hr97JTIf4iqlUBjJlP9l4KtVHCljofHXhtvY4jL6xx1aAKcZ+
Cd0Drjf3Kq40Akzru5GOZEG5qS3Aomt2OY2Qg2g62aV+guSHJ1rS2Y8X0UWQ7KCpYUUxZ9Aihg6B
k0Ot0zTBgkrD1d4JyIc6AosQY7GK50ez7pnGFArULZuON/yX7sACagljacQP8eyyZDqmYWqn7THf
nlI+oIUz5pylw17lbj4xBZy35oB4uXRV6fScjatYhah5yd62aakp0cW0XMGhgS7aVkV67zrYzL2W
Ae/JZbIeUmZOTsrvOvd3NMz5MrKMQJDMpvcC8/LsWw269fywkfhkVyGNCqjRYfT6vcJrDQt59sQ0
O/vGlJJK+Q7ullXOm8u4WJ4sglKEJB6Lw1tGTdSTVSxuDfIQkxYvtjXXoebilSRHq7BdQZKFi36J
Dz5VoEkzVHWZXEQzlnH1FZTm60+YRHMrkridA+HlT+ikQa4buNY3eKvUmiJxDvkbL0fubfzf24Tu
WHlj0T2Z7YfHcKtPVcuQOp/KZpYsweMIBoCFhkZogcJ2u1v7m6kihr/sd8vNj5+91SpPWwHlLN1s
r44KP2+qwBjMo4NhZctmNw1vKAPhS6agYngk4AZhqIdSwtB1gfX5M8Y9B0123PQmYGvZUQxvoDTU
h55s9IrYhXg5axL8LreEbAf+h1WhN+16z53VTcIXkfex/9P5Dw/CFR8Vm5/jaXhH+RntzXfUtkKJ
WitaFC9jCtk5v9eGYTGkhmWDIL/EkE4Cscgn+dFafTXcvDdIijhAkaP0GliuWpsO7HVJg958gSMW
39zSgRdm8n3tTwOycm2v/MVR+AKS/3C/kKIXFwkpsKVoZJcI/oa1MhiEbsr8JyMmIDCYndbxmyX/
OA23bkuE9OgIsO98fHhGtlF13xvW8f1M5PYoCGUQsiIXUF2NHW1uDV6IoarpCz5/1Q8Ku3EakSsx
hp+udn/eNs0gQN29tVJ5Fla0EfddvpeeLtHB5O7NWI41DzggD9454ckgaTnl7A3cuaX/ItBsb/6w
KeTsRbftg8zY859BlA8NFLrNfv+Os3CSPpkmyvk8rZtAdK1qGaDrv5AGCNY5rmTlBHhbqfXOAwRa
3pT0/RY7gvgQ0JJp4AK/m7YEX/uBQDUsgflnsB3PQSpfH9WjSiZZQv9GM0peBrn8fhlkdUW582Fk
MappdqxpikfKFnOd0euJlLlAlghZeNTqBAHLHoVlZvJ76x5IGYFceYLUrafaFV9ON1H7HCZAts20
Zj1TuGY1TxTiU5grr12zkz2Ql7mGRtWBru2geKr+B/Qg8hwT9NO2+kwIVydbcWxrnMOJK3opDaKl
hYtivIFi82NDEqdHxn1/mBbdy3HTEuT7i9nVmBRFhgqXEhF+MZLw7gw/xkxWsSEwP1DrxN6iPCKg
fB5MJ3NjGvideQZwnhfCcKaQT8vsnbEvKcgna15k9EXrkuKJfUG4XvnlSw0VW1MTXFUO64eL28qV
pF5X7o6WNAjFdz3aBfO/4baeWh1141+JC50qzM+hQ3wU6f28qYMTm41dRsmjR4y0z/1oS+v8ChlQ
JDvZcSy/tJzTjkw91y89dNA5rIf2ZeIbA3s3FT9AJcs0E78vM+NMKVueCSGNPiyHPJKdAP1t/lRI
/21mfoH7m7aXAfjMmtjw59hmDSE+Dg5OeUfa1hC91NltN68ENvwde2xnVoqEUhpi5VqjG7QjCPfC
6xZHFOwYI/oFGQiH0Ql/ErasGw29pM+SdQ/hUnLSZZIAocaj7ZwNEuLxRcHY5SAunmrkSkTv6eb+
LBvNSu5QBIUmmwgg9xNXIIdVm1YIpkQ6YEAxudi4tYPiMD5DM/12n2sctdiH/1JCgV7g3dQ/TgXM
WMuHlt1PYPKL4COF/F7/5QcAHlNU8RpvhOS4rutO/PaG/NCVvGt93mjlut3Spe/0Pf8do6WZ3aWB
w1HpUrqG0V99uGhGS6QAFDhvVcajPKmy9mvfc68U3WxkgIpZPL2W63Go3Px7qaiG8XNCXRMCMi9x
nor6953+ZgLG/hRwrKWRJ7WhLrJzceuRNRWQdI4ri0yvN1bJoutrSOSeDSM95Ftla+4gnbQ4AUQW
m4gn3qrdswfFsvw486/s7mQqzjrj6PgwYNzjK7IG8uJGr/O6HkzjC/JINObJgEYFBrFbOK94TwV9
ipjk/kBNRNhjmYUZODxmfn2WcoNrInAEnXkYRo8urTa6rygHOmcNojFDR7ftSJlTh7TWzYosKSHb
9GIGnBoiys735Lgt0hircqcrB8fDLe9L1SZsGSMELN82FOSKbp2stxXnOhnjKUwbkLruyrt5jSB0
fnGRAnnuq/7h/yzlng797/1OTaqUrK2mrRfa74PsUq6hSM/Qri9ZejLe3xd3e7sbMkzy+f0dQf/k
PfFxkG44PhU0WkmA/Kf7kpXYad/d8oNBCF9ylC9pkS0BcEG397HuhAiqlTQjo8NRhC0IYaZPMhjN
XqMly4+g6BPdOqIJv8psJaA3y/IqTiMIvNILrjsMO2KHdDuwVvyyxhjYNLUPfxWBwlD82vi3erUG
cY3wRXVZReFD9E14U31Kq2gt7IfzHR2jw9c7i9oeZv5w41KZ31nBsuNqJbAC7H/zAPtXgXdBOnca
nf7emPe+vsW6fbiyZqgdD58/guQ6x0nzAFoU5/I4vMY44qDiy44/+ggQEoFGgV0g3BhWIStYGieY
3euqv+LnnlKtzPS1G8DihtGOD7GU4xRuvOBRN3JXfWABleSdckkyyN7PuCVHwFxMZAqWd1+koI1Q
GB/DPjwc4l5EURkv1+2+826fY+71tvtIqYktUxtntAj+Md8dMjiChkTsTuucgfgy60N82SoKeFLF
tDoZytTdW1mHBae0/SaX+IjMGwrHMCjyS1xkZ71FnaAT52pqIeKZn6q/Rog0hyMp0U5k25KJ51ir
bTjaUB3SrFjNvgPeFSdy67WfLYDhMYPuSyv5Y4/GlT+a0hRPEGAV7Tln6NrcBH8ijfYgYnuI+eBV
Ahy4+D3vF9OnhnVhxXc555EexW8RWq8QqwJWIbQmRgtxoCCNY+FrZQzbwp1pkh7PqBPjZiYHqIaR
g0RXM3zi40mgqakQ9tvBC3xA75uR9TZDFDgZ5/RAndpLDJ9UPvl8cJPVdu27wvPqht5rIQKKP/9A
AknjDZjGj+NgYjLjSJ6q8CFWJFKunjOZ8/ELBSDjU9Sx15tGtBXlC5hUuTDFNCKMyRUF2ZyNHUqD
KA4xENE+iFne3mm158/XCbiIl859Qge4n7nUO770YJSEqTM8iDUUZXPgiDuLxeCluAm0k+pjEhZC
53Pu5ib2qZJaX0PHCzMtXInoT8zWHx/h4hrQXbjFuRIwHBXdVMN+SN7G1LKw9lxUovZIrt1W3kr+
c5N6hf95VsKs0U0x/oH/zbnPbIYDXwLzSS5zaPi02QvF3V57d7NISevvHUDO3gSoUj82IzQ/2kuk
DcQIBvtfLWQrLS3r8TbxbU8vTvuDamgTZSATDsY9Q3/cjui2qSeYj+kPtWvy9c4ESShiiI8OBQvM
yHtKMK+rZRTYdmbNpH/5QpGZK7bM5Eewm0RVvG+SzFysoCQ6kwyrxnB6pW0JF0SLKKRWFnpuas75
hLZBsO3XTy8xKCNYwuM2l2XaNVKGdYkQxsbSVhFAOSl8hAe2pMPRBzQIvWFy0NW5SGTJozEhe9w7
2dzatcXjyOoS+fveIPFOxoz9mh0tgf+a5YFUr6NaIotCKhQOae4uNGQR83EAfF+aW5bn6k1rkUng
+1FCLZ1MTRorNAO5S3XFCxtv+hpnayUZHdnnkUztqJbNPybkjuwKOGlTIAJA2B8BTHASdQF1++RH
DnzeuTzOqfFT81nTKll9TjxQbSy9lhyHya2WX+bO2p7ze36XszfuON7RUfuHsz9tN4GhPpc1PWkD
DCAjzrkEZTyQorBiGu6506Y4hgdeHfgLBzu/tu+AgGXFZpg1O4LerIYah9EMFqsNYlmvma9aKC5f
MfaYiqeN9TvarDzMzP3AwDVTaatQFQ7kGXGV98lwimDH0ekn1Yy2cSo+abSfsBVwu0mBC9yU6Jbv
y31lrRQjbR88U1mG1mMg6xiPtiGpce+rIwONYo6V2h4dP8KXlvxDDBjZIy62s37FKum6V1vU25ow
n9b+ng9zZdLP1JUiY1bxiWMURUv6slA+Fqnh9qSuv5JFC5dRhdH2e6U24q0DDsgzeOwdks1hPz0w
S5/LHWd7JCng8xPWg8TbBofYX+G5MSdLmnQJFatTBF6sPcIszyjivC05Bl78nuYJMXgnKvMmK3WZ
ZIPe77VgYG5LrYPPj11qsH5+ZGzML3nT+WtZM14twzPa7OhLMx/4hxV7djbebWooQ1ZTI8/r4VHE
Cv4u7wI+96nm1iMbkXoe/dZUej1XaEsrPA/AvOmxmFyVdJ6jmtDp3WUZ/6HWrfbKRSX/JSby/t7Q
p0ZxmKZVPQ2Y/faaLvqS1E1ovywzN4T1ujtbIw1+6OOJKkm+gH+ivyb7zxvuDynZgf+FP/9o9QOp
0nbtRcwDni6yg844AvdXydNFiYbfXPGZ2skG8lJ+/NENqoLSmfSi0Ml5AL1vVS893ikZwh1cGAxl
5BxOwZvNVsG4wc46XOUnhqcxp0IbY0qTdeej80wlpbAraLpYOF23LpgPhR/tonyjhHoFv9bPMBLU
cWJOTDOvOc7+QWJZpPgG7l11cvjF4t/mWxc213FFsN6+Z0MIsmnEpkXuEH2bSq452OPc00wfZtqH
CMOAOGtLByzta2huCxBSLDez3DG2ypfpigqNNbaX6LPDifN/u0t1zi8q8Csb5DGAAzVLkUdhEvhr
E/otzdpPd1perEwd+Z0eHAwjPpA/VEkcvRTJLcv4UUXXOpmkFbZpO7ki3AP8ECowqn7cjBuB8Dm3
IM1Lv4D2ltAR85DLB4rJI53FsAckP1SCA4nGpWTnJl2VfRAqpRsgoMPRuQJUuqbiz43axsSvE1KL
BJ2163rZqbuB5L5HHdBn/XH1zOT9PI7h29pJ+7oCdbZ6Fp+pHt69ppfNtifChFXQK1syeas6j7d1
9dkElP4nXyopH3rS8eJJ4rqYGr/X5cCcY3D5QgT8d2S1lUJzyVsKR7dKRsiAP5FgN0KwfOPzKKuy
2mht2d8jscATinEzjjnl1T9QFEhUzOpEdKCNbuVtmd3d/erBy53a/rLTtUWjcg+7D6hzPLTLZRac
VtKcKErxqcuT88yyxJOdWlb3UVDQ8bhd33lM5q6fEZjj7cwdTCXIleRHEE1HPa3z37GnIHQ6KwXA
bDKXSZZOq1NhFoUfC4TzIg5XYuT23IQxvEanTxhons1/tN7bhIKeINyJ++PznDKl9POiai8qCTYA
lZF6xr+eASPEGdxoggXyCV2DsEUcJ4KIHi/qjajBaFKd5LKZ3PAhTou4FZD7g+pOfgJ/omCppf6k
7yNBp5tVZfKI30grVO1PTzL2BEvSM6NQ2LOsk9FHc/TOW/RM+u+gxAlw0GvBJD/Ppz/z9n/fJYk9
v+l2x9QMAgEbi3BP9um4UaSVXwUvEdkN1x5Aqvg7102Cpee6PmEDOXXMsUge6mHgccj3zWxhew8C
pW0zLM9EPXksd4g2oAFwKNb4+PiQY+sLt8hylvzYsvikeEh8d4iJMJWuJUBN/mxf27fPfC1PcrdR
BXbHXUr/CRrz9nyPBRtV0AwKuC/hp0LPt/oHSsFqG1ZKOX4AdgilfHa/5ngXXyUk2dQTdiczkiXK
nfXt6E8LXdEafXQTIubjClcjulSNHtT0vG1X9etpW/jzaFULGYPqqo8sCdD2Nf/p4kkZIBsvLaWK
Edfil2NYKhwpbD7OTtrVL365+Yf3nLKW0ldZRxRl9x36OkIt7pudZGUkLDNEQUVywDAfaTB3FAIe
OGHMvVasAIONIOCyaiZm+bwqv7znYcmCHNFKuRlmN2a20HYJBojG+3N0/kI1i/v5mrQEP04JiCaa
lAjBFeq9zWqtnC0LVYS4GzZB5hqsTS2mYeHAjTPgt1E9C0KwnluJtNMLVOyEnK7ASPzU+8w1OKR9
An6uwK+7U4uyW3BXEGt8Ugaw8eln/tVqLcz0W8aX0RgJPMdW2WJp8HfRs7rEvAa922kpzkYM7f30
2gHyaWyBEfkxlyeaQGQeIphUx2MDQEW990sX/OZeTnktutI1MrUH/BlsuSn9Hv6b+ABy5qCqloyS
a6m0UoCMWTCJmic1QqufA7Hdociw9C4cT88poC+LA//nTVF2YlRfDWN3t15BEd/pk1fZKEyC1ort
HyU9J/7oxo8GTT7dHzvluHjD6JAnSACPiC8BW9/11YL43kZ++obO8B4nXBW1YChiiibnXES5h6P9
5x6xOwx9hUpPW7YTfJhEQ4NPHBItbzmd05eMlfeFrJ4pIk0iX2xinI4I9aT62RFZi3Vdy8sCjpzC
iFXjMOXuHCfZvl7pfkhn5vDJSndPNrSikIqQY4NNXnVy2aJ1i4DKVEcpGw7lommD4Tvlr84+v1BI
4uxQ4gM1NObi2nUXkIkgeFG45Sb/8UTVAu8yL+y4rEIQDOYUvgEREXQshFCmxKklFjbSF2AM9wis
m/2crvX40fuLtn0W5llw5H4X44G+PfgEydqUfshwQAv1k3vsv4EXr+jlgpAO5BWM1atu+qjkWaCF
S/TSn/juN/2y9BGZka4Rfh/abkfqnO24vtlVQd60BprkFU2zay3kvAJ4ohw4LNtlor6xiEtZkgas
041ITBifMtqVNclOkZCJpTUfCFwy5wgOa+1f8/Fhm6ymVKB/YWbZUUlfLs++VBVxaE4mUKSoJpZI
tyiXrTH3mbbQ3Az5LEu/C0PJ9VDgIkWWEN/MsUHflfC+vL6Qll8TpG4d13d58WZxLBVfk7uI7scL
4dt7T2OQD+nxpKDfvMOXDdEFRAHosaZX2/bXlPniCNcVu1RPHgSnqXzJV8KH8LrVnidxXCml49eG
jPqEWEWQS/pXktQlgPU3QxO5xRx5eRemT425qLlssIbkN3B+rb8GeToX6fF+yo4PY6/ctndLIFwi
ICDGHhPCCmkFTqeeXKozV0pIKgoB7nzQlolTIpFWAsBcA9278dFfU9P6DlrV7QnQC8+XwiqLmDPm
nYm4sQF+bM3judyaQkP/oIbqlV4Ne8OOBVYH37LQTrfrwX3HwpwK4EvxpfsbEqNwguhhWMh2FW0f
Ni4SQ4bd0gAoFr7A39TebxrK9vG8fsQBdp/9+R1BoEEXiYusQJA/In8ENKVRMgafgBcV5hwHK7tT
Vv08an6mtPshyJXzGjnYfQ3lhuyZXoyrMKc6loC6dZulBNs9pgW4FUBnaB8cj0vSwE3AiVaUbioc
5agzIIAlMy28bXVBYcJ4DGJZfKXvhZHXTTpC35RCc93aC1E+qcMyKlJQSzu+zohLlUxa9eNx98Tq
xr6olX+v61HhK1d1O+yluKZSbmtW2ajx/xoQYpXldXXPTpdWrVxoP3+0CgU6pxW4zWGV5VP+Ns9Z
ozXUnDuaPzYyo6oFpKTQNSS1jUrI7VXexGYIjCTG5wjjc89D5WrGZcdMeFnhXKgMlIukXSGRo5h4
GkYKrdlaqpFXVMA7UjdFOFmyqOgx5lijh09PZN9WKXkgWsfiv8YJEeFSeS9pikE6yl91me6xgsH8
+DwPE1TgBxeX/LWfCcroidoUC9XlmD8fqAnx1xu1MLxAUzodaqiXQdlnAYS7XwiT/YfCM95ncC+s
EtVBdm64+qo3h7MXtcdaZ0xvTxaR6n5GLAFjSZ6AqR0LyVym0AXOiRV1AfeR+s7sPs5lT/o3Zt3E
NZBvwPwo4DKwNHoc5yS9oFY2287a64oPMFFnkv/YUKAQ1B+fVLy9Q9qNAQr266My+OI7t23T29DI
zibDm/KSoKfgbxskqkRcPCQQRh6mbAKdWa89eJQOxJMuRPh40Ldb9JtBXSxPToT2twPjQpoSIrkz
0v9UIhCk7U61ohNLIsP+m6Li33GkC4dr6Y+vhCfYyIue/kpHbcMQ5rqmyDfWb6FVhPg+E34fpuAf
SKkV1A4JJR6SNJXUtFKDGyyP2rBRlkyYGpH7Q95KDItWz25kPEU9szGhwHWLXXbnFdizK0TCPHQe
a9RhvINBaPadqre976BuPqhADw6iFVaeF82k5DZP4603DgEQM5UFEBpw/7fMERmx72TqIXXlauQb
fRR+kJlVP1AWqUBJncS/MkDI5ukPTwMpsM8TXJIfeg5OoOXBE0b09hIwek3weestMwt/T0sA59aP
fUEmTgpvo9WYl89r+RhTHuBKeWhVdMsxIlyUWUMxOjyYSNg7o+89mEbuoJ2sXwomfDFvz93KUqOl
M30bIrNkefYhW/72tOZR2TJvFgp565P8leffdFTYcSa2au0rxLr7r/Kg7HWrzUooWO6zVe59Jtfw
eOmKVIfFA1QTrLiz53+TNAGr7n8TxUpylFOeGgsCtY0XnsDYJQGzdb1+UgoDOzj68ZV1RQ8T17SK
UkNZuoNpfmi27miUt72Y2Xeqgx2NL8wlgUxmYG4trOsSeYWIeRLNQXpqNLvG5HhUUGTQ4r6QfQe4
OoOKrY7TV7OMzBO2HUiuDpkPrPUToe7kOyNpvKNZoxMaos6PGAu/FiCg7k4swfpr4ehnAQIxFa5o
4fHiZ8kNWyoHrCqOfpSfyJ71Tvb7llk3NLMGVRqQ8evdbE3iFlByGkqqGEGQQlL5866UMRno/iIW
CCD3s/i/KK8ngFVB3j/eWb7bYBUbRWKFoFARVujrDzJJ1XBfurjBrw9S5ceCu2hilLw2OQx/gp+X
y40VtN4zK5bE9v0tbhPZuZYftAzTGDNP/nbuD95C24x3s6lT4L165QszAXCifpb5osfwm8CSxnLs
uQlB1r27X160MQdLmhrT+NsYYmMfzKkjQLhyb7NIDYoYYMGcvoFCY/4eFGf7H+/gyYV+zerBKLGg
6Rd+/YKNZRjz/IUv2ITsZ9s6ZmONvoViAGHBNYkb4OzSIXRUTHYDHo60Rs3H/VMYZsQ5lc3ZvJbl
sc2Cw6PNpRGAcaCN90uvsZfOx/igtktpum72woc07q5f63/7bwjj3Kqr1rQ4VkDFBFnJFHbCBn/u
6NNx3jQhujis2F/C/6Z2dZY8AeYslirYLKHO8JJTcPpcVXZ6XT+2ZIdJFJs3nsgFmvNIPyr0Qg09
rXpkn318AlgTiUmFBJm3obRaPsN4jL23USzgrcTEht5NW3XmYQNttPl4pqQZ6KeJRP3LcxgXlkNn
0BUhECSeMHV9ieqdgddp3PvEj3ZW0l1YWkGoun7U9/A44O1ZIse9sAY2h6c4xKRFb5B7BJV5B7BT
8PrxbiQ4eXzH6TZ/FUtZ8zSggFEtXyAjRbfuBidj5yrnIpdBQvMwkiTZbmsHtZiHOa8SDu1TFeOm
U6Jdc05clxs7u07jusc4lQnL28eEnNSmGd8AFtWQxQtcEYamJbl40OqLPd61jpuxdoMAnX3bY6os
x9AgHamvOwwXkjmdIETHDnHREAdOhX8cVyZx9gwN0nj0FIiNVsXF5ioY84TO0pk9ZbJtMY33gm9o
1SP3ZvWGxM96GLlcVmHdW9hjiAK9QFjyFm0OPnDPmf7M5KgBIx+PlEq3UyN4UvhCRmsCFb5PP24M
gD7a+0pw1S/9V62RVeMwko/X2BmeGyPO//iTVaCv5bH9KdD0QqFXDLMv0YuqCKW+vd6irBMFpoMa
TXm1p9pomvOPoFb2Ih4s5uFMj3UTwFLFMQqzi0XeXLVp5xHSE48Ek88H/U8kInltnqKBdQOEaUMZ
0yhP2AS7fmhLk/5q2u/f2+sQPXMPvV7MmU4YlCzD5aFIbe50RZ6Dnry0KBbe+gA4VVI4meDf5Iv3
aoYgmmB5FWAgGLoQFvnlY6YRRJQCZ/CPDk27oQu4Ab4tcIp6U2jPEzyEu9AlW+Syv17uyBbLRcMl
F19NxreHmL5aoKUg4DFbNKuBQZBK0RNspJcf3edydeNaL+PN0ODfaHNeOgeqYb8AJrw5Tx0I5xg1
KMAwo4Eh7M33PJjJ2wnoo5gJN1LBuT8jrpejj6aDnG5dPUzh/5eV8s2gv06MoAhMyCuqi1G0lhVi
On16RLgJI4SoSepDMYtu6+z6T89k0WaDfDXs3DZgEeEHHMWAFv9hD+Fx2sj5sIcWfrcV54p+PXlY
65huXOqwzQaF7pggIuNRcCg/kI/lu9V/hBK3GWU2g0gmoDxf8CZ7HiMQeiLtURH67aH9HfbpuSG5
0t0L42j6w1MDMPhrEI1B2J8fkgfd88O5XAevf8tbIITGtIHFXvY2bMUXI7IfOBj4m/ClTWoiVVXg
Mj8VLvP/FN4A9sjY9IDxirR5gZkVhNaEAo4J0PBAyOr1A2lousLANWzxFx3c/WaHPCUySdw10CVL
7p38biHvDrEsOCQpzgVFlkcmFcdNIa0fkzPAAqcUbOvsikROJEZMum+WN+BSxNtyNyfHJ0Q3hwIs
HGgA3j5MqXD3IM3GAx+9izb1x/9ngmEFiurImgYbzUNo+d+5NyNVWg3FH1iEze00UBWgXc2uD/Ae
mOLjimi95XOcQ/NuX7i71yvSU0Wf4pP/qQ/n2Lu4FFTmVbJki/yr/CE7pI4Nevum1GQyEB2pDiN0
kBkQw5jP0rf7VUUJcRtcobu/EUqox0BqOYHly/Rwh++HiUcJJUdm7ECMjGgeIdgLbmUHxmhpQybL
yZqYp58VOb40ei1B0noHdjdGO9RmsWJXjmZFWXTxuMUJcm/SVctSunIXj42KguPUK00oOw8Iebli
yOLdWFXnk0Jpw709GKB4VdkTTwxGQs+Wey8tC1lA4z7jDKISuGNEcHVSZ5T91g3MixG34Ox1BGg/
GOvMqGomdDBQ576RTcWSHri2Ylpsp6GpjXtcv20SLzpomTGyuwFd7xhW4V37R8qj4Q0HPIuLz0nE
bTniSVvGpuMPNPgIkBdXSKPiFSypbYq8ViyyypAs3Ak3Y+6E1cTxIoPeLYahFn7PjKTBMrbP/Z0B
BL0G1uL4QBHWL7Nil0rrR2LChp6et00bb72YbQ5b88Y0FB4XwgHO3Euh241sojYa0atcYb35r/3y
sb2AB7NhqKOGX+BSoLru8uXxX2olKLTI+Qm89AHMFcah7JIFuwqvPxVdr4CMzRWlnhbs1EyyXWYm
83jG2Tqq+ilMHWra/KeQwm9CbRY/s3GmQ97nXso5gRkuhpCR/jTe/S9Y2bKmbeDQqwkQwT8isa0n
1ysXeO/3v1V+BVvIsOQ+viWf8IHDMUifqqrKizsCOK0XtKb26YQ0mXEvzdaAxMpMGamQC4h5N3q0
bvr6EYaIHawBxisVT3Ev388vqSels6JS2G74mZLCbOX5xIKdJgdf2uU7cP3Sh9TPZnN4BaqABMWR
MdLJ9zLGG+xzZcpT70tH5vHjC+voAxNYAzXMk/239E4r8b/ZyMHvSGQFiGu9lgeR0IZEdqDUMazW
Fh0s1AQuJoL87+aedFLe2f24HbS5rDSkP/8BMd1lnDKEzeMmzW8YWemwoSB+XVgwZKXfye0w3Yom
AbMcoqj9TpFeuTy1SSkC5lVYrPPcsbZI3NKKsJgIItzv8TjaHeBhm280UhmPxEihtXGNnyp3pFq9
5BsYepHwmxyO/AOmVMYxEnOgvFy00TB5Yz1SFPHwbXn/NPOvBzxg0379KDPA+yoTRzT4dBUzildI
zzrX6/YZtHO1dmBfKbivnQnQ7zOGNP2K1c5VR9UATpPYy+fdZ+9dB+NELJsAszCHx2mE9x+q6IYX
oh8cOnYWNe68rNIx6urx3bJMWPGGPMQqHqwsQ3atzbhh1NVgvTggqC9G3xSKapYusNVXy6D6Fbpv
zlnVD5I/YpR/Cuc/+sUBtLY7GXnDGijMWsz5R6zftqujipi9iDk4J9utOuECh7CepUaOkltlovHh
MgNUqyNj2IxEEHN6+rErLkjKir7wZfPnf2cLcw7ZlxTa0eLmxGMYlWaIEawxQAmv795ruljWHp9T
LkaKOES7z2IBbxQUmGcIjW5JDe4dgDba+GGgGLoxlIdHjeL2j75FhDkZ6M0QV95Lz8HxXUVrC7jD
i2X/4yfrdQ/+2nFaMc+G3VNss/7WMafDWguYpKzNABZ4RWWvSKGC0w5THOtuljxOV+tg9iw+pqcP
xBiPux8rc/V9UvNxGcOQsBsVy+VF6I9IboBHyHl50sWxDBHt/rn6v41/AzcPUnXJ7m11m3nvf38x
d2WoNAN6fFSdey6PixXKuuUzxt/g0nB3w2xUKbs07kdXC21WiBVhexaJ9BDbu9+OmGPlPQs2Hnpd
trpSCipXMZZn2f2Z3ZhIJNtnYYuAo2DSQ+tYa7BVrBK2jLCve+iTZz9s/9Y8LTDRkNeJyn/P/HCn
SjuwVsyTslubm4247RwrJemmWF4giZJZEx+NKowIGhFfaL1sfXGnFbzq8cFrxX5q+tNC6D9W6ueC
tEb+45EvnjlAfpfpYqrI6/J7EvYf5v8OCnavAdc3ju493vMeJeY8ABartZanciljV1PyQ3C2KlxX
CmApJ1QI9SVjpJb5r7+GwzhIrMxZjGlG9+X++OeJTy2nRU1BXMrrGLROqgR8o2en3cTd4s1JDILJ
rHYWX8RgmvkJcagjlnah+w+P/bc94LiC1L/ZLqDA7/s0+zvM2CBM7aS03qt2skoQlxqB6hUFuUSu
Is6A8bcdVjUjYeuaLFpV6GGXcYL9tXvXZkeL7hfAYyhRcgOPBBNupSLdFpDn/WT98DMeU/AP5x00
RF4cOL50xU49BVki84C5LOZeSqahk5Q9zuMkQB5c+7UVvbmc1PydXeGcHwg0sK+/LLgdCQtzERi0
86BINIhBmKSg2cGooybyHUOn2EyNHxq/9Zf7Fn0mWOEDDBlorZ0z9LGwK4b6hNaG4nbWoY+EkFaX
Tgwb0zxSy49+aiFsaMjqmv2ajOQy/QbQO8Xargu35McjtEcoWHv7FaLknnoNTTcxk6KNqrjHoJnu
8D/LdvXocg+llI7xFzrFUUTXZ78ZV+pMVbThaWMc0m/oPjwBIARKOnw1MV2BECDYJfmA7WVLInA2
9QSu9uN4TD1Uf5s9y20/IOGfuQ17HtTXEbV7Pm4lJUAiYzK26o7WdYjwUeU3JsovD73Ur2my1G78
lyj/PN7CQZiQWIYwOiHA2AWAS9DZ0MsoUCw33aSFn8G+PnGH/G915XP488uZbEevuk/JY+ibvLOO
jYpbgQMsTrmQK+1E9tM5kkZudYjquwoNWxTSoc/dLmHJuOj6KJQ/ly1JoekCgUlzUFq/zgkxp3eK
AWOTDkIIouBzUynRXJHAgo+NqmV+KmFmmaK4xSvvKjd/bixbExplO+B4OYOsz+SLGf3pnu93cJAx
PjfSjmBqOw55LQd+8WGtt0qP3CnA7uvkHHBg4z2JUvzT3pGGrESGGM6H3HOQxRGiCtS5oIzxjqNs
lHuy6QlkPykrOBQ1Ixt559CFo9+m9JXIhEXG1PLu+9PCfdO3ybhvRownOaf5ac7mpkrZqb+EvDFm
f1o8gaQlK19BIlKbyWfQ470pidxPyRPSs25JtOEtM6hFVuKiYKRa69MNOawQNTwk+rR0aRPrqIus
wu83wGBX78BSj5UxFkL4eXDOoJF3j7Ni1GJjUbjpAFYkAHftWu07wwSdGPjfFH6YNBL9KVUARAfR
owlir+LeG+TcQ+GN+SlgrDM7Nd/+Rha/f7ior6OYqwHOHsFhD1OmaCtpImBYDbo/fotu8vyUF0ox
AjrT6d3lSZUPWzYwvjISdw26s75F3JlTZmnaLfA6Aq7pdtrE38r8M3fntaZMqAvVlDVo1nZ5ks6/
dXdUYgyVlmSdP8m3gmn8dyTTWLBUz9cP6zPsxlENB6RrkS41clWbzMhRIo5XefGO4TTblvd4HUat
ocgKDGORGldbkaar+Vd5WJZpbJXuQAH3l4TyoveJrEnriTj0tVnEPG4pc0VoTP9IWmXHUasGd8eO
YSLcYsrQjiEfxTOovv49H2OwWMNdusaMF4MdPQvc3hew3/Qmq+7h0FcqJCjZr1o2v5J7zsvlb/tp
P5qAyPpR/XAXnl3JZT0e3UwQUCEDhm+qFWG8HtNAe46ozJL5JSv/MyNOitnZkK6Z8ZOIVCJfMLYz
rB+S2sQr4Hjr8yjIiLyuxETYIwaArsVqqeW3YJpYYlEVLSjBfzKQe6wTuRzm62+ZMsE82ik+102z
NA8blOpE0Ef/tNxp7UsnSTzfxKv5/lsGIkchqjwyizVBbrLjP9S2scQ5NAyVkTJmglZFMaXytaxb
L7iWKDhnIKNXUszuMgyy35C7Tpqf/fPuHGMrqnR4BQVYzmmRCKTG+NZlPmnRvd3112NSxKyRoQa5
ktu3JYeeJhhS0mH+Cgas3Ot4TqMOuffvto1+ujiWu4dnfemcM2qpHo+55fq3L/E5BKTzaKXnE8We
RP+XdQYKB62zDE3oYcAd9Y4rdtk4Y+HvjmgCwWqubeVkceNMIOwXOUSwgHGRnNlpqpvv69vJxhrg
0jAS/g2E9VpoowC6t4cRR6T61PY7k/9TMHnTsnA8wFv4kukHDWt+PCyF/TiG5UwDV6ZbXQ4O5KkN
VWz1f7o4bj4boj3nHbQGnggk7Xp9X6WUb1OspJbQKmnm+CbeCuHWzSJVB6xIgohl6rb8/9ZTsZZ5
yLnMmj8A/z2ymHnaP1u/MpabOJ/iXSWv4zAOPnGs8vD/Sg+r/Qx7hp/sKZh6NwcbV6CUKDB1a2cV
MdtnLA6z7yOfVf6pP2ti6VArFqw5q0nzjXk+AGhCyocB8f61By+Qfv6jSQUSDun2Rw8ANb5edZ5m
JWIgCyPXwF3TzoQWOKoOyFODMQESfwBmV1oOyNRVdYFDXNAoTGWoRBaeiOcB0mkaj4LpJ7MwT5Bg
HeEVVheLFjETRDQIkhJuYj3aPz6dlKkpbKEcqV7N4oDYVNsShXQpD6BkCzp3uePyQfURdNOMK0UR
FBMczn5TIajkKD9z0WpNNWjOwTAyi2wrTE0NkCJHRMs6O2JzgqpXk9AzmjSn9vmjWMEl2qTCV5ZQ
PzGRsnMiRERsCHwQwGbKQS5QkJol4gFlsIaLYjnetWF5IeVNFqP9tLdyze96Nqm4JCAOgR973ZA6
B0XloEGzmIxSRxtS3SIO/ltcoNcV2QnrWOC8LDaUfwuE5jdFps77BGzRflxyz4ESRC8cxMLBu7n8
SuVT+XzGKAVKtc80zisq9w44JYMwoi6r7cGgoatIJKYNhxN/HryXOx40ISx8XfctbLeYh5gbA9ek
d5TJtT3CXaHT8BfSXpNZww+4CFxN8VcPQEXTyf6sU3inJkKcYIyazaRX8LU+0pJlZ4dA1f5/gikR
ueSPr77Cd4MFcmde1ng0emY28rz4GMKt8HxqSvHSba6KGG5f3pB9Rp675thO7Ca4d/2QGyQn0hcg
TrKCgIz5mrMslYQ97s3eJroV+PCf9ipq0lemQYuv1/wagIxHlaholgNtLYOsPNCNw62eYcAuST2i
ivWZJGn98+cLN6BRzcz+QgJm3Zpe+z84hEtz2MUZvPci4p40i+fOL/1iSBvf7zsYFtX3qsMy2sfR
wBAmhM1JeRuYX3ktoUbH/opyprOuUpZP7XMmwRk5lNKMDu6Nck1kz1M8uRtruTM4T5Txoq6gxiuW
T3hvkxYOnHB7hv4ZFCUXDdutmsePY1HE4ZzE9SIM5llMyASDkXW4nCyq9cADkZvkdnbeXY1PIj0k
TgkXsy3TfydmuAoWmJa6Bmyc/Zmgetb0UCJLN9nwWIVVNRpSDjmCSVYFn5zgbuYuYLC9cg3l10qK
O+oLqR6ywse0oc/9L+KvC4/LxMZpL5kq/rmNPjJovwWwQ2l7UYQ0WFbnNLFOnxHYnCf1B1z6wSKp
pzt2gZafpjp8PUGyum+0Sy8hgCZxRw9YrxSbpRREDOfcvelwWhUSLS/2dvNWT5CuR+ClVOQNHYPz
CDPbfT6llLTvuehtxvMlnSViPtVkRbAbl7BXpH7FpNRy0oyVPbzvufc3/qFs5Ny0bueq9vj4jEcj
VzbPURAVqz2xTV1HUxURvDfqxcF6y8HJCWXY/9KmoAecRqsJO/bR6RFSmff+yPb8tKSRf6XmErjE
HhVd/5AJxNcc6S2NsYnqesCXM7+Wh2Q923cyTEkScucwTKLg0OJ4Nx6Xn7yrQls7wS8xdKi0Yzqq
u9930PQe4wiFgMlSlzRflns4v9eTuqC9+lb8R8c2F+4Q2yIQJ3zlfMkwjaXRCZIdwS0NodhI6/m6
czEKWNa3bmFjkP2cwYOBmxBG4b4GriaisVZAz4HSx65t/Xno/hqoEeLY71Mf1+XZ1QCvu9PNx2hY
tMqSdldRTCzkdzlLZ+Oa0GCPr09zKkuxlr+mMDrrmzzG2GYpoLtMIqwvc3SUbHnNbeM2TefN/L8Y
16kIGbzDQEz0Q9PLE1iALJLC5/wgXG2jH2UW7AIqKGCnosNmjcrrKMkVMCrZHpVdkRQN6v22CMn3
5jOKoTf74qWcglkzsb6yp5EgUxNY9H8SSIT+o/qWBs65LWwEIT7nnRBtLmYoGI2nKhjDMansjRX1
JEL3M3Bg9PzauxOjyyixF2yXUTRm6z9D79Rf64bLTdCSTNFAe0BWd7z7RDdrQprqr08L2W7SEcSG
zYgWMt0nkPGhFxZYJ7d5tNHBMQdnRdNU9Swgi+xPF0qqp7gY0DhpTnh/eALbRTMR9ITNwxdis3A0
Rjd6KCIquy4hpO5DymRm59vP3SnbL+y9QL59lZPLnebznUUC9MQbFVrZer1ZasGxlojI92Qshfb7
HJr4G8oEadR160SpX4wyOkqUm5GIElnjDcuymyr6mcQ7Wu9EpG5wYpobOjWAttF18/N9NHxIldSo
m5UviTzDScuGp+DQNalgJbvXDMI54kygG1XSQmU0UBOas/SKUv1EZsVqscMH+guyFJ8TwlQMEuaX
m8KiCnnNI72GvwcPHsVxtulBxZFuTYJ6qO+khCVmpEyKou7ZaYXizpb0VLQ49NSvtHXahI0MMvoQ
sKamvwZwHN5WKOm1E144HJWZNshvshuFYLvdsiYL2XJyYzjNLG2U2Uas9N5leedymAg76xpesl25
hkVSEu/vvqojPUeFySbH1Smp6hfibco517oJWcYvaZRyuF3axafqdmNcpAfPriPxQ0Tm0vV3o+tt
NaL8H2Y4mtwzTyNyzVU9NqUGbOL8ydsuXdKQW9p684CaO/Mlky6LaMK+vncObBZr3XNi9EIwYcgm
c/+UnvSsb1pqj6D+mjQTqulCjFS+sOABOIbIaYu0ymfBQw3JhpEsWcZ5q+DPfNWFw55kyt/xesAL
B9/fvBhv/5K348XUcgR8DuLy4wOf3X1V0CASSJ5/GWcG02dBQiLiDfRncgL8Afk3AN/5w5nsS+BF
2e5L693/GyeCpzRgi2HaaD2JI4nUu9kjaRdcoyA2nO0VI4C5qnykV3OWItE7vay0r1qloVPMqFLM
zAttRR7uq8uQ52w1b0pS0QyNgpMvcjF1qv2I+mP1VWjniB1Y9b97ZHTbA/GgeUQBkE1EdxP21Gzp
fybvaFwrg0dc9Ak0QdXnZCwqKSRKDwI37xsUIQpdEFppEyqDZLKvZ++RCx6nnO0m8Yq1hwP2mDvG
gy4Kt4Lwe9XxhD2trNNflhA01JD0qEdE2+pVYWMFSwKUT9WA0zenvhkUJuPRh+BwFaz4yFLxdEbf
iKO2kjZX9Pq6cxSPPtbQmFb5/qGjnKpaUN1Da7zfri5RxOVk1GCE5yArEsWhHVloPgOVUhIU/5rA
pyVTvB7+/c5UI97nxu4FD11/bJhYUCOOARk+vE9Hpox61ACLca2GPDK1a/Do7jstN0yg7YwYchl9
GntCfCMJw3D9qUNYMUQVL4dm6kYMY5ClvnNIUdsF9uK8P96u3KwoRj6luXZpiOYFW4Y9BcdSYRkn
5ELSeErQ/DiHAkRUfDBo534ZpSBsv0yRc5O6i0MsJZoOf7ooD5Fh2HB/La8zpQzEwzvd0uvYGozs
1OEsVHWZOh+En5wwGDqvcvY5JpH2xzIF2iH7scQL5h9dQPAbFE2huzFbzXEM9X7goT1EBEQTHwl8
XbIJ/D5X+a2G1Bc+QqIC2oF7FGPl40LmrKSmDE4Zv0YMXEl4pc6gbZChGbj5idjGEKSGhvfLMsZR
juQ507oz+JkVkMPaB+moqlaneWWUb1Y/NPDeh014mWQ7Rh6ATfLMXTeozAAuirFr1ghshHEOjvXT
HwaEUbb4xCyb92Ozsdp7EVS0Czg2l1iCv2K8wsTU7emRAu9AFg74Dc2AUao2WrwFClO5Eq1uTdsA
zzPP9fYvLzLt43OnnCY0EO9GvOcuNFMrOGYn5GweaCOR3Ig+YBe0ci2GAqIiwWqKz+pOofjGyE7I
ZIiKF+CKc/1Qnn5wxHjoOT4KbFulI71W3GhGdMxXQg+/pHDEM+R3jSvUjAkeJzscpBV1xlRdJmll
fC6nnKN3FsAqDP2DpDhMpenoMwI/+4kN9Qb8FJBVRzbPhrgeBb6HGCtYIGhg3c+ArOWUKmA5MEvi
UEkExiGeF5VlvzWsiocIwgFBSU7gjZoeR8Wy2uXbWGaPxV3nErLDvbtLkLBx44rjjgCO3GbV154a
0/4CbHbKhxZFxLAXxyS4UJbVtA0I7lV7iCoC6loQOATiAgjogbDrJ9zGWBsmcEzd1gnqpvd/AlSu
lTLnzWQYdG42IGo2gsPMhIpS3EQpgSOVENxrnMBo7WPK0HkYaPP0sOqCaxbJQAOpjUbNhknonf0n
TbmNYTLPQq4EioyzyPTuEDa2esCmuNrBX2D459eyNx0WmV9Er5b2zXO0LibDMXT/mqpIFLCLMfVg
FAaaWbqvM5OuNYx1G0uq89ebAnvsu4XxBPI9q/qvJOy5K07hjv7mmZLbbjk8Ap91sbqvqxddrSZO
bLH7D4kN1htiWQRZfri3ToqPAdhDnYge83JdDf9/z5PaSyGKuWb6WpfzjnKuh6P8V+z7SsMHsBJC
e4lmOVq+gtZnLL+tVi87xoTUeOg3/CUajaVQqvTbJPnltvZjKlaArss0NtwKmgLD3KAYtdUzgHU6
LZOJRQz1v+7zAfuP1UYzVpyCEbkbnCyok7XMUfdwfjNYWd4mhfFPwbxODXJlpTd1Gs8ki7n+1WhV
hAHpigPJYsF9t6UsHXDKeu17JO72hsKx6fkuGYXRj78VtvcuvQjwcgzqyT7wxNbedqcANlEgf3tg
JbfPHCpt4eDFzppKH3VpTq4Ek+wSIOgo27YZ1oJT5NtWkn0TsqjQWi3ld9rjBM3u1E5bjujY3P+C
4kwyIYrKVp1+d276mkqiZEm4jODSa+fNeHkY853zE/xTtKvl6xOqmM+MY3+x0ysKqDiOlLbIYL9T
9mgChjzvclpSO72rKzDn7PSeNWCJIANiKPpyodIvQZk8lzvM0GA7AVIgLN1432+rHSyi/RAO5K2U
iGjANx8IMx591ELsCxlYqMIUKeeWpyea6W2l8gpXuqOrP1Q0U5+4vDXi0HkEwJMM31fvNX4JCTwc
8TneLo1ThNMxCoRQFRoHDSQGx+oYCuMCZkGEzo0jItey2dDf4fr0Yor614Md0JYuC2wIVRv4ZPnq
C9pla9VCzJTjwYBVf8OHHma0CgH3zsUFvFiQ27zhTreSlnhK4zCBEnV15pas5+WjklL5o/XAlQbG
z/ClOyLFoijcyaLXt15cU2HrVggDvq2Q241Vab7KXSjEhANZyzmIzXpYkpOkM/VYfFfFDu54+3wn
D0WYeLv50lJ0i0K4wBJyx3vLSFiwrqTJTXng4pjbCM7POcIRMwYsXWdpsmwxQIqfP7jxItaI6nUb
kXprZCMnKHSoT+9HDLvJXYtXl8cWyqPPwKNesInWqBVardQst1ynBZSXnqYFE5uHWn82HWhZGx41
q4TPw7NNe1YJSURuP7Brs9djLktHKo2J0Cd/zdewERb5v3tXdo0/izuZzo9ZPmkF6X1pJGWH+9H9
ZlQNksH7ZTgmAEQnykxl2l4nUQ5mwS2dgIBRyVduiq4M0ulYQGBU/Ku+KG+ib0Z2WkQ0X/iN2pAr
qiGY/9obh2RaUQscxZu7b3EO2dCKGfkPYFv39SkYOMZ6QFiBONxS1c7NfURc+OYIoG6aXg0KY4ga
job2LFR8SEke3bEG52TYf0YDDAvo6HwVnw03BZyR8Wo5jJGQhUP7Laq42UuwFd57MpE14zVmUN6b
O/Sr3DZsBGMccwlOplD7URU8OtZW7gy/BIu9jbrrP6wSZEr3ctr461qRNUtyIu8u3b+fUW0GMh4+
1rUO7LRShlfLGDvSsflzhTAQ/wq7QPOErT+6hD8xMBntZvTvlxFQ+qOrdiriXOJlRZrobKfFhhv7
bNXpSoezOMtsZ73kG2om8nqoERL9EdtWjaEjVEL396+11dlojnE6l4SNl/QkfD4mD2Qiw681D99s
N/mM/mEI+Oz+FluVuLCT2wuYtCtfjK75X1Vym4Mwjn2sR+Gg9hc+M6Rt1pXpEN410x3k4EuaeDFq
2dgpramNCMNoTvbHwin17FWpyhpb9Fw+rDheXKTZdjAqs8cYBkDPj9GRRkPQgJQt0n2TQ94LXWPV
FrsRxvfXmBMJnX9uOK1t/StADPKzsosye+lUmb4Ec1liz+LZ5F0l+0dTTE6N7HPMjcHTX+kiHUsy
9oLw7sE6z0QGuT3sFCklvqr3b5ZIvwRHQUf7sn5tR4eygygNDUiTviokHLEYEQFS+IstmiGlCvth
jtdyOtjweGLZ2fHGYqygPOn4uTGOc6iidkhfwofx7hewLeWf91uOwqCAIXaXFPaVGIqiRf5W0D1V
ft+t6eicOtVMxNZfS31m2WlqYT2BTDYQtUL6KOO1/NVdjF2D5o/a3z7ns57jCQce7jQ8cZV1bDR7
10MPZGQboPWK3c+CY+oNuADSF1vQH+vKNCJHDIPo5nR+uo6smsiyGOkNWEIEt2ORW9lMtWz2uz4Z
qbbg6jSuA1PKbcJIobcADdRQ/VTTiyQW/q9Qgy3f/bNxJW335ZdywpxqZucKYIAt5s7Q8J+vsTcr
2UePuvPISJiyOrogvOc0dPZb4NMtfk4edW4+pah+vcyk30EKzaSIdAP9ErfPPO/Y2FaOFOSFba5l
+igXiBlTpzZS8Mr1GfATHguPPlz+Nlewcq7V4tcIz7LaRLXZBWA4sUUes0Hu1CPMWLmIvkgGl6aL
91tbPCKrd3We4oYHR2rK+RZIRy6Df0h/YVIkCcgZ+kvP2oFI2BuiSwClOlDUoLHViQHnvwrsTMD1
iyQbFchQcFH8Y7QmjVqYj8O/bTi5AIarf7e7sESs85mRvSFPHAtUGX5cZ2VPJ2seLHYllquio4B6
Ss8vxUMhOlEvx2UdZXBNrrhTZZiFkONKtkDXOe4KveXbs3K1i7ByrlqtW86VehecDe/P+6fpeQZK
IgDcTGRV3ih+Q/DrLtDbwrcgxQuRnjH3mbUKF5EmE54tiX2HEElN0uWnNzIZY9ePyN4ZWqe/AdlN
4AKyF8m/LywlF+l51erRa58zrUBHPeRZuyYLY3pBccxljviD1xCs2j9LzNpB0och2UNvfsoFZHp2
E+bdSo2Wp2LJdHNHfrTWJrhE6Q8OGkTzo8sYKpzatXUO0TZ+jBVBRepqVcXROpcMZjhsZGPBJO2W
AfhXRrLF8uhzT/lWAMb7pEKAKiNBw3uI/PQnMrIeZGqO+oF3p2DOIHeG1Eusjvvi10r0/6D/VQ9I
K+QgRoKey/pA3sKQypFmbn1jJVPjqvBv0d8f9kkcttOFCXMkOdu6DtwZXt15rdZ+uoxRjjhdS+X/
hTdN1yWvsq9l5JN0AJIRF5N9Qcugvgl8imx9qElBN4qgmBE1aBP5UWydlcY0cjbPbggkIDCqR+XS
Nj7qcU/UzBfxppLUVtIncsp53tyPcJfYVwFk+qxZmGARMvfL/kM4egsvJ2uwNuLur/97+YHjfR9r
U3D6QJsqdCWy29W1qgRl5wiJy3YQwThEi4xv2YCx6OOkspTi5jrEJZHm6gxV2XvbkU4Cw2iGB9Jm
zrE+xI89M3tGaqaT3HjAbISfBy5dR7xqEMRj+VL6+BkfnJ0cMxdnU8QG3+S4uEi2mAdmSV86DO/k
iMELutGQezapIIpoMqZvKj9Pk1Yxsu7gW5hFuNFVzntPDtGS1YzA/nUpnWVGRQykyJhyH23lXqcW
qgm7fpJn3/NMHQgTWxPeg5cSmmnWyP0DshAJa3PNnQZ+IWJtASYyWfYqW8OO6q7/MFYyf5OqSDcN
SF8OcdEQtnUHQcPNsKWgPFe2w5jculC5DBgOuBV4U12gNPuk+Zw8l/Zlu2PSIr29xSCC/Vol2r56
EjNJRAxE4FL58kFwJyQ/Yo7vgVyDa+i1yG5tz9DruSOebtzwUXLtiFQ7xLQyw+ZOeLSCpUc9Yxxm
36n4EtzAstMTrIni3CC74wKniDPUXzYyQbHfwtiPeOSld48J/BoMz7/IGl/KTkMoCyGH6e0+ZoFf
tD8Dwi1Gl8slYbRV6bdeHav8tc4A+G+CZa+P7dpV/bhJGR10tAFSBlMpXS0TPSSKk7tjcqqkc9Ce
kApIY/Hm+3jix2C5gVVXqpJ7iXDOjD43EdBXAe4V3WdffQzG7xxrOmN2KxTR4dMi+bMTxGilbFOe
nU7F2tsQjkcJa1+LLFWAX7k+WQ4H0GCrq+0m1EdHWUO+m49pUbXwiLxSZGmHFpTM0IwC63b/kUkQ
4e8Dk5mPgjM3RYzedIPkI0sjTJaQzgxZYsfjvIpcQREcTrI8dUK8EsCI54UnueAiaD32au/u4uc7
wphLWZ3NrPZ0/TkgHFr/47dABRxpijQHzkMkP6fu+CuBTIN0B1RIiYWvX692EOKDSil/YtJsXgCo
Aat98Xzovm+e7k4xej54WQ0Hr8E/3CH486HeKdlXygBG1Xh2V4icW8l+jFmvcmOPP+rB6sNVRwvY
cQ10sHhRP8Lkf40+3V+4uD4kvaPC5JszLnTO5TRlQtHcHJ6weA9xMsiekX6eDdK2AmIfJ4YgEcXf
4vgfQKRNMyWY5ZniTVGXLuyGaDpCxUMOBBMf4q9cVK/u8s1mFEbBfh1B61qX0LrZVdC3wxiUVzKk
HdDJel8RMehgVGBouk8w1C4AvD5COPgXDPE0RSvW03SUpR6is1kBWC/6mFY0DfNrmxk8u1P38eU6
ymqgKseO9GDuh+E2qyETANsPZzWqBldPF48XqYbgg2VqC3P/nhjlGQnleN0EwM8cMqVCP2nfbbeR
Xt0AbpE9FAGQnfjM8RT7n0TvCcCzvp8C3TtnnrIrf22ConF+QaVfO1nPhPccSacZGakvFAh8AiRD
BIxhDNYeCH9fqXyRPXzQcKqDt2d6u9eovNgUT+ddbv0YzPgLRycoOKNaVMy1OwbgjqRW5RD66ZQD
nFveJxvCaMW0jMNA3AGLAsy31FL0CMBm/jmYPxJjPmZam1kFx3Utay8SgerLjfnczWcMh63K1Fqk
0Pnsb6r28fpzTwW7yVZyx/Abb3aGrV8ToxDMsMqLPO0h208T0YG/ruyiTJxc9e3R9u9uNtkqQb27
41tmpvNLZsh4blhVsU/0aKNnfWb3lGBsZaVHnDb8XJbdO+QJ1jrkaNSvRyWR+YUS2DBbOEaWBe6k
LwZYesjxPrhCOkeevtzPkmmNY9/iomvRGtS9RywuurUguEK1MUe8mvFdhSd8joHbIYhOQGvVzhQ8
aXmL4xrobsRJ9XAZx9sqPL4fxJeb259pId7GgzA6g4yh08kzSQAHwOejc3AY9F6A92d39DeuyXBm
Z9fxOmahX6dvsDWqnnEQccVk4AfjDmJugQRTMr4bcKSpaW/nkzveKBbfXb3+XBfebuRNC+D2YAsS
T5evkgVlRImpudaR2xPfhqlk30EYUjlfxvVqCTkhMYyxvFUFR1/bPnlf8/zXMp4qtHW6nHYm+kaV
buW5lvagblRONhBoZo1Vb1dukO002octuqauhbpxHS4aY5wZUPC6MNIkTrDrE9bCMgF6bN5G2G3s
gfg1zksRTyENGhjlYCL+Q7ruUiDFxAmMblSW93DIX3XxZNW/mXI+pZ03cA9I6j++wCiLbCdH0Wtt
srTN/T7c9OgoWfhM26v8eymTwojmbab+k95lIJVjBbVd2SJH1p8o3ZoAh8TvALcUBjbloKtWAfGv
jOvGMPAb3amnrcjyehZh9jaVcJSu4JD0IDUKLNO2j5gXsXv3ThDVseDh7+MRUh+JtYWRErkOFxte
l/kHjnHwLDG0CuUgNKQFLu73nGplTDA3RjY7X1yXI+aBX1PpY8BK2X8TqEfzXV7K5qbjfLmTdEMj
liKC21wZSGzFzcus8I6Yx+A2mAWjocNarwBWfuUFFGNtyENI6t8TFcrR7MlF8jX9KEp9W4iTuKH2
LY/Ahabaxw82M66jLrbbFNq9rw6wLF8yBKAmFtPUFkoz0AA6h+R/WbNvEms5WIQXfbL4t+BMdna+
MyMBwBgmdQmiTT505N1rcVjQN87nkfvf4xQTdehNWh8fxbhJpE4kpAJy6LVkfN4D3xjzTsDwfZ1s
qCPZdYumfrwtDHFMMaILRJBbreVUFySA0lOWa7BqhRMcPU8BCBcL6iWgf7oyFIuIO4Vmh/IjzVJT
9xIr8JLsD1dyB5boVT4HaetRG24D6kwVBasgT64Tk/LvakGm4DloZYtrISVnkEapxQkkJR6hyAe9
avZEM50vx0ZO1aLgo11JfUrKRA/lhew7J3u0R6TRUCRw6KJVqmZpwnsCNwbiENi0jbRJlllkUqTM
6N708pij7WSeL9FrdLJnc6RyFxGHD2O7zvhVkh6Q/gFZgGoztU/vFdpCTIdVkeEECpYVLqiQxbs6
9WowXZvni9ebN6QS4coR3TkQJeyL8cVz2rQXGVAjL2Rrfdn3Svqb7ywdOmucy+2mKRNuGETMCOR8
svdYh9A4YYQMkhfExsrSk9KWXQv1+Da6SRNhnzWQiMqbi9kKteqFzgGTDOemTD/pI5YjvYGtrwMd
IfzoxiRVx/jZCsND1b/u68oksmM/3O+xswvQ7+HVMcaK9OyQXBnxHFqzpJuS3cn20ey7lGxG6qJQ
lt28Q+/bVH55+nTHwutnoPY0XvsD8FVyTHnmFCOJAqrNkYV07svBNdJQ1md/VvwagITNtd18XNPx
9I3dnXc6q/qYnQXFI8H/iYbkPYuuDgqq8SlPYX1fjIVYbsxKWvWmSWh0N34Ay7lrJo9xNKKFjLyZ
rMXd32dMib1j0pp+kObTEcJL0i7kc3Y2TYAjAxAhDQc9+Q4PITsAeA8iKRmQzh24jXCBiY90OBY8
k1wTS7WPT1do4UFEcVPuZCZc7vNeyT9ClIOTmr0LAiMNy6umuHs/w7u5eUg206X+4uB0F5/Zqc4f
018DywL53rFMrgLUbTH+U4bgY1y7ii2KIItarG/gl/QRBQSQTOKtIbJ2Xsav53BzDxXTgK6aBWLg
0N6GV595coZB8nA8tFjYOBHHWrFYAyIqR3wKWj86Fig+8+V29TrO111sWSYu1yF++ztgw1M2iyIO
ENCKb+uznE71QxBOWUN3RKqMMntWOfgMmS8TUNIeDRjy4KBPIj40UZDx8RjCxhfhqBM3rAX/IsOO
lAU1tgBjn+V2Ne8XtDY1mSA2LuwCC9iEa9nIng3kQA/OmxdVQivCk3sF78AULXhPERrOxW4C52uD
SHdvWvv6ujFIRosmHbbOrEErMEh9FPteMkYohhZ8+nr+M6FqP79ZJTC9M/ktEpb5V+d+EUUh521f
vRtu5aNFafKlquazJnskhDq63R18L7/HgPmd1LdPnzecpoYpmuwmGP5DJMuWXxFQw9kpNJcJWcjg
1v62xd/lBdt/QnnTugLurf7w78gBBajgC/d7CVwhRZrtZi6TwoFcamw8IVgQdOkWxkbWc4Kpp0fA
9KMqdASYAvV+Ra1NGdM73Cdf4S+AdVu/S9O8e0lrCg4oKKUE/ZdseoNKeCZrNi9V2WaYUkD96P6i
E+83jtNsK59ZGwU6qsNaZyKQI+4gbdyxyOxs2mzRFn4XTxZ4KU6Xa7elcFnGjumlqraps2Yek0K3
vy1IfbE38tjSn4InL0nYwhyk7RT6aJtotD7P0TMvYL9OrsQviXjzk7FnD8rkzVKgpZZ8bisZ5XIB
a6RvtxJ8kAFfZyeuBMQYgzFL0z0FOS9DYSLl/vvxPLEWIzouVUl0kWxqPpCdLo3OYwZB8A/7Xe7e
ElN95zsa5o9Za2TP65v736tJWQv54qAcdtpeIj3GQ2wkvSyOlg4rUDEtClwe2XXcCoRf/K1GZClR
5cfu8N3rRNUhWdHsEW2SCfeEJ6Q5ZFrX6REyxwy3ONSb2M055rAhz7ULpt7CIKIn5zrUf5tHROkr
w9vSGSHGKbWnRdY48bLRRODmKtdBk5FiWH2K/MQiH+Ew7F9mJ40+NVcomgbJCM3slL+fNxpJfsyz
L7wSOF1wg/j3FCqcp0NZA8d3lGN3HnEEYRoJR+3wAZGQnoa16Xtlg2CdKn74shBGte5BDkZqueJl
dYT0H979b/Qc5X066oBW3Vtekmjlzn02jBdp8iGH+V6eNZT2ZG8UAa2kngkhp757DFj42vqfCG7p
VbuYK474X5mjDvb3sc/DdKNnY7rSi6im2ygTkYFBJVkxw494y9BuXZwoeXV1LwNc8r8x3mp14OMV
THXSKlPzRJfXAu4IYKNdw5d/wncDLzLrgAwrXwx1CmJks+AEHCH21cvIlv4c88tMT9Ifkj6MAIDk
HlWyKMHzZBrIn9pkPMJ/uiyMie2SyWSTcO/3qfxxsSv3g6f980w3Eu+pLkR1qi+FUffieQAu8dNC
3SUHYMaJv+Wy1nyUPOGWDe9sL3Q2jVVa/DHMngfJUjMYefalYUb9kqR9HztbIM1ISBToJOHW5V9a
PnGiNaLU3RT2KC3YwPVW8u040jhI5IIZowNFxv/FNb8DlM3aismG1H+QaUy18u/yOj5p1956d5/y
AGBwj4gei39uyb4JZ0jz2Bi5xk9ouSyZ16w3A5+M6eaEp6UeTv6+0mj3ElUiL5344GhfB7H3k6Jw
SwCY3m7cpO2heCCFTiYpw1t5Dol52xv4Ei1gG/DHOhTgUAkRlHGi1UG+iPKCI2XYsW0e1VreVAbU
qQWMZNZH5ko/4jB2qDJVC/pb9W3jkxheRBk5oxg3zDKysUZyeoDe7WG85FKH9NRSYsaH7WAZqLQ9
XkUAC85kwcU1snG7Q0h0eyJ3xLa7hHGWP01AGk9ckQfMFLxD6g+eX6wZHRZrfpDNKbX/DuITdL61
eAZLXvZQn30bXTASBGHf8U4D241znKKlFINKg7Oj5ypuqWnUw8YySfMOqdR9Yd1mJYidDY7pNrg+
rTtVs8ZEPnVjKHOHI33V9URgQPEXwnZDNraBetEfN/e+MxFLxcyVPltnWkwT6SaSVDmJnDByMlBw
MUWvB9Kbv/QP5AvgCkzweeJ3jMQGZSQ/NsP2zfL+JtpPEQ6hNoA7ZNsSztV8HLMmV0fUCQcMyKLi
GJ6Aj7aPRGlcmyJbP5h2EwXfTBMWXQBipaUZ4Q/PENgolnYMgJtrDD5hMmroWHnCmtYt1jTfFTgz
hO2JHrs9hvLJiBdbgyknqCcre/InZtdvmORIe3oaQZTKVFIh+5o/a0FR7jpvYD1ax61syEOWw0Sg
qvJysixpBDwnBKAJhfWPPSh8StfscHxB3mimvQJHqnxBd+FZpssQ2fMaVm3zRVHIvKWbbuF3Cv3c
kSz932LfqsZ6fi4B7/E2CH1hc/KcNVdYflFTYWxlrtVmzKstZn0ODVmaZQWjFsNBQcNLUqaVFWSf
DIKv6eBuon4NpH+Q4YTOXa+plDlbZYmBdn09A1hPJSKfOyxMVEuV7jEv1QOHWDd2SRk71GBAZa9Y
0cL8+sCT2yb+nhYFaIzhsIdlKrRRo02a5y/SFx9KRNyqSC3cpyde1l+9i3Ab9AltKUm4hx20GacF
0QiuLJSKpjzFMvsOestguEeDktq+L318lIuXmOshRPZF/Lylqw+94QJNl9OFOtrtYCUvK6+UpHg5
cifbBFoO4Zymuqf1bbikKk6hcYJNviCjVgWcOv/ZAG4+q283NvD4SNtmhz1SvSjHFaDPa1SMwQWJ
G/yDC4sbo+iQXSeHjzkPmvJGRLxOu2AHfw9NVYalkC828hiwEDsumBnO/lHqfjioTLI4xuptJxJf
jLJsrtifmhFQCCJGO/F163GXXIhVeGurp7WU7yFi2h54lMkuewm/RzcIai/FsyLvJ4PffIuy219H
Nt/QnIV6czZ9WNcSNsuAH5cy4qEsmm2bniob1THy/GCLyivmP0ru1VHrquF7sxk/TTK3rJfgM1ym
r9ypSlVizo/Vt3RQKcpWnbOfMXvIne7NmdjlvaDXkkdJvFepoxaIlk3Rev3f+4r+ySFaN2mIJd0q
ckv53r6/vm5qNcZf5aZiucWl3pnyAu+bDcDB+4YB/klOcbkpRQ3a16JwbNz1K++z0fuM5pR2MQyJ
D2yPBJ7w+23KbpNAxFBDPA6JAcLg2Cweyb9N8GjuQIJXfyQZG0kPANRZkmeIydiYvvTsH5sKSBiD
rdk8XGFSjCjpACQYuIBmMsafeI5pbo7qcOi6NTwGmk0CotlL+UpeG678fxCE0R/Nul/h3IC6JuyD
pTtiQyOTXpGAOnTevrVwz2wsXm/t2yJ9IlT6p1AFgZiGJBle0ejXmCAwpLR+JPeOcka+AIQtLfND
fYCeL35LNFtN2MfbOGUeR8bkL+5PYR962TjJ95H58s7kri05CAYSr72+Qxx1TSObzTeGdkO8fE9n
lJ2OOU5WbzP1v0GoYzcdFPTEdErZxP6zSROgJfm9UGTcW82NK7XTzT2BvapdxGvPNCmtJiHhet6V
9nc7ZxBijZ+x0z2ckYmQH+UWypbiXTxLvWvGepJ+hpUqvBfNT1cdP4s6d8bWKEB1XjzuaxwWQPwY
e0/PRyqCvv0ZBdSQrySS6k2cTfI6lYN32e39UIboYFMQyiJA3SUgNZhdNqlgx54NmUviX6CbwDno
QO7Duu7Kc5JcjhGS8yIES0kT4WliAMRGaSyDEEds85kS7x9kqJSY1rPwnp5FYdCmXfti8ITvj2dX
x8fAGS3LPBTB9tOL0C4jLliTX6FdpiO7srozMfDrwC0MlaeWmmOJGAooiQ2CZ/XCeoPFupPBYqjW
WJLW5RE2VwXkqGJZa3G3eIbWmRpLPHadzC/6ZEHPAavRNgRYPtBg4wkoSXVTOLDFQcMHSDvM5AJM
HDDATV2qjh5EOgALMN1wVs6IdV860CMT/3qOcOkB9ST1xBz7c+kXhGVbe3zmRhqshklAyprCwuS0
bmRh9BrzcpLLJoX0VbmLe15ZUaqanUWzbNQRg5yBeMKrhyyxm17j2EYKTOF7uwLZo7G5rmEZqp2r
nweOrLKw2pBfjz/m+DqsdJB9mwhJ9tGXtq4Y31hCrFYbx0Cd1LMXjm624So/jDcMdsCPD1SiwEN+
9sEByBQMv8SQzmG2O5DA2YmZiNfFUy22wlDEawh9mvsjhqStzHYOzFh29jPUPY+v2YqnkbGFM2Uo
c4P4U5byhnb0SvhcSdXJ8+kN+a6tsIc/bhH0VYQw2gE4b4um63YtQJNvm40clSsENJxH5+P68tce
a5QekYUhUR6TTSJRGNvdypgmgSt9TIZ0hNYO9mQgsGKST8opQMKrH7vKv2+4kLo5HceYBCk004Uy
jBxHYbbP35ak5VD1JYPRp6B9JbICfDs27Hbf/Y+f5oEypAULV9IKK/RD8M1GkM72jNfkuvfrOSW6
KRsHpVImTVMbmTO0Rhjo06JDTbmSrFX8FZOCSr6o8sts4XEEK3DzSHe7n2wg2FBBJLA9pS/aaizK
AIGBBOF8/gklEeQI3GTjFIm2pkAtt+1cXExAT2Zf81nYA8AdKTePo0evHWdMmLkl3zexjBTIKypV
agoLU86FG9g9g58LgcUTIwz4GGGbukiLVHAUj/8N2hhDlnBybDwH0shNQx72WCCPxuQbjPrJNgVK
6G+uVu/kj8kuFb7YWdmIvAviT88SHvLiGjUf9dgnPSU2Z8kIqFobS+3IidojvAd3ZOO9H0drohfU
wbAFlzJPcljlMYn/cdbhxWiiKSE1UbjNQuKQGeziKg6x+wv4xNG0Sb+h80njSA6TiXYMEnxahsxa
R1rKh+SgdAuDl99X66UtM0VAudASyEjkEHV0qsJjRzi+pDB2aLsdWXb4r5gUr+Hoe3oot5udfRvQ
labehjif+8fJ2EUxlDl77rWXiePrSplPHKviWJiLqJ3AYYtN+7RDIPNWHksc3ryiDgK1EBkN2UiC
faMy9zbay2y6MV5Ss50IaWwRVCVgR81fOT2cJG63NOCTzphg604iEBw8KBmFnmkyq5ub8/FnwdFD
KNGQqsXdGFQmMJqVl2fw94YIIPRr0mfroCuADDDvHheYs3nQWEMmF/gQ6GJNkqWs3fayOqQpRFM+
E8CeLwWnwqmQH+/B2pPY6j9OlTJcqot6J06ydAYVLZYs7BQ2lKmgfsxCWuH2W0bf+UoMKy2CLxTq
JmwfeQ7CTqJbqmR65isFhEcMMVDRifIKmHvpEVNr4gIAJurWs+ss6ueVcWQovGnHBAwvYUEqfP/I
f0/jeFn5XhQz2rMH59PishSp3P/gDOGITak3J90BBIZSUfHq2szZa5cvGrczmLWIv7Pa2Pb1Ekpe
Z3og4HYW7c/CYTrUBSC51CHPvVTQ3sbcZG5VG7aGPysf+C3AFESWsPCxzyQgUhCm4P8XrI1nOXd/
YMzqw/M8xKcvuCIkMklhtsrkbSlg1zqYR9GeGyMjsO8RihFDgXPb8oZSl9Vgf42h7vC8OegSl/OR
gyVACJrnY/qz+igdID37iCaE+Ml7REXo6NY1iz5fss7NshsVsq35Rt+kPna4N1ebjwA8Cmh9r91w
38iKGBzcKhj+VEDtloxu98pl+S/cVse+60nqKXbKlhTHfqtjCf8W/AEQlx8sbl1TZJPNJ2IrkTup
+JfOWkWFG+Ba/2pL16UIpFlXTQWB8d5oTHtDXIsttu56ueCi2Ptfg471wCOZjl/u9T2NVJSsVU7I
rR63TFCSsmF2DNZyhmT4Kuebvuh2TLFWRkhQjUuCfiFpvf+MOCZaA/6n5B1CkYfFfvF6UaVOWUW3
mNts6gTOcG70x2uCWLFMbVRflCigR8Q2uMf1ggdKBjewHIk8E7A9VSbyx++AAljhDhG1ecRCFw4+
JTVV/Gkxwx7wZ8DkR6ptsaa2RYJR0DNkEyipi0a6/V+IFJgCyumc3kWH70X4TqNIdI/6Ya9qHvVr
z4GBajki2TK6H8F0DwXUOX4qxzg9iM+f4lxJamdjpb/s/DRS5/063E3Xu2R0bjknta5eZQtKbQcD
LKIi8ziHdnUW5123tXDDTAbhj+f1BkHrxu6BPl3rWAjNiAGAZEHwsw2UKV5SIuA7uqNk8yHbuBK4
MX7ENCiCZyRFabMozSOE0O9plM27z6lot+J9NcynlGZ97iZj9m7wbJEHC3yR9VSsgqdxWG3/t4qV
ujyp7Jj0KFKNIQRaRf8XbsN/gPltK6NMbgA2FZ1qw5N1nT0phsdDftW8yMenBybejcWC7+MKy3mY
EoOABsvq8OJNMpY8iLaQhJ2sPLAx4wZDugoIC7reltoT9mdSIXmNyr8FPab5V3QqdsIBQHKGzJnb
30gmrDLHGeWT9gCmhcnwOX2AGI3sRaewIXX7OLCLC6prJfvUIMmcNHueaEnyDnreksbOHUHHRVmp
OsO+ALZEF4+9Fkrh07AF+EgP8XhmntqmPBJlE8pIXqCduEvnEVsQiHl9xglaBQCuSpiL4C8Tr68g
C4VUsIes0gXqY7hPvmNVCIMUIr+gbu1xB6pKJLhVJbq8EOwBmhLYVGM0FYaGrZY9jailV4uyq0WY
uoCpKY0UjnNt7zno/bffnQiEdIoBJmpwXaCR0vx9LxPEHzxZlr7USYakXVgKNnCPWywVd5D4xCxq
EJKI4iJSqe3DnJOYZc2d323fDgBd07DUPQg0SFZHrIIFq876U0IEvJ7R7P/ctSgpwKpUaCvj/PQs
9iD+rdRJHV1XCdH5JQHEwHlJev1/0l+OSwpfMvVutObbEY0AD9drEzv8SC7Zza8e2VpB5y76gkqq
n/Fm4/LfgxjvgxkGQEAtiGMXIL0CjxzaahPxRo7Atoy1OLr8WVhnQs93RmMFNAKeaXr5EvauJbgd
ZODzV9zV9Oz713e8LT/GEFkqvs4SSnUkZTVGIj/Rjhz1/ElvH5Gnntgf+VPwcVhBhU32z3b3zVR2
g3jtJBluBmkC5un3vbpkWmeXJDP9LXxbTHS1m4OPElxvb3cJ/xuccewDyiqEjw98K64X4NBhpUzY
EQpnbA/cJcC7eLBae4FNm4ufUMVNs+CPeS5oXFO7j/aIe5jahw6RJ5dLEWrq+Ucr6tao0oCnAz00
EDtNshH1QWRqcUDJ9Iz82LG7fshknss+E6GzQL4OvRGn1XFN5pS/WbnIGzNPx7x+JXyTivyO47WX
L+Cmc7W7kWcLlCjsyRQo3/txsIFb7TBUNVm2Rwk0PXtBvTGiTLyVKwhIoJ8xAqMRM9s7P69AwlmX
VcKq8rXq7LB+v7AqAhr+YsUAQ6j1guYjsJqzB+oZchcgVoCSDDjck9kzx7jpQLuLKU5piFol1/ae
vijB7csZt+yHwtl1B7IcHIvzBl11hyXalmWkuBbQodUwrmN8lPYAhWeVkliLFism0EXU1bh2gynV
l3epyOr8wCeLmIx+sCJaD2jJe0aRYA6mXyokNiKzoObs5Pp+TlPnxY21TCnp0w4kXm7EYMVngXkO
JYgYdndMnyJUp18ydLer0EtARRXiJvpmthPGuCdAG0denDkmeToA/sBIKaV5zu2z1OhZwqwE+X1D
LVy/rhHwoofo1MIGi46uPRaOopT74qZxgOSQsRuEKXjXDbLByLz43AfGjvR0PI9c1jCJp6nGCM5q
anGOOK714aKp/fEe8wZItcii29sBCOnUO0uP/FsINW5VwApUwUFBvNNg2oP+MIRswFfHKb6F9Ziz
JENDxyqWcQAsBRVN+V1XncAxQl7ANNug6xBlTLJTTooiGGJKUQzvJr1jhxu5B2M4Br7QStZxAZUK
K5UAKq7dFhXpPictVI2qsRi35F/DJ6tYypyqXrTiRgwEwkdGC0GJJVcRCw95XaueMjlj6NOXu9zL
hw04PQZZ2oyZtNPatAE0UUTU+DROwnsDNG2KilePj+fdNwN+rshDjfzUwt4vN7HmKXslHJLBxUIz
A9pDacg2s98posGXNjw2rOLV+Xmuki2l4ePqT3dvdSHy/tbSV+88PLnsL0SOpOt85g5yljAKx98Y
0Ynxbs8N6zmdvCt/UBD6IyTQZ6e2efOg50oH/Didbv86718VtopSRBb9h9jOBfnPNKpg7N8YpJyo
+vKfB0B//nIhQOwLsSm2HGTDbFVojMfbgapB9+71iKeCULqdS4ybrBEnh1ToQ4h3iJhOgHvMDvAD
N29bd3oWQVue2Jg3D6qLFB6Y4Wtd/DrAti3ncAq6bvpvZvpykBAoZmpacz1wmjTrGJftpe0qy2NN
Jgwts/Y5XtvOVPGrW62m49X8ax0PPDQK8LmvePTkqczNI7NGDb1kyZ2jwGj3dzryrWf4mLNr1UqR
S0ehYb54HJ2ibknteBoV998OMsa6GdMnGq/Ryu7/t3RP3gT5rIoL0IxQEMYc9ZD+hRXJtiyEmI8W
WLjeNuOEMGp9+9yTNVI5La7bDNxReco03Xx65ybH2aQjCLlE9LHJ6adbO8qZjy5OKlTOrFoiX+pa
q2PZmHdXsWdxggDq/bvACPJ6mJvpoJCp+3U6OGXqtkO8vdPj2cfzD2F6ao1YSWoxoAWrc3lpOgHs
t3TE+KehtG9HwROjhDQx1IL8mWCgFSm8WsyTQwTyIyfDSO+ONh0CStGEK7HZVZNoyL9QHvC3QpHD
XXwGMcylkAaGK3norPfDchGl/1hg2RuFtzh0E63MxcGqxDUMqXN8ZqN6S/Bdt57EO3+UvI1jRXHf
K3mUTHSJF4K4FX1Cl4/n0oVlBuRCqejHfNsO4ciULTefmKE8VHLUbwMiXENiKB2liC/sTjfVJ0iB
H5Ds8irv0bDNMr5NGAloEQk8JdW2Y75z0yCgQTRSZamUvFe5Cc62WvWFR7LH7BOveAKbO7iyi7Z5
AizqzQoyu9dX2obpGQo+Rq2JT0O9zhAXeAQl6iUkZnx++iNKJiFTxUxxObFkRmYNnAoUg0vATEAX
nQiu4iXZYNlZbnpXerw0dy+oCmxOKw+J6xqHjBQtaq1VgDY8Zf+imZGQzySP29Hh4bBzFu/1Z2W6
ugn1Tc5kI0R5jtrEJmCfdtYtGFukD4BOHWO8H4KSB7V7SMzC+aXAVujEsr97yqR6cVf2NHmLgl+R
Rygi4fv1F3ijYaHj/ZDRyQe++Op8uC82M+063Q9t8dgi+cpmn4CD2g9VsRcLJphrfNOsSwPLnKUy
RGo4u1vvVBBZfeXi5TFtClD9GiZLKzrj5gzDLW2BpyCYMpUIzWd6UjkP1h1DnXhWjEOOJ1cA4ZT5
U7e7nhMJH+UDvUzS/Ddwz6uiVx2XXlT69YRBXEG5C5qGkyAQmeOJePwzsFOQnMOcWx1e3/EDGsix
dh9umItJtl6NFa1B1w9d4mDwonBnFHouTUsACJD3X0dhm/gQ6uCnx/sOg0/eBnfa3Ryqqr05sBP+
fIUwZaWS76yFSjsepFXxTOvIcB3AWVJ69aGsyhGL3AKBkbeGI4K70mlYS2kfdMumq0HA6FBpMr/d
QYUeXr48S0VbO07MjImUaSMC5PyZ/zhH4IYPOxuVgc35YhMtQlBSCMpttADkrJfbjuF5FjJS4dzh
wY8s7iTR/TvwDDApFnEc/PrpGQwusZJlCidUs0BfNaS+i1Cj7yf4wvVEu8CyAyMah+GbpxK6jhq4
fR28nErrMcL8po8HrhpZpg4p67ICH4LGy07xURG7Z81VljJ9y4Q3NRjhhSWdJ3dkDkr3CGurZO2K
ckG717tHfOdoRr5ilfajlXpnj4y/wRLjQ8ZzLd1xGuN9voEB1uhbvtCHvM1AEVX3mDpXWT/quPXz
9CNccQ4hfOAYEa8DW95N2WFNrVGX7ZYzdDjCtks8P0ZnRfUwIw9+t+igSziD9KENPv/K5lmT8icj
pOes9GRSJEOJKUG/rLeoHCbTneCvDFeRRzNoedq4dzBmsgUziIkwbnucMOW27wt2W5IAgHKlgldm
LHd+DZmJ08hG5QcAk7EeqqK/G4VlVxDflETaPU+HZKwic/YNyPLh5O16h0BuBSWNWfF45+WpRmmM
7cuG8Jc+dO1AyYbCcClvc5ET4SW2vrV8FcanZDQahGVXlhUmZz8qxuI5i2o6/cXNDGUHdl8TVWY0
R93euXROPJa6m8spZ+zIgP/2jsWIxKcw7hWL3Bq85askaCZm48DaOdw9Te8sEYC8F03IiUnO1wMM
iNwR/hF2ORLLZ0SHPa1wkv3nPuRlOkFGm7Ox6taMV0/TpXoBBGq3UpxOJm+B+/Pk4wUCN8cF0XKO
rZdUQP5azs8cl8jn+fIszAzKjVcbjWrLwnQHDYAfy4r6hjxnF9xYE02DtE9KntkDLOsHQSi90j/0
l4qUGL/3caaSEaBw90wNY4f3mA6V3j4ucwu0sVpNZ3eZI+3ChO3D/TbJFTmRmnjAyGPAKF8Jo8jP
pPxS9xXErIsim/NjwQkMmmuopE0VDt7RsZ48w3Js91MyDceSDPQRL7iRFXZEr0SrCPYUHUsKe4GW
Szn2jouxuYDh+XEy2GVpfx8NKDQ/TBJGP9RkE7+/KJYR0eEjSorNf6oySOLgsMaqF+MAmo5e20du
Q153PoOviZ6a2dP4Q88Ad+/0b6Qn1o/MFZlPbokSun2B8y0/OOa0MSPsxC5cl8017HF+zYdBMyWJ
NF02bUDfGmS0qyMhTr1cTtKUZ5fXsBbjX5rVDWHv3UiQc8vmx8kukqu4DP4PHyX8OTQ5CQDpIo0d
avpIdA6jBiYm618EQRGBkJgmaN2KRlIgU1HUvJ5aqwxRCjiZ7xhzztNoxLn9kpK6u41QFxYLk5YB
hEVtKEF1xE3Z529XDlyqPLs+Jfw1FSGFqWZMeLB2IPEoA3k9pVbTdzGQ6PQGKEhP/7xMD6i4t1gG
7QJxFQ+qRGqa7n6CoYVuVfpdvpVd8KttT1cVWy2YcULC5Hur3H1KPmMwM49BjLJuGUxXMdXNCl9n
0seNSzwn33ip9BJyG1H2S5Nrobza4OaPKyzGEKOEYuY0kzpZ3DutAzwaoYUYDCvVakgColSEknNx
XSuxgazqy9wEhAY+FVAqakpzpZb7aY+zOB6yXmKY7fRuIKf7Ii6iqWzlc3+114i1Qup9O0O3gP0N
MId93DKMBl9N+ApOx9bxI4AW+nhRswJr4lLpjpAXIxQTUnXdbtWtb7e7XlSagsgChFQ4kjeebaqE
yFNZ9UoS60EwpAdFfS8eOwz+AuZRREI2s9ph500wMOyJrcpBqSNCJBbbRsE8edXmED27GBwh6Tq6
8cTb5EvmwQNvlFnCa7rrIP8aNbS+JtdZ5y1jt7p6FW3G3rnyoKtpoVbJJ26O59FdEvoYtE1F09fN
hOzETHm/v0C+aDw+Zgip7xUh3J2BzlC8e52nBm4lDOhVzrxrYtfVFUmF7i76waKKfkW38Klx+V5T
k7TohBkbGaA8pxNkTDwxGwPx5TmwUx3a3a2yD60n7Vz3TbBt8rtd2E37NzBd5YsHnrnpZH2iVCyS
hiLy/MwjuA1TRtvuWnbVSw3nt7fp+f7Off3ueEiuqfJ1mSEhTMU+JWn2B+GeYz0siSHsgN/QXk40
JWeEaFklQxTyjEQG2FzDcNOEdMhrDh38jfLbYkXg0JkxFrhABxlJO5BCTIKLDhg+SkoURFbjHFoJ
LQEQrgn+I1HgO/1+MA2irN+0DhMB880lUfawNoZtz7pJRO2GGcmVMxRzZP5V6apYzWQN/gPEt4ZJ
IsovmhFOkQf+3SOz4/kU5/2aLPbe9uxe5uI45+W6ltSVhDAsQOa7lOpmgx3acqzCmC9fD0JB7Ije
CweLc8JdUuhvbGEkcTU6I7f6MPG3LfstQBTbskgKlFHhlSk4A3Lcduuc2mNi100y4X1RvuuiqplP
SmY92HKrn1ascAZnEPJdjIRH3UGH1rZLHEjdCUiFi106+NAyxcxKC2H3BmOQBr3mYgB1aPJwzPiM
ZtDtP0KqhYX+8BbAI+N+hyPfi7q1BzJE4biutCI6yYnLzEJetcddpm9sUKbc0Pa2nddOsj2zuR4i
ACCfeP0VsoJnAib+o34xD6Ml0xEAh1mU1/QW1bruVmM+s4km+EQbi2Xg4YpcV61ofRQ53SnVLOul
Ejx7tnZo1hVXLHWLGj9ZZpkZqnQKaq0DtvwzsDo925Po4Ht53H9Dx9iSnIZ6a2Fl4Ng6WfG7yQf4
HcV0nVwExt/Na71Y5o8Ah1eOm19IW9Ty9H1reNBzmFda5zViLevn8IHWvu4vzyueqgRs3D9YU2aZ
aN1H4fERh/ka3JzlqHWzg5AqRugOQYz4Bv3d8vmE67q2aUqXhd0wcgJ2a0Frt5yKhnEVxgPJy7eb
8VLBoHehqFYOUWWNLLSiRo2Au6XjN2EaEQgM9OMDFv19OZKLoqYawgfF3mKKHXfS7wtrJRE83SD0
enauU1PXcRm1TGx+ze43ciDM2SthHHD6eN8j/J6rHlwygoW1Z4cwpXeCo056ZT+oQ0jW38JPkvbu
Z6fyUqLdaWQFcUExoYXgqkjDuGNKo9n5ORewq90BX0okAH2V/G3jexF8RMVmyvcTun7pj4xas2x2
AQL/Z2AMARFXjHw1xf4pnQVGgtKgmDF56xgipB8ZjuiG0T8VYSLgURl3QDFlx/EyfP951yCBcO3j
59RNJAEnxDUA5iDBXxdGCEPoti6bgwcucqE0XrHZdfSxooPKhagTJms5gwWkQu2vmQ6RQcUQHugY
RMyDEMh73kMcOxz1ajTBwnaTq06IAaHEMCLkCDVNvoEJ06N5AdfH9T/cZ/PiCCzYBB7TnFkDSB0F
oqz/XTiZh8p3qcsyP3Xyufvy20ASvNP0vQBLd6/jVzioJRAbKUro49Nb5yDBaRvBSwfixkuLip7Y
8aKjSeJdF4Pyd3IpkWIr10iKYECb5LFF4xgMkJ4mn/LU6w==
`protect end_protected
