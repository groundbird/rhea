`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SBfzr4OG+Kss92GDhB+efubXS5uCzjiib40cGZlEFPDPNT+pOpfhMHbdHG1nbFM9wtj+9CQrtkcD
h/8niKwehQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mt/Lj8iu8VFQwXx95kTY7IBLbVHL9MBZeQUGRd/H+QQFpEC8iEvYdwuls/JnSMmhOJ2iG5c6Aay2
u1AeM+iLROD5Swu4Me+XK0dNgExJRPxxJVAavNlLZ0uhtWo8VYBTjvIPrVm4lD/13tPSa84YIMlb
64IZtXVHxlZ1xtgwhDw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JCLsIFfMYTZz0usUN8rJQKev+ydw+fxgYmK+qep0Wl8QpcdmqbvncpBh7rLw4TELgLWM72+RX+Cu
IWh2h87v3hLIw6LmzAQFs3pjrL/0oB1BXefzEQJeeg/c2TQCWNKiYvOzwmNesJQoo8gxzTjOc2vR
AQzWmuJ1lN1kT7rnF6pB2QdNiQLE24OI+tsuorPg9wUb3tgYLmQMPMt0LVvXWIo7jDuIMeMc/vgY
igu4wk2k3ml5YgtywiuQrDiCJWGH+CgGvip8VcJjDM8KZvl7shMcsH5B19/0FCqZFx4jBCVThVvX
5k0pvmikEwgIRU2DfqHnZ0stWzvXcwTm1ZMPjg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FBNdP+IxBwXtudukAN/KtNbUgLpqhNXYu79lLsOAhlaSkQCJgurztMExZBUZHDvMED9UZio2mu51
WlDl5iYNVX0dfqy4tuChJN95xCdto10XoznCsoayXc5ve3WiekjTQgULj8ldunSD3AAK8twCgP9q
iFHJ+EY9e4UGgCq0Pbc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gsuz/gMQPMDdtXyFHgCwtnMRQ+kML7JVa6S0X0TJd/CnW+9xdzZNfBrWdxHj6SwNwuzJwJzhNOOA
3pM9d+Mi9ZxN3f87dGEigB6Qmi8E2ql7SWoHZsLJK7TjgaSz91SHKvnP5M447Xhu+bJTkJwPdqAN
0twRElEXyfYC4XFxQYiBqsDv2CAc/FE2T0hZ5ZkQXCwudML9MSj0DmEfqMD7YIkHbL+39Anw37eG
fPXi99Lmxn+yqIGLwMq/lF4tajdPXAXPrdrihJrTU8MTm/76qUl8Ix/r5fL9tL7ONg1iN+cqKNNr
CAvu3g2+kH26lv/2+EGOeOkPGWRS0UhajpqYiA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50640)
`protect data_block
Fmz+ILi3ywuy2TrYL5y9sa/ekwyUgXe1i7PEL+DYFkgQC9xbdACkWIb6xNOn50701EFIGa2DsT7D
Tl4roF6tKyBijJN2UHGHsmyccFFt8LFrKyOlTWkf5eXTogcTzZ8GIvmQ86Aw/rwBsHDdRMcHwIe1
3oPvUIknbciCvSljfoYTtwRI2DvPfhadjdWBpyc0LfEK/MvC3QOpEaPbg9tLoRG69w2mw87eCZxs
jNj28bljr4fjz0iQzZisy03JNjZzqS1j4rILaahGP46EdLmF6+QxGYjd7pj+aEne9ZDqF/LYgmAq
742sbADVvpCV9MofY7bDU69ARM6nHcQRNGAfF0ne9SA0kfAx40XW8dUVqBZMK9MXRL8gLVfsza2u
pofa6cKHLk9nXa08iQscsELd8GtNcBCVGKmWJg45w9Z1LEIXMNoBgdAs6GIWLl8i+Lc3RbepbuBV
cYV6q+bXgey2nTW10cth2hQF456QFAbBOimmKb++W/GtgliOZ4WtTisiGj6e5CnunC3e5iGQM1cI
FLkRbA/1nU5jOKetjoaWSth12HLI4WH7yCS7PPA6z3NYiU6wjGriwelPWjdVLmmiA40GgRfRNlWa
amFFKKZig5lqmMlHtkViBKgE/ANr3HIFnaeSLWd0Doplx1x3WkXpGOW8Pn2YGu4NG4hBenrDgJLh
l0da40yVjjLA9Cd+obx6LceFcnqEWTdfqW9yaU1JoR/eEC5/EVjuW7ZXprb/GQJ9nI1qiYJy3Z8u
z7jLK+zBJcdHNE+iFUAfobwL+56GKAeGxLFrD24N/KW5QbdX/7pYF7mScFiXKLE1FxlfJrU08saC
GVQ4SqhllsAHhYaJ3bd06Ih5QDoR3lGkGwEwWXaIRZz4y4KSOEsq8/OwGNQp63UVpj+LofUEKBRC
VnQksqbWAfM9dQ/swBpeuInhzBgABjcQRM/cMf62CLSDUyP08KL5wtP4PIVI0CRGJ51FRCQ3SVXL
VhgG6wIYhgeuZ2ogH7+j4NewV3+OV6Z8683Z+NB2javCL+vtuiRuaYbzvrYkHjlzzgw2IiMs42cr
xIGBxJPWWb9qUJYp91moN9j5hm4Tg0wwNAVciY+uLunj5fvkQ0HjwZBLz0QFOuKz78reMCYpKkz9
FVdgkxdpq15HUJwIlwdScy0c7D9i0SnnmPEruKPEKWA/dzoWJyNNzW/11aKeoRIt8baxO2k5h50p
o36zO1HLyDDzY2RsRtH/u1AHxdGgh5XmMVd8iFoiXi+jSMy6LctnRvs2PplcGiHKXldoaQkaZxJW
naTwpKM1PcrkLEr2OhJmn/h5bBSMRWqtXbCiI5cJJi2G4f4fqMFswmefdJPZ5NVQIjs4CWcca5dy
pWW6C25PPPJSH3M3Uti/KIF+h7nFbLoW8JKlH7MibZkRSrqT3Ie4vxR1ZtECSHQTkuUQdrhsiSIW
9hC8bgDmTw3pDm7YN7MvcXx8vi1tInvQzBKGghNESFHXEAlOutGX+hLZ7l2O3nsV80ofMNQDJynJ
KdVTYHvvmQWxXleY5epOVYUwvOf+uIfsPn+2jGOmWosUcbYQFTKm7Kqv+BNwC5FlShfA456N17o8
SX5h8An7RGT60dn2sE2AV1dP5ptimjPMYAEE9pDjzzGq3jWFvdT3yXr1Ug5+jWSEkRH8v9Svxuvj
UbqbjXTwvtXoXdXRfk2SHzqFvqeDJDFKlgJcRA5kiMaqdAspCBY6Yde8II9NKUxxc2ksy/BCL6dI
qRKhkcVWUobXROs9qCRXnLCfic1MwvPq0YvRzZTTxRc1ySTElZR4wvTMk0Im1Dtl93JFjSCTMVKj
kAXJpbuqi7/hsqdfPAIArcHod6IYmjSjBVE4QD3ME59RKoSK7BcilxkxyRl3oeB8nJrYHik5tQaP
1CBjCmhJb/5dfDFaUw6MUeQhFGB4+608Af/hYiNbSBT8YdF91/HVoVAQPJUViYNaDzHR72ZX0By1
Kw3QpgrtmTfxtWzofvyZZ0vNFEpjuoSK0C5wcdg1hYF2zwYrvNAoOhEQezfKhnJKLAcboRJRZniw
MgvT42/wH8OTSPgEAe3KlzlDJOdOvQd3DDfr2ZX1Uo6UmYiIo5qU+c0amvy064tDMbxbiajguUQw
9kRhh9jlB0e7MWexh0gLBPdzM+sZQggdSwfeIRiY3zjW2USE8kDwcJA9PF/9H1e9VSn2o+LkVg45
UogVrqTiskCX+Pqw+prm09jlFwoyFJa8LECaDinHcynsTJhCOMW2JM4MM3iLt9ZkUNfp/zEBhMY9
LV8/c3m9ftERIoa5XwbsAk5Z+8bSFq4SDalaqY4l/Ftp8+9AYchKGxU5e5VwhAfQKWxGylj4lzSR
rbzQAyAwuJrEkivP90fDc4/jkSIgTlcxrjrCFt0mJnlIagOUZIiPqDN+koMONhn/E0bmKZ+t/4z9
adJBxB7EOUabiIckXx2MnDd0TDfvLi/27leu9Unr/tDQeEYZD63dukooiPUqzeYO2xzYi+TBoMFq
VtxHSs0eq+gx2TgW/B/uqEql9Jqkab0HXofy/v0E5qvUDono38FD48OIWOxpHMcQnxhI5C2+0U1+
d2TkL6cD1qZ53opzUXzFZQ6IexEV7bH716lM+fwzWMPj2DBW38UKWhep+jKDtuXNwKBVPxxgVOzc
iN0WnjI8yboVU6A2LnW7OmsexpFdnc5fDKYjX57R1+sIprrxyEgAcdmaNGVUWVw3kpolBjxUc/2O
5fO1gulRBJHSXBBOvmoBCjPk9jiCAaXKYn7T9ndzShBfDnXMdbFCds1tmCpMynaYDpmhoMR9iRoU
jOyLWSMOsDiJErPLSbVAeQadCsVjhDedL4bj3WZzUh2cqUPbuzIy80LxeYyCD2k+zL91n6ffpvFi
5WbuBwltBv76G/hZHlYBYgz22CnW57hHPArgX7Adk3bxxQYk2TC/qmJ1j7Um5bnKkBF15kQ5o24t
9zGqV7tJEZUIasFb6uNBdevNhViW5ETfKJhqPWT/+/jM9U6vSRmVVMVxegN7FMciv1ke/84+DiZd
Enmxt/lfl+EhS7/UDAiEvswhs1YweheLPkeJArRt/N66fVHUhAz63Zc/axcmp+GNiXzDh0yWrfIu
+gMIK/zIcj2upqcO4UZFK0pAyxAKr24kECesN5LjKwO5E7pPIdoAVpSRaeXwYZqWeON81TAVvO+a
EikypXzMzJxGIzo6vQZjchKHtG7cAwkyJtcwofAPLDY+G8ARIPI/dN0zNiyrZH6bzOFS31NQyjTw
MR0TcCrrfo/pz1vQwYV1xg+8bYURhohAsYa6yQqDMuI5WbFsLTFrJMxT93hJgNsS+1YGm8saujVE
mn/H3GOo952mKeU+Z3mgzaFzqcQG/MvpY5MjqQCtgb0D0XV4gZ986xGdBYgmAs+Sbebga0858666
vDdoE1GvMsSIIQjf49Ohd1A52qNKn5raVF2CyedpVBMVpMCxWEAqFlbXoESOiugiCH511wZzdgoF
DG/B6NgUVv9GnJ6FKVRZiVpFkO9FQz+aJjENayD0XXAP9+EG+OkIq2645EYKORYOrD1Sg4QsjssO
6wNfHIHbM9uSlqnPCnZI5t4R6EeoXptA5pNFBa4VGSvPeIMr11ElRBWd1hYeHublCMGEqSu89dx5
YjUwWWsSNx1s/yvCgZhCSR308FQHb7Zu1UaxXvDYIt8UB/ZBBq2m3jdS5sKzGNoQt2810PDgZJt2
8/s1eiYoyULzzMLifGzgTVtosEkB6+h6ufVUX31F3+UH1nbx+/ZREVOAkxXZW+dbxO5TV1eaXFXj
iUh6BZ2PVQRdAtifP4ShEnzIh00BUkkcKN3/H80XyO0Pa56+YoxXVlv9fPhJ0/u8Dx0LXhPHbiq2
n/iHuEJYMjCY8NnqLwUgy72Wkg39fqwIwD3G7tW0KOmWQhdusyzDPQvbhRTxO3TrDtRV529r9uOs
XhmcscYqYWDEY6zl2Wqf/0UWVTqLN+vvOq8KlyKlPI20YU0x2zlamh9e+HXl18zNehoX8uc/xzMt
wlk6INvc77cylkI1fHnetsForXKMOdeH16ObXYflnngZ2YWFhLqsetvfIk7RlCveHPUFdGE7TyOk
lhNy2BHvV6qlI4Lgmf3HNVlXpyPazPlwAtv/Lpt7gVcxI5QR+yl2HhcU0BoRsusXGNV5XuLItrAW
aqDIHEmOpnmfZ/tfzul12F0DqJS9GBpuDFe5CFwaLqjfAP7pcfDh9LQEtpMc+jdw+cZXJOMJqIlk
dCN6BbXz8SKOzVkdwQMRAXziN8gyWZx+cRn3rIkH7efUXwTbJlG3uj8n1m5Efwd+S0tY0L5SwbkO
yuACWfc/2LoP8BC9f4VoUqhEQPTQLtshvUtAbdTBuTGlcs2pH2WlU1odM8tJEsQxi5PePnjJNqlA
hn7+/2Xu+vUDARwAYknxHzIbvbqhgpmeMDzlIhIxvALtdjCGjH634ir3+lgqyk/KWZH3GoDFClvV
tuGRkivt5N9x7zXbAWcQXkHa0dhlzsHbb4i+DFKXwBvxb2apvFY/SxNNXOD9Nai0zBostpcEbdNe
kfN1q6p2XcW0lzC6tAq06Zn1mZ78nPVpp/bs33nCCGLs99qLKhh2ED4o69og3eGih/XCINY5C+9F
ee1iFmGWB6tKXnCTmvS8KxM7o+I0rQgNHLL9VfSPtLVn0wtQol0Gk10pNZp9OQ6m+LmfLZRjnlz/
GdfnF2W0i4m1+tzgCQeyp3cdvSFgFbpE3wltX9XpAZFu6gCj1mZl1aquF9O213ElPSSnIqy90P9y
xoobwbJMoJ56egupksJPpAl2ia0ZnoMpqS8GNjQWdbcJ3yEZ/N8kBj13+MCcqcdAzNvKOIIsHX6r
BoPuIGdiiZcVOLpQfY0+qFzQ7LQZn0yndpRmIJ8gyMeqbUBIiwjaXRT9Yl/6R1+y8MxOyjTxtLse
3XTf9dzAmSKYEtGuuw3/Epmj+wYRyN6VsCfMENFRIPrhmTct3zlAEaqGRxFQ8xJjD/lL/J1dfyst
j3lUZo5fGX0jbs+jRpuHOaAtzjzehlzSmQ30uoQi8lrqWNFYwvHtLY0u7GfSsyFtDO3yQL1Exvz7
92Pp+dSOUspA0G8ov9Dh1lO7eJ26dF3bMWBvPGXzAbm85u14kTBv59moNsbV0tSjniBpK3DOebn4
yl5S2B8hd2D5/bCegaYch0iB6/fxA6jls7drpp+Cv0LZPFSLF2S6V2BUJRx7g52Vp1W2NA//1fDS
e3X6YxC3PbcZwtpclv46CSUlWDPkmX6d+YiwqPNFykvuDNTazvm33x0MDzDXu/YnrIAs4tW5NiL3
2Jwi6ZfK1TVQnZaZG8LSjAaNIm8M621p0Kvi/KoNsCwFKNLzDXzMOsEz78+LFCSGNhjRoMTiinQC
tVSH2XRUBwtCUUxV+H3O4mR72YS+wSd3HUEAZo8Sa/fXZtLaLypisXTq7HV52o+Uz6QNc6MLDRUt
tOEq4O8FzAYUar1Yxv7CwCh8PXpf8xQdUFzdWReFOqJUX/Mf3nRZqlCCUDUeAeYP+pbJEk4HJOVw
/2ezdu4rkcVyBx6mxZMt4LC70FPjqIycX8lXdgaZHpgW/PKKUqXCoXa7NAHeO28eKUxaA1mwX1pT
CqKqlLmyjWnw44H7+3Dt6nm9WSnJWzvuVZJLrPB5G+pGADbhtOEay1JbvkUaH2ezBdn4ily38Jng
Trm8SPGxMun3K3ahwQUvPJRuDV3PALhsahWivk21ZB9VdBpeKpw1xErEmxOvvoErIEr82Mf7h+My
dNlqy2ZkbnnpwLmil3FZWSmsDm/REmQgSba8T+yLdfrTECjGxqsD432bLXB90FewIIkqf6LyQD92
3OwevCbNI/9j7zpGXyinH7baQOHUQrTs2pyaKRr2VSQQhqikO07KgbAuCxl+DWOdT8Su09zdKw+k
1xQc7pejzU7eZigGDjyzvdJ6H0DtYX6h5ntoc6AMPKnfTUjPCaBczOoPYW1K0ZBoLTdwG+eM8tUD
EzfqqFuvpSOa8kchqu4a3MXx9nWUU4U+HZUt6EJKkK03Sd/Lr4DuJyzX9/IJeh91KZChZgYmWAzw
J1udQM1PHIl4Iv06g/2pHsJlC76HhKgAFWubnrYJTMXrjCA/3L+D8P9Hk5Y5gLfzaic7frgnuGiS
BuceCscMpJ3drjrYSTAvj3pbenrJ29jMDtymOVnz4lV8xdF9TbVhueeyz6C0Jwx5khNVjJ/UjKD5
O9NLN8aaEL2QLrkBrfH5tQUpl2GrbIFR/bgBFT6ioECmhXbZKVWXG8jiCfgUEf19vvuugWIX3+wn
oXlNzh/+LMpUDQ7HWls6ApZKEgDJRpgwhoIaERliVfZAM0ga5W1ezPKlBODAngTSxDWcKkZJhpEj
Gi5WTG43A1xt+YcDqt2JePt77w3U0a/bINoL26K7mqTbf3IHQ901F8QsoquWzd1zeXpJ7TBX4MI9
3s1m4l89YGig9qjs8t7q7PtO2qaPkCPJBt/MO+TVmGdBYX6q+L76O+FM2rcR3NpqbeGj3UYECMIL
/tgACwXocPklEcksHOhory3dQTD8MpOxWIlKNtWHXPAC+GPGAQRVaYpRNTHDDIbalp88s8zdJYC3
94Ri/7Odap6yixAGGS9aYdVQ/jciXX0AlKSfS8BfabSjrg0c52zdhlxOKhlJQOvdPRq/ePkoN0lw
ot6L4ASRMWdAXX+657AjLD8c9j8pPaeTEUmba4TwdaUn8zo2U8PPR9hTwW4K/bPt9BGBc4CV/0iV
E9zr2r6UbmXPvOZKVRh/uKcJ33AfvAZUDQSsYHIqZ7UCu7DHGI5GjTEUg1kZ2H5u4G9KHoF0Lr9y
pK7QoacSNAX9FgYoBzKeY/vaC/uqs4EaOXFvqoJZK2l4toNEAjijuGFiaLEa3PtJ+QJysK8PgQU9
GwknsTDi8ZHsK6S0AaMfWW+dudoTi69fRg0+ftvK7TBBv/AOfHYA/B2Vc9mid7KIrJ7jvnkeH5Bt
GV0xvMijhwfwYrbB+9FXO+KUxjrVGdCaOAPbQgD6uo5vNnhJAYPGnTU8zVq+RDkCdoKn2t8xv/NN
WhQQ21SbNJOP4GzbUlraO06Cdq1Vfw2/8T6Q1CCBrWHqQQsFOzIjmkgSsuQvYnrfmETerzuwqSp9
7IAojKYCFilRVCrQZjbKjQVXZTfjspsKKqtzkjJeQ/X2nOl0w7LK/fhZ9wXWYhfiahKBJD3akgO9
WikIMWKdGtQi3CJ5SqL+66k8OPx40dgj4hsm4yVe1j1WdX1hWNe1uUTLN59QRqvG19zmi7zoI8So
Y7Oa4JoJCiAo0NmodaD6fsqKdJ99qVdQD/vxQMgTpiNn4CCpnh4YRGUNyI/0dmoL4Lmdou0wTjeb
HIAFl9TN3Afs02egl7X2I7xoEWmLrIOIt9QO0P6Fu9AhuFRxwfWQAfc1B4VBRjEsOCHbf66t4MGq
k1czZMGiWY05jkNOhg9d4j0yKf0178iRHOPLIrekuSuZ1V/OYc3OU4ybbS/CQu/AjhwHd4wfdStu
qNKMAVtybONeMfVdJI7ELeBB32RJrWYzJRAkd+r5Cijbq5TWnZlGAcXg0rgOa+ZbSvsKJBCAXNk1
KlkNc3kEmjhUABug0sJYZGgGQAsJePAMhDzhIGGijBKW+7F6TzqbQFYlN3+6ij4VBhsFiUs/x4K5
8B3daSxevZ+5utRTzlRTM9l+0qhSJY11dJJMHxC15s/pC/ZTetGrEJ3YO7B+fHnojbFtxA6hHVkW
HzA6ediRD/zMSrXBMpku6iEXH1j/G2bxLkkgKOIdEvw1Q+v+umiwIdVwKDuPXA8FeZkDDNLiVaVZ
zqEFD9Q6FUHA2uYBhqRRSJwD96aHPS3Y/UTl7t1IJukqX/e9RYaTe9a8yLCMjE0tj4hIDE8/eGIo
egk9l0AbhqIXdIitrYNMoeHL2Yl9nrMhmUVhiRcjy2tqNAJiNeLQrf8Tyym0sIX9E3HQhyuO0AGM
Ycb1Fu+hSe+nF6+4+cVohsu4iTWpax12lLk6Bh5rInvSYZ2Zo2p2LPSGeMIRGnnSby8OZmMz4/io
wu25NdHeB8NAmTEmNQ0XKQv47bo3pH3R9vKZkuqad54l7lGmgUVYxW0NAwsMmL0hm117ji8GKonY
OUGxvuqYNYsYb2hp3WIkL4oYrN2IHZQvRThBCcwk+0+Ev97YW0CiVx0I3G9L8UmVKOAgWU2rNRZ9
A21LRlAfaZiMtErkiju40x9tFejKyzvOP3ssmBSTUaIybNHmFSmVJvLCGiYAeKJ9Mc+2UhDXSmz8
8wStDotPsP1e4VS0KcFNkOdySKdA+wo+tzd3JFPlYszlfYpVNRPe8/gTeBoYmkpbtJ5Hh74JcWMt
6Yb4xkVtcXyE3i8JNOiSgb84OCVHA4SnTjGREt5L/HzJuuNWYoxZa3VZx5NLymyjT9R4xvs/4Pzf
16neD8Ah6mrNQ+0/eiVN9imU5Gb49Yb9Q/qRjhwqtXGdpv7Ak33DUMlvr4LtE9ve1WTzYS9Xkv1d
dTyG7/Ue6gdq51+GrssSckkxaE0wWUjy74T1oeUclmrOuFnfcOFPzFClcFl66sKaaUN0YBMZ6A4p
O0lpOvFsDGBp+zj4WUlUXXhlS6hS8I+HzAhh9ZqojwtJ4TJBslMqwvI9V0W9nUpj565J6dP/84Gh
2n6HOo9Hiy/dJs/oLEkq45DD9njoZEh5/E04SQbDPEoj9MIoAcfrIZdDAaKvPHdrLu00MOrDmHzW
OY5Gf7/Ptw1gaIOcguLxMes+zjR/874EPuGYkkMd1GGbbl1QCTToHT3smjkVWRoJzdv8je1ZgzXE
gaO6bbsNqni1zolarQJchZ/A7mlzNrzNfxuuYWC8ShTvSEdhg5yw4Iy3VPtH3G/Nj6jS/33aaSEf
nVNVJuXu7F43zbtwat6sZ31TJlL7xhJrRkXlZVquXzeyn4nUWJT1Oa5iKlbwonv6eMfO+u2ZCWLY
bp7jxyrHF1MHwwjnG8Py9Cokm2IAnwCmcoSlL2ZRsI8GP1XeF3F2qHXDUOsTxyQb2VmnkXhbXquG
bnFQAov99EKoGxqVGGAtOVDxCd7CztIp6PvQwedJYrwn0Wo8HnPXp+Dqq6eDe6CNVLxX5SVJfppb
5jj60vG95qWEy/REPI+qutNgAB7vIPjiDQPFWivoJf6lgmaXIx8hiSrfBOqxTA4eQM+mHjFRsseE
R922ONn1ntfzJRLGKLWiUYjrOlmpZZXa9CYZwQemp+3JjwW4MI5z3iH7uwvc301Ai0eb7gshCmlT
PUQ9Em4e3huH/AAvBFGcrgUdevTVZm1QFeVpacCI020EUtyDKSVwkAeaqMuyNWMMiMqFF7zQkrTr
qS0Yq8AoP5vJmdYVRWmvuD6drjS6ITJNQCriSsHKbFeThVQgkpubq+jAheJRFC259Q+rbgGpNQvn
x4V8PSTmbUEdL725U/B2x67fJWqg+L4pBgkDK9gUVa5U0x2dePngdjHgvMZqs6KeycSfbxtsrSC5
qwFlWgTEKgnZdXJJpWUMMhzIQkBnavkg1+M3BbtW3Kh0zoZ7JNW66aTgK1lKGN58VOcaUOk8Tfdj
Fay6sjNw6SgGf9fICbt7PXBquvrwbqAz5hdwiuyUv4dnWyanp1pVYRHJ6hhHkPrd5KZsYX9gXddh
eN/9d665f59L2n/6H/TN4tCyqUJclzVMQZpzzinLwkfa7cDU5vKtS9dK6uMvLlr70D+LEJzl5SM8
gdhFExuTkB2COGSnkA7zzWugVgyHokddmcOlogWMKGCM26nTiwITjIlpVymtVoOvtW8hYRVLHf3U
wBzy/grOS1zJTvwqxJKqe89Hkl5Ay1CRDQixoPVJStk6V0Otsd6h6ZDiU5cbQ40Cu4PdR7sq3Zuh
4PO5xk6htOUiEyMf4WjTwOZ3oPb6ovpF5IziGk/r2SplgHkYLnkn2tWscQKTlm69fbR3WqmuGVO0
qJCHZJKUiWmPwNhQzCTHO9C84Cdhj2eyuTtLWJFT0NFGa5mc167/QqNpRV7pftbigXdbrYPwtsPL
1nCVAF4blI5WM+LKblItuiOWh6pr/jK6yIzjt4MWjLXTgVy1Kn0vKAFUD49HnDUNS21bogloDHcP
YcnmbmGWkaWbQOHoMziqj+47rEfIbt50WHOJM7Af66jcA+aAUsDCX68hokdRenA5PvgjU0CJu+hU
LBCEqSbzTRklBoN6yscJ8YRo/PNz+MWA3X9ql7iC3xKw74RaQoct+uUbW7NLC16w/EhafICOeNF2
IDhMmTh8KxcgDQmxz7BwKgq645XUFz++f3H4IzwEmHDoAHC+M3vTDijiZ/bZprhZWeIMK0ngLpDD
WVfy/7m0KxWcWSgm64zCt3ILw3eIT5+BXAN8x4RlJCheypc/vuOy+TARz7y/o4Zw4XzdyuesfoIX
M33olA1QEPIBAlEog61HGJpx4ZCHSI8Q1FJao7kG0zQYfOGnnXEZW0O7/9rYU4P3NoX2hUC4stz0
VqQRMh+XsLsH41IQGvRb0psjNCcWRzdQMgFGUa/zsbDlSn5TPSF5XHywwKAs4vPK+g7loi4eJS0p
efmouuBJwDNZubjw5Wi7YemmZBFGmMIaBJMdZnYb8HxNfxIB02kOM9RQe4XFPUZo7SSuDyTN6sQ5
GCAG+grZdQFsIAtSEtLzmdkZKJ/LvZDiWQlfmt8QA9U6Ygmzk9yKxGUs9MLltYOWvcNdnA96zh79
3rDvHi2x3mdrmPQ/KVCat63s3X0RbJe4sBk268ob03IE526dKic1S4YuWiSmx7gtGs4RqlBcNrda
5rU3hf5cMKyfchEtbbDVGcMfJqFqTwYt0fTzZWucVK9Ifbr9mufwMiXOZDk2P7y9FiI73fL/g1Uc
gd+Yyt7cimEf1Po/jCLYZ1HHpNL2hkhaFSrplXvPK2SU/j0078t03ia0v/hXkN58IBum2evUFYiz
aOSNi/c8gsu0UaNtETlOvUH0c0zsQr7YAuMYYLkYboV9O4URH57TDAvcu63swqH3Ui33cWfElO8o
NKFQCG1Y8CUhTeu49cDr4unhET2m1aJOS5bPRAUdNdP0OXjk13kZRUJ9yiSNor2UXttifnklFzjx
/QFNNd6YTHRm2MSmEEKWsRIxCQtMp7Lw4dMx7hKGnq+tnYT0XbbdR27DF3fD4KApFlquXWRaUurd
tGzDl9HmIejEqqy36LO+nlPgJp9RhchSJGqE6+vArA7w4O3cGEiQf0Uwxizsn0saqD9l5U+lzLOa
WWDPbjLyHhhwb0nRUd4Xep4+QXaOLQcTG1Q4IDfYK2gwQAzR3Jg9aEhCerHIsXHb7uyNSKc7peY3
Vajvaa/Eu7lPGTKU5ys7Qmnas1Gphdam+R4FsN4YlEx5lowAArQpocI9j8wCcwUnwvTVHQK/xv29
nLlXd/EyFCdL/WC0BfNFeinEoisJNMqjYH9loF/CORzN4W7VG5k9W0o75Sn6X7dEwShyC270eEiB
iHtVRA4g14PdOkccKe+ENTDY/7rSt6t6SBIkKfxkO+3s0qStNnVaoQsWLpB583e86WdERSFcWaJ2
mAmUSZ5dzREiCoigytAuzVDECIA+vGbalpe6eZUXTEpnBjm9JFFrJEydWh5rAdcLHvRxci9Ui1Qm
9QXFMu57Zd2LkjFzYQG0lEmQE3serb4zDLeIh/2CbW5Z1PzOD5t8yOdEW62Wd4it7F9En72R7K63
NcMH6dbGWMYywb8Nq9hxPR/4MTcFDmTdsJ6hO4A8ACVxG5PHMPTvrfbjPDJ92zXCXjgcqOiVRFlB
oAaUAUvXzH42ygtFjLYCRJesJ+gYvq+cNxIzovWkhUABNyDjQ1h3H+ydQU1XQQ2NK0Fp0Wf7231d
Kg3MwDNftQFhQcp4ktQ9eS4Vx+9KjAtObd6ycOpeRU2+1JQk31QnRx4esJMOXWBRQRd1Vx/s+t37
h1AK+tr4XUIZifLqYWnDloO8kkbaCeXj/jWxJdxAZiOb4quVC4iQnh7CboLmEz+Kk3K+2sgdpO7X
sCiP4PlcxQy1pkYzismDXjpbAZRaggqfnONfBWOUiCkwXRxfPbEl72/b7Gw5ukG35Gbc4Zcxvx78
RYPWXNEOpknSTx2O0kLymnuDqqPreQYS33hYT/Z8iJfFDyd3zFOOAv96jWFOFh7Ou7jeX3OiAMaa
wlCZBOMUDtoIVGS0XNJsAN7wAaxERNfN0Cbi2pE/uO4dGNPIDLhKclAzlKPsAAGqFhw576qlTt0L
CYbEcsMuF7RM8mF9mODKtHA/2hAVeSEZp1ldRvWealWiwsXRxy+wk2YvE/JNK6P5orU8obOA5w+k
ZaRV4+e1sEr1hFGbzrFmYTx4E418gEP4Loq0rb68uxYx/I5xe18H5TBmyYBZYlQC8nLFc78qVyYU
vTvr7CUpYwMHWdoVqd43NqX+ghGSnqnvZ3nA8XSSc3ldKSDHvc5dMbVF9U4lQYGSv2aevhMMlLo+
7/ZcU6Am8xYVsDaWJPOdrVYG73N3YrQHNRulFvfjNN1LEG9uQ7dB8hhPjkLEKbqZfLH4zAePdW1O
GBcocbhiKv29fOgSMRC6cttvG/Lt75VjJTjSDU2qJb+PK1d39Zh2bVzv/nKUSjl503n43vavy1Pv
qpN4q0D5ipjnvMPguvl1etZhCtMSQumXGdsR8vbdc2Y/ZqcRpqswc4THBWRHGPklSXID44TfYV8w
/VSdggUVdFHX+5r42SUQRzITt+x77spW62RznUdJ0IM7PlctJSWAhEExj9ojtl84hsXbQA3sbgmF
wayy4dTFu6NwfV2Xdlmkxfk6hj1oAXSbliYfN8ds0KIIV/mlhGoLxtGYBNSMXNnEMoyu5Me20q5x
a3D6OrrJU38E4qT8Nl1m70g6Cqv+ts/y6kh61Lr87a1J5eueJHYPZq3K5sV3KTVWQBR4m5hW6oHL
txe08fYZM22qathiuaY1cyKz9qZa159NuGtc15sguj77qaa4KbNK2wGWDX71l9Jdc229GRLiKiAw
tRdzraeVIosBwiheYdxbhZ7SZf9DoC54tzMlcRSnmS5zUp6/Q2YvunYcefQnRyVadq+RBPPiJWQe
uIkRSP0SNnW6Kp1ByusniPEpnppndVfLYMCE2PGdh+ffIuOy8FOVPXx2X6lykTV5mQvKR8wWoE1c
nMi1b7w13t0H7YZV2cYjDxTFm9DYtAG7xCNp1wGQwtxN0MTSxh+yg84JvXABnpo3exMMpIlGqPUB
X910HcK97j4KMV18UDRDr+XibYZzTKzkyYbvTqzx2A2QTLGkgbs9ro+NPLbidi2K6JyD9WeJoCu4
b1rbURm5lcSrYF0oPpHFBo2u3VFCyFQjH/ENRxuulmMJhs0zu4zPhqBoOGGa1GQAFjLhLxk571rZ
IZvXugVmoDrYxPGqlW5et8neyMWpnI4GNqMb6xOw7cpoIO0X6K/cVDCnFvjG8u3x1+COLxbWJyAe
eRTZD2ntVtfJOamjILVnLRv4bviGISPFq/4N0gKzde0+gpd9apEe7UfrB0/Pm9UhhyP8AskrZRyK
5WFR4M+KaIWL5M8BM+safBGJSwAYRXBgoc5R0Rp4bU66Ka4f3OdFWYfwKLVqLZ85uU3cCNs1LYdd
bMe2swJjrBJDUlEgH6IEkYxu/k3Kgi1SRLN3aXbwof45jPNGjewLNJX5RJPuhMFQGfr0j6tvkhvw
2WxPfMVTqfiiszqezRygh9pTQ/zPfLYdZ6ZHhcR5dQ2ZAdPxSyK7Eq9pFOQpL31SWeDUUUw3yslH
jMwBZw5qRlgLn8hkDUvEBK+HJh70IalFnJUbP0IWsezyBprgbbiP5+ojpxMog816sRoa23EsTxSI
JWl6BX7EMdpmmOku1D8bEH65tChsmeJXuzdOZFxotSd+JXALesKadcHqPwHyD8rKVay8Xjlf+Aw/
073M9Axz8p9Z0U0nj8h0RAJGjBjBz2rckm6crZ8Tf9neGbYk2T2bkuBPOg6CGhmXZaybAPIUYQeh
zyK7H5ZgQAhPaeiV91152XfgIT5uaVJxVkEsYlCHEhHK/gEAiKNOkO0J3VDYbDHgA4kjdP5sJL5d
Y3xUwJ6uGt2iKN3YZHjmbmXKXx6N5GkqpdrV9wLiMvOS9D9Sj/D/as/bJ69LyrbcGWeejsKhWaRk
2T7Enxy1n5olLop2/LnVfYw+M8RyHOVfpdBqc7uwac6U4Zc8GkoYL2E1oRzOPqE9CtAL6XGx6bIh
w8qUIxX1CXeBwN/UpcVEyHNunidJa8GVpOsWtX5PPpv2M5h7YKhrDD3EdTc4nf+driXE8TFz0zYT
hSmHGL0FeyfQvlSBWNzFlykErP2CUFJRZs6QI/NIPYDDzsEEPLM1+pUXl3XSNednF5JrZhDfrs+M
qOrnjC3l+S+y+STU2w9mqeRAO/vldZviBgN3xekkmhyl3OqvYyqjYXMSPxxfv/Z47e62+YLd7igq
GWJRS1+q6TzmwveDJD0knfh6ilDKXg2KntqComt9hJVR0yjGCMQ+YJDZVh9HwDiZH5GAuPBUCvzS
WcFdQGj2S9XTSnWQ/NDVj2gQTIaqhSY76g4ziuCFtD4p7mEbCHuj+SC5CmQnnOwjjvmR2AORO96A
0v4DS+dre5mOUQk2dlEiJnodwmfEPoQHYNsMghuGzt3PHrjkx3Qajid+Tt+8NF4a+/iuZD/qwFk0
GUnK4pCdG20XTP+HvqRz3QcZi67LWIsUP/04aKrQIYW0f7EV5FYBWCcVGMPHmmMuHE9vYlJZz1WE
wllABzM3THa8nQZb/gZfbrjAS1vwn62Ri5QWdbuRagrZrQtLSDJ5rnveLm/jib3w11X1y3ctKUxi
MJl9Jub+UKow+/CyW/l8u2gpZqObQ0Bv4b6am8WROtwYgi5DzAiNbOgqwasPmYknj+iuTynrtAAv
kBYLDkqJXLxOPU09vFqElE8egkCwDYqE+agfWWac+liiQCI0Fh4VWFkW/ExS0DjguVdBSR5rRQCE
MhP+2bNU2bGikTZ2FzGFLVyrhDtX18VCew9ApqfXd2rgN2YCYipvCBKtQI/K7MgsPjoeLNVWs8ks
rN5PImHkGLCZ6Eg6u7lHbWHdaCBwwRe0gyZQVLIvkXAg6BlBwwSWkWTQFlCULAoEqB7vjL6SHNrv
j4MSHRukocwt0ykH5WW8HKjwxOjsIC+JaRiv243wBrVWXUnNm6iMcGQSdHYW0VId7/6y1xmjdnHU
MoyiaXK1fsFbS3/42jzJ81Pt3z5v2icKfQi8TExdVWQzAADzIwdXaY8E7cCesZf/lQ4OBj7MBiJD
zokVkEqKAaVMGMCmzHDIR6qaA7mEsrynQi4rl20axhBYDJLex7CwuEOslIhB3RuNdxH/d3mOkSNU
y9wE470RDA+SiworR3ZI4csnQLaFHr88fpu0b1kZxQ7HDrDd43feTJOUXG3JW6wRy1h2teJf8AvX
wbeA7nqYu37OR6CRC6pLyz+p3jwUoGYuG0ZiC7AIgcsn1/rlrm3uO4l7XaqeFUjUivNs/0NeffEG
juLPB4pFChX5GNr3NHOiiWX4zrdxKw4apy2IOknxoMGNHFM/AT0ctZrRxI2FDMvvmrjZfzhUhqbV
NpvZ58OneNwsH9yHwjBazL/Rjsk09dq2N80Z544WH9oUJuTWXp2WUTzFEJeewLrfhJmqne/hz6Bq
nFfqQgvU8aF7MeUJ12zy+hD+GZ7IqlXplIKrairxEJE/8vzvsGTAUhznteVSanu4QuEDH4+tevIM
vavk/d2OUsdfQgk+fXyNlAKODp/l067RiDVvueiXACeAyYu+ukPHg/q+1dhV2wTeYZDVwZDTG2xZ
TUemKXYfeS+ZlDupHFNz9P386vvPAYPMKkhQzLKY22uzkDnyfIRc4rwSYCHDjwEh7/POxrKou9m3
05dMEroQu6YGS+RocMkxY2zQV/zvDtoZrlcO8h+TXrg8/cvgELBhwOyADOpz1EV7VQReruxL1kXn
MWIN2jElvwl1i1+5Jnt1zkNtDvpuSA+MPSzG9SLUhoilqYo2vGpMBTdtWxxEkwMpuRLiOLN4kux3
FfvjleM7BPJJNM6qQ+TYxDa83XA0c+/lppLGDC+t+9vWbRrNeJSuOa2wFpxluEcxruXtGJ4faUg9
YTBwUyhsYXRcp8C6+70dbtTtRDFAv2lB72+91cy4zksKmb39o3yZdzASBEwXdqFWOyV8Rf9ZFwn2
5Ly4omGiAh0YMCcNpNh5+5M5k8E1k8dsMNpidHXLsJySXLZ/yVU8PW9ZAy4FUGQmdyjEa6D65L2F
TgjbygxpAw2/vOBMcjoyv2UdYh86Lh0FssLRpdguq+OG0j3CfteHXgDxn5ObS7yVz2swV3/32A7z
GdzmcYVG4ZUOOTs8OrwB1Rpe1bQ1Me0v+8iBIzWHOndd1zWNxGu+s3/nGjfjuaOu2m9KCReSTocO
2CJGytSFgoA1hHoB4TPtnxuSX82bNIMRAaTSWSGRfgCAHdI+EoyAC1m0/NB2iMR/kAOlW2cJNCyw
3SiJVXhPwE14ct13Q5BkR/iPxSqbgG6vm7wwKsO39vBqu18rfqp5kmncnO8kU4ZpdkV+mmofiKZq
KJ0G+XlcnBfm41tWkgm9x1XdXdSs3BVpSYWlWPhTuraRcn6F+j7A7eIc5hytGaExnaWt/hJ+MO8y
34aOmxcG9ByZGNkse+zc3QqmxrzYWsuKQKYgOkljoYQQF9eYBq8HDZ5tLY7+Z9IPID2d7H4BQ9fy
rmeKSwSXH7oy0kxkj2nyZRbuYVyNSPQHEUNqU797JKeymRAxK6aVj92TKCBX9/EnbYv9NKdxWDkt
n+VFG2B+K0ECMZSqaK/ihwL78T2mbWoTybTyZa2KhOoV0aakQ95mK+SE7X5tnRvfgNku2SYtwUrl
6kkqbrI44EkmX8oQdT/F3/To9juk2deOR0ASNjAmPxQgKxdspBjoF9sMkV/cTXk8lfGF4KEs3BbL
8OpsTywR9+sbXKJxNR9afZYP0XY1COr9clBZs4+qzekPmUjSskf3oGdkjKuKbe5lcIsGWLZFdxz1
odIorYQTJaOsuDH34IHPLZUEH8Eui5mSJ7aNm2R7hank7O1DT1uiSax/bNMvUDvTUmcy0jmLnMm5
UdOtL/Z1mORj4uo8VV634ZBr5RzidDzm2n7aEXdmsfZARrEGcBsbrTWU1wWZ0qXE+2vrH4DCH9qI
D2byMenXPlGpEVb/kAXDzD6SBCIMHjtGdM0tRfOycvQDtQgqrhtz/cUzGG/K8p7BoSkDKYdp4kDU
EjeB7gNvfx+uWg0Gn0aKDzHD4jwgCEBpaFqgXxtgvkld1tmHNF1qaGskX3TXcK27B9HcJq4bMSNP
QAu6oC3OkI+RFVGC4Tm/vStD9QPLlLnsBPlzZKybX2i9XuJ9nPCLkVeYGrJ/hOSdAkUIJOddoNP3
eVj9kuo6JTdIWN825FOzv5uBWZ4hCjuINOCrvyQ8NKQ65gNntVLVfyl7ec8Ki+HCBxdh/AQF8fI/
kGiWfnflVZjo5HllpyIKMx70Dev6S6qTNaszGDv6MJmCY089MrB3LnOgALH0owsav0eMYT5fQLwi
bYUyx2fhzeKtKTKO7VfNLrabKypVINqIpYk6PlLa+bONOWefVpPWzM2mNNCzpJgD8QrlfOog1YKq
wnKC7R5omWlZbaJX6o6lX+JM7FZCuhJidTqWpG18dUTTekXQWw1OpwlQw/bFESLwrtdnFVtD4hbD
gqCEc52dtpefXbd6ONVCHuzVeVued0S3wlKky/Djk1Bx2Gecdg/qnOS3uXo3z5gzDsoFf/d3kYYB
4eXIl2Wnpa6Wg+PArOzv4CBGp4ZVubVhCL7J5c3hFCVGMpB+00AiEWjAJJEjzRCPR6Qtb4+PCIKu
zcjo+DbbprXkjYCOqtkk2PfyLIi2tuUDdsWTllZ/xqYzGlUW2rd8IyV0pTm+kywJJqw+vXz8GUK7
0MLbVISw99yvYm8L1O8hbi2hcKVdnGi+woNSLpd0KHyWinrWNoQx1Z8aRgfhEXA9ES36+SDuQPBl
BL+3+UHVJutjfHFPsEFQd/Cp5YnGfjQuh9SXHQPEAollIK40hC2hP9xGfQu5kxNveGEyyQGD0lan
dtU2qGwz4m8QHQ0bNYJ4t+inLLpGW2m++rcfQ20JBxT4H2+vo2PZaAWznjeircTwlZZ5sXzNBXYU
IJQyAkvUKvyjKDoqZ/qyIwNTRVXz9EAXdpAhk31RRrHnzkiWpi8m6RHdYYzebdHW7NakzjsNHSDb
lTisoQZ2iMp/N8v3KuS9m3p9rW7jcAk7GnMG+MXZoOBapXdsqf4nLkQ613/Tw8rSVDIYe5IK9gVl
jiUysSY1PReWhwiusG6gtHfsXQN/UT84NwAfAKe5KMKHyPy9u7RboonpPMQ1lLwzbAzSRT8SVcRr
/X+2qJsgqBCJuWwef5qNCpHVK1TmS2Z9scCBAg9L9taygNs8lbVIyl2QzkSlfkRsZOOY2ob37Wid
qNjeaumwiomeoTtZwlJjkq36rLS0xeSiCDvaO5N5JQ7sN0qoTlGV4gUoH+DiYC6B58stn3Z0tN7f
hzLcMKE8eSmBKVTY1+f4D4p88hAfpPwTvM04/tie6TKNHmEcrm1tJwnlt58BogsGZsVEXC2Oo6om
Yv9ER1EPx2BQkSDp5ILQyy+v8ZlB610k0sAmK/3bToylPJnrOOAvCzHMfcHve3dcLx3+OjEsvlZq
P35d14/s7UxdW3ePWE8YvrYq3KwDMHXX6IXyYZfJQs/xVSQivbO5hE/t5quyW2iN95injdlmKcyO
PV8KaLqbfo3zGrPO1UtpleitiOuXWbHl+1I8wrNzRnU92N56i6JyBPZbIc10hCToKouO5/lE4nv5
/XAmogcz+SwQrYTsaQ4S+TLO1TGynWr+GZU11E+U7NwX0VaPoqYkXuq20iSSHxUUC8G+Y5EJDUUc
9gyKNs9ipy0q4CxGO/7IN9W+WH0sBLVgTgcPB+VDDtNJNDjjDA5ikFUYRbZj7Gx9fKCHJashY14g
nmrc8en2r2bEeG9AAX1HCfYQtY1jPjHLUiaflBSMvSfuUiFyGYZg68wL6Kz1xm+7zwc7OJf0KlmE
u+oZ/kNAIR2kOHn2DA6d5wh47GoChwJPdJHq5SeLcD2L+I4A3ezf9ktOCYXFSSG96GSC/Chs60xj
2+2ok8ggQjemMu0nKZZEcCtw45ShLgl5hmYBh0XeI/+F1EC7YxZqxqH6plLiopH7UtxEX/lPXTuN
6P/aqU1FBIVuRiVVYMMJOJRG4yhVVtSbCvOLQVjO2qk+tw2oyUz97tz8MpJvEdsSQJVndjnBKV15
7Juv9Sk9wb82ZA81Ya3EscAZFIWezQt4rKHXLfB+BNDbUNZNAf/pBQvXZg4QbtocMl+ZdkxB3KJ3
LB135MS6Z21eZCAEqtYl5+MRbKp2dmWQlks7DVIC4+M5UMV+c37gOnWfL+qJmQKRKUod172b8GEw
FPanuzi5RfiP3ypj5Ds7O6zEy/jeIZlVy3sE8KLMMNIpkr9/A7QZjBRLNztx1ueV3sQkWjfyofOi
WgtF7I2zwWzGaws4c5fJD/MkubujQZB/ymdXGH1RSJ4L0dnZuuoZLzWdDzD6dLhhbViuiikMcaHS
qCP9FfKN0bCltxvjPpnXdDt+utFWp0wsd2FyimSMsRPZpldeM0DW912FOmXsEAv+jDGnkonBE9w8
Jwfn5hUMSEkEoj/i2z0Mssgu7/KGy2vFjUp8u++PIYrIxtq4KxGgk0X3qH+hJYAG6gcLsey7iuRI
dwA/VNd7ex1uxzAHKktdviCvZxantga7rEG9eM7p3x8XZaiz8lV1askBsGSObNiEac/CLDG7dtGM
fDKbW/XMmgMSrSLOdyxT+1P3+LMFq7+EihmtKwTLxaek7mXSGXueAWc2FpAED3gPL2NKqQLSp6Tx
FCKGsGU+KCUuXZuZmUFPOZYURbCuwX7ksG7zkQcsA2gUx2ZlJ01aOuCm5rCum3QWOXzGsE1hQsWg
8OLW+F97yVk1YqV03R6kpZDGfskHnnGsnTPVeWMlDKeOlxvPwNFjEGBQhlIiCYAjBovbSfXwOiGX
X20j29Cg9RaDfbNg+CX/QlNWTt+wBN1ro2DItzol/C9Xb7tM5QrsOaEziNzRC13jPlAkk4+5qcg2
w0GWQ5nl1OB20j4PkT+hmrROcRVukJndRhS43r27kr1YfkSmOukd0TG26N/TPrkSi1lu/4XuooHI
qnoCZkUd471zCEL99r2xZ5+/svDt1KkODnapH8i7cRYPEcYP4NYEPyeFOEJa65EGT8k2L+esEF/V
Ch1GXHXXVAN6+qIYCmuWLUbT/J1tUJ8dZLkn/9ihOuOctTyrYKrvs+gXGaheWBNl2GoM9kQH0YmQ
FjGvSMEje9nqNWpLXwOLY/lQPOHVabfqjXI7YUbGzBm/T4i8UyAedGYZRfAMBj8gLDtf2Qke4Z6S
7C/J3c5xCNz3NShU+1UhrzjH9KuDlfnq1c7NAKPrRlLpT2Me+scEQSlVt/JpkSCUA9snFhdRQvAJ
iKr5+hcuMVggF6bXSZIZw9HPozohdyLITbpZTWG1hGaQnWrsdLUCHlAYEC2OQzdhHHitoWOmZEFb
PNGrh/Bt4baJtawM9I4K8cMF2P6qP8V5b+snK1Xm9BJEdVMeS0oF06ScANqaJPpzyD2ClKFPlWOR
IhIfSdkp9Sm2hLMkbR5I9opyRN2y7Zin3mxNOaY2S0Ahn80XCiq6yNFDN93B/gtFgW1LfgPFSSox
/CRq5FsQvYlvimAoMbCt+wg4VpXYBLutHNOFuYVKv+OrC2JldyIDD29wFpyhHF2hfYLv/1h8WPgO
LzD0qkqIYrgL2t/DyyzOrBYIT76j8kz4RlgU47RSfO8iYUoTGg7VH0ZH/2lpmcGgchBBsUME673A
epWXj/E7nJV/x0pUwFVEwLvqwPURiJY7RfKUhAnEOKVrIU8900UjJPOTg5SrvRmIBonJcZmaQIqf
6m5j3G7FqqUEwCBrJ86TXSWWritL74FUI9+WuHNGXcSNjdkL+jhvLbVtl9OGDlf8vmIaIeiSbdpY
lFha/50X7miH0UdUoIcQBBPSqzmSQ43s2bwxaAlr4h4dvUBTnMrfO/sBQZQuaA16fr6hh7mUJedG
7fu0hpOHjbkmi+9YDtQV8zJOrZDHgHx7O31KoAjgOo8F56dnr+pSBbPtgFlhtmDo/QBUgJGw52GB
16zA0YAktbwAJwOJE/9l3NR7N6ByoZ4S24RL19Ubs7kCWqsml45FWYm9Yasg3tIBPswGWT2uhCLu
Cgyvvcr7GTzNsm+xJy27YV0cL8Y/YNATb1U3+iH1BLcnHhJZVeTuY8pJdMNQE9h30hN84xcXOj58
ZaiZQPTDidYtudvDRW39jr93HQll/LHMidJm6fQPOlbyoFrO8gTEaLk+mafMNwpFfM3QOmVKHl4z
Ao6U+51bOpv5wVEl+PnUh/z/JkrU+Uyr2iEmsTVEtYplvbyiJNyACHZAbBz0WtmS2M8sNEKKsB4e
AvVJVDBAcRQrGF/E/mwnT/5RIGBGNDZTJPe0JPJ+pYDLaJQOyPvJi7pm1DCDrSxhmiHTPIfsVNCU
0gLW0l5l7VQxcH0P9Lrl/DgG9+a8R+/mhMQUAXRcL8BRhWAmewhoG6nr0Re5TouyXTRlOG96s0z9
WzvfE48tJDL4u0gmomLSo4TMJrg57l71Msye1RIpwZ+wnypJdD1HVSVCyynUKGrkv1/thTo1zQGH
DSeX76bu9dJGkP6QxCE67KQlLRFyuiOh7/MTg7A0i51yP5ykhFYu3nGXH5aDNA7iXMXAN+WGFByA
C6ADyxsczrDNh5ztVwmP+nerLXS4Nw5iocDmTBTovXlf+L1YHx0KV5BzdDMSmutv7O/eCCTyiCPt
r8e3QTRstu7RZ0xA9zxPWFH33tSbR6ihepfkfOQYDF3Kp8VzCwzoqFecmaC2z4q06T6zuvAD/U+z
sIGpIG621ewQNaAumPn6yO+bt7SxGCV0V+2LmFy+DybuX+/kHw1H+xhRyswtpkbbfTuI9KO+fDGm
DWMuDX1IJshwuesI35o92SzWiXsL09FHozhcTP00zc3j+M2K5gz1kPVLEOTrPzxsCuzmI8EjPdyc
Zfr9YiRpn4qdqxIXLEVCptMLfcHWKILB7sMfHHP+y0Dq00Pt2nkp7qIq7L+zdlwlXcGzQWuvJrUE
BKh4pRH2hQ6Ntx1qtWZOngmcJ9+1voyBsyKxtyJ/mqoOZaD3ZZpAeRPXitvxw4MNHsSUBloaYET0
eWHmRg0KsLyxUb6zOiIPLlDyRe6YQwCYzZUm3Yq0RV03Gzu8XHxaH5MPvY2SKsE/Cx5NQYK3793m
sCDV7d6ADGpv/7jLcm84kVPxw+EsMo2hoz5vNJFvZHAajyS4roTTeGZUeu/QV8/vYjRcmuC+LUKS
utJYjRhtAeit9Qmrv0Pvdbd2tXqgtkMrRW+CkW4aO/P2fbagWofg0qFtOQgRbtGm57E1GcjcU1Kp
lLVT4KJ4thpuS9GAqSJufXVPPUTh1cGJqnbGC7AqwiBfkcPoWDvmNy3e6OEQsyjVkFhE1fqmiv/J
B2sOHxmxDlwAEBq0UQBE2Fd2EF1YRg8s0IjECjwngL48UUyDM2Q9BgGwVcFgAzjkIeli6SjNAOrp
3U8gRWGQ3kpOsPpszzWSXeTuro3EzI9J6hSm/Naeyzfxr4+L94YuTsrG/y3IeEKPZDKazfXE4vyc
99GNfykUovRiTPKeXwt+M5t99h/CTYnx8y9FGw/59O+1Llns9TnWHYgav/LX2ssmyg8kzIaUa5Jt
PQO9TEMF03lNJ04yjqy+d0w/CSfAM9MDmFdVSEDWeACfIxRIXNLScMMpsmawc2u6O9C5bW3cp8gQ
3x3KgfKQ+9pam23d8jy1f1lXu39HHV5Z26uA0LL/67HoK2lPag6sRKQkTpQrJphhUlc0umsbccs2
E9ywqJZ2wNYXxXuCcE6CRmlLOv6SoEk4n2rkN847tgmJhhvqGqrWYmVNxFyvk+v0flY9ueuQa0hS
/IN4otRTF90UWcM5ZiDMYhSoAD8UURhpUxO2nWygoeUvcJ5KpvOsh+fSUbbdaOTdgQ8PHLpVMxM1
U3dEnmmjiKE/qv7hSY+w2zjz3XPHDK5o6d6+mu70DJkU08dnBRlo+rqwBngv1G+7JtyMu6UGO6ta
mf2b9LjJONeIXLYk8P0XRt6GhN0Ja+rcT79/eeBUwOfPsnnGo2+3+M064Ru2I5Wd4r0MENuHFe8K
X1oBmC7eLHZ5TXN2RXVJRp2mD0DUx+sf+FF2CczWXz9C152OvpCNjK/6+vNUj1JH33Y07kJgZ0Qh
qsYA81AkEXw9OIyEudWtP6/N6XsOqhH4kypWg4BCP1G46hRs9YmS+URmbH9+tr5J+CJ1mCQoAsbl
MBIKWZXc+HvXOOGwfHPmXvdwFTHEaOanC4zONJTVn9ubWMGndmoFHPAFfuuuNqWIOSduDJBBqtSa
bnOnL5X93WVr9Hv8pPucIHOJCYrvFsTArss+5Uzu6NgBWgQ9499hhk0Yu1TXs7ANLhOHQbX7+Ysl
5NED2jp2rZcIPrQ3l+NhO8yJNggPLMugLgOvm3Xdx/yxb2kAb3U9jUIzM5F7bh323q4o9Wwx+3Zn
KFpZwLsYXlwpnP9OoUH7DzZ1znbl5MxnF2GXfFS5jQ2L6OX7Erve30sXiR3z+3VMXiZtGIBInEWl
NjhILVu9HtTa5MLHdcaEDSQ4D3O1OptdQZf4y3nqQW+wqwb7ySYJ579T/nFDGRZUAaUL4k/WMYPt
xB4HIHHAKprN40dPIKSHOh9YXrMzRXUVnicSMHXNeiSMbuaHnaRDOaxvR3ZCL9Lk/Lf7WSL85Vqf
l6lpf1BOuAALH8eKNRd85S91ILO/peq6KVpJwj/rTeGQHwsAI5EY9dff5NjpuXl89DxKLDwEUAs0
suxk6bRLT+fjFrbdABtkgC/FjU9o4dOpiMZ6Vpqoe7jabhQVd/XF//yHEAfzD4WsmCBphwrYwyZ+
+rCeguRic+yEhpKxfdBSZY4hIybkvpST+uzylrV70OhdN5G1iwYbhx8a4pL+ALX4eiKgsdtpJI/f
lQxbshtjPqA4EtuPMOQeIlalGBjU0IYcKFDtbz4iFWgAk25io36gE+aGtCAVs7u911W07PqxV53J
bDInX/nYQlasOIpPTodiE6itV6rOtbp4WUWeLAjXZ7qwhh8co1QWQjmKJrqPnzeww1IRiQwPnBrK
PfXQOQMwh6qn3BZXYAYODaaUHGwPbdj3ivCpu679FkDbyDeCPKBqboV0yrR8ggxXVajV9jpEepe+
2qer+PpLjQ06klRvTz0B/FAX8gwicYmBVOqr5oNI/nX++3vPZRS3h/ZNSVAOwKhGh8DT/Nc6g/3q
hy/yG1LXflLGvUiCJEnhDJ5iRP7ftBjaops3qQwea7jj9EIiBz2PdvWyqmLX9wq+9IJYyADVW5+h
47C1lVRDFrlF+cQAlXRuooiJTWVm8Lb6ncYQ8Fny/gCncrek6WFXZqms5zMOY34mzKUQLYJQ9CVx
QrG9hPArzzZYc25iQHxNXX8Iw/45ym74krr4nCzZaHqYPy1DFPdjrEty5Mk03Ctb/rNzr3w9HLvO
NMIUgr+4U4R32jFEkN6lWATVblx3RhYQ1Ya+cdEVlxfDsQtycTohhu0tbinP6eGN+Ih4BMOduxjK
43AoMtKTssx0lWQWhHx9T7PwPsAHAjcYMyRgV5ZhANoHQik5ypqNkO9ELkcT0wqNYQed+LFLKVLp
x+k434q9s1gom0mGniQoJQIudsIZxzP7JjoqZ734GGczFCwOnh2eAp5EIRTzS6rbpgT3ukgIoJGe
ELkmPgXT8vw5orwAkvs8oD5ZjQv2jczc3zRDs8IwtxShI2djiQ1pY7DsMdpm6cO7wU5eWNYcuaO+
z8r1VxyEX4DM804hICneenFn6PYcZDWDyy072FwfRjkV3Q6OSdt9hNWvVf4PhwYhRWLvzTjuPFF6
VYJFXAKKX+aXuOeRu5XwL7AQZExEgSTP07sQs4wqdrJA+im2Dc4B9SECFAQyIxynA0tqoIqlmY9I
qEIle95Hye7vuniild/9kyqqnaX7T5z2HNIfvKn2BcQFEe+phbnZc2bgCtLh18wZdfwGk20VDXfi
5fJmDXQitYIwz6PHaVomfu7PGEVJxPQXcuMqOijlmVysotcJeOjebrTatlTnn7o7cxBmuwZKZG8j
vPPXQGfu9fF+dua6sH5c9ggshcEvdhFljzKqrKsNHRyVUB4PhmdRaV7w1hAMtcGDOhHMglZTYFK2
WO+QIFYE1nPLTPwE/GGLawfqGNnGDs+2SEnA/eYVl1NFnyXxpYwEQ/33mNqxf+wmh41XJNcNCisu
7T+QCG43B2JWCXZNsuax1wdHENtaFLT0Y/xPS76/4lIr9Sc/F7YaqFQjhaY9BvKS5jgO6dArFofX
L29rKHYyDDAdyVQn2pNGD4hE1wGDRdz5pPjygNFZe877cQhdkPu2aWzwJouxmjOxkQrtaKl57Cj7
LIKSaOz3KmnYw2ZwX/agCFSarEPlXVOo41Hea+LY/Rg2TzgQr7U3gwAmzPizFmSJ5wvszDki9s2x
OXFXitIiCfhzmS0edUnw3F9CkNbwjCN7H1SsLdGZwTGx8H3VqcptgYn+WHoVsljMIz1wj30xQbdj
IZdKE0w2+mj1AGJPeTC/NvlcjikjIFLVM0P8JZdJ2RlSZZLb9Lwhl4oJXby+jGtyogA0Zyl68vVe
Kdcg7Gbafq/oGqvfngon+Tyb6fz0b1LGXsbDSbUPiVaF0b1rQJsTbPab8MV+gYudYxW9+zcW/zRg
JLW44G+m1meaLEjCMJ1fjwf4BactwlIcQ9HInKj9hvC4N8sxhfsbVw11HsoeXs9uX4/+Q1NfKBvl
DNCnusS5Q1U/UF+furv8Z/EyaADROf4I3ryrwxS0rpx9yUkS4uJumc6qvXK1X+8PzGx7JCCenRlG
zzoNLbksRYbHT5eUhgMHh/4ohh2gKdOvg3lNHTf6z1A+9LbzEuZENGQgXENh3lwZYZ1qQpTDHrvY
vVqHvr/6JXKl525997zEcsYZ3Ph/dTDycXV8+J7L42SKZiSNxP2OArhZkDPNK6H/r3FtTVzTnSZq
30K1ABy0phETv2zVecDKzzv6rEHSZIP9NGwfAO5mEIDiFKUnqQNO3aRrKQ7rkUPjUWbzAxMLWn4d
uC8Z48Lw/ox9M7z+RPFhU8VTLlldmf6TYJj2Lwq3mhIgA2qGFAGAt6VqzDzBiaf8DKQVCzjACYLo
YjAe01lWYoyB2PnyhAH1xNdK254WohSrqYwOMN/H1HUA0rEfBbFptNlxgXmNTxJDEW5I0/E+jnb+
9j4zQEbcxUrZKaPTZqrrJY/vgDHTJDUk1eKes4Rein3AawolQW7JtM3JMQZuEAhqBWIGJ5ap4e1T
q+mgHq2KqHxKeuVl4PeVwMM2PH8/n06szo3e2X51S0sNIJ8dQrapEnRbL/WlRxKZrEvCmB/nbyHY
aT7hX5bB+c6x/mvYZv+W/Zheou9GLBsxDT8KDvKflQZw3oljnI6GO2/TW5UMqn5LZ43KLJboGkLR
CS7PJe+bMVL3JHIrYinc6VSg57KO4bY+xF7/ilgynS5Tvl97UbR6x86KELWKeAJCnj8yJ42w6HpX
ttfxzPj2RoKsgFe1D2MURKa3jVOCNl+8O7Xrj531b6GVbj48PxWm8Dgd2nrmbtPAZ3LMapHkynWp
R0Qkqi0tcjtA94uEgVSVHYrgorYEsM+qkGsnfPlllRNCOwunFQzCFJc8dgJv7EGb2N2mTXS0PtBm
JuhjUeexB4i79vZLL8kdAks3aJQq+aLwoP+UkWg1A3iHy37QB/83FOIid278XQNOGs33hFQnJBUS
Ump8ZjdEeLuRVMq4V1C3q7PyNf+m7eIFiuiUBLbF2FmeSrALG6ea4QbhFru2GmzQ3TKgx7BDy9K1
LxmbmwP+ZBFkoypTIlQr+qBo+Yhb2RMyNlMpyUhi8SglJVEu+YLHOsTG9k7L785Z8yU+Hcj99J+k
ciw60PTQza1dmd26L2bEOXo8uIsQfCwkXS9TkRc1doNp9/nJUOpn40d90kgeO/386pJ7WWFAZtjB
s4QcXrSiXylpg99nQ4C6WyY9pq+jqfhqD9YJKzSip/jx9lsNHvUBiEaM5Cb0oPUAnUS3q5kp7EsQ
fc85exUAglTI+B/TbasBl/Wh3zB9JlVbICptzEMylxEW7Wwr7eEY8Dn/e685733k6tAOhSIlMpkg
ns2FDttgOay54EPsL4e7TFOtfqyLlP+36nOP7+YSEdn1cr/0SlUQDIRZDIidjUEtDbNsTOf1QRB0
BjmtHscgaHDP6FzDumfi/4puKbUUaHjjnU8aSCD8EPKfMnMGvFqw+3ojvD0OVIQkBrkn7v8xj6Q4
tQlpIUK6Bkbi/T7sD5FAaaU54acOMQZf8rUCaajnBWYuqD2XxVxB6MTjy4pUxkBnw/s+24fXnivm
W5UFXsQ0ISBx7pfgU9HOqfJXmL8zSeG5fsuxIzKgNjD+sdqkzFtAPL1JQN/LvDCOfJEGI62CThpa
0DDS5275gnBLBv9M1rJyyQIEmmBsmATjv3oNtqUdUBqlIaQNBVMPYRpPSHGq6Xt8bq1cluMWtQKv
8mADPi2QmYqGOe+JbEeJazdDphJrEmd5WwAQhmG3k39ZJwcEbavE2efXtAxjc85waTG3IPe+S7ls
hVcUIkqUEC8WdBjB0mv9aJYgeVNo5JiNRPcbCFsUOTnvxOej8lhZgTnPs23v/JIoHSdQSeZDnOrj
2eoqhRMVYNelhw/HWRd/ayRp/kUsPW6vPLkQAZiKpWvLNFBX4RBl7efTh/4wmmqhktsVxZMNM7SA
p4ix91a38t1Ww1OR/CIbZFvpCtMiAzFqprnM74tkwX5lYqCaXgMBcIvZYKWmGvSwP4BDQ28qCC4a
ZMosUbeWd7f7UyQRi71mp6D1V7aN7vxP2RVJn7Q6wsw7hMY7TZkznvbfZQeRz4o8NAhLsQK9jsSX
edDpbQu5LhLdN0j+ikXLygObDidcbK6EQwGZGRvs/JwxbjjW02V26xz2K7oLVOJ/B8FFxfJd6kwW
nuy2u0GsDvgXoZ1ss31l3jZEcHYY1sS5LaP3IkI1tIcvRFiuMWGp9HmMZvuhhUYyJ4ZwC8GemW4F
JErVIiNF/s5RYsGa/X8bfoWfyM3bmoOyuoSn5vqGiBBVTtfgnaGp5rYKZRn7yK2KvdQyYsjQDizw
PnVe6jKb/kJ/cdju/KB4xao7eD+Mky1N8fDk6iGQymcIy+3NjRy8wvIo3h65yqwzMLhaH6m4BThO
+AuMhPu43sZ9mqLYMeI6V1YUPp5N4Gkk8dkbmDYEdbC79JirQinmXTFcQqzBXmxdWtLF/ymK/OC1
RPQnZuhyx1VAbpQno6M2gyqnGRn9ycP1YeY1M6RV8VfnOHDPLwhIGSzGYyus74+vTKXIOSYDkYIu
aP/eSLdYdO5G5WasFa0CTovvS8IjcLi+NjvnJd1OfhQkxXm1fRmSABqQEv+fBjScnTln/UGy5QPk
4J+uZPnp4GWukuc+1fQbNUJY1Hz/8zjLwQu8kPvakXMH2YuTiVB/I2w2TX5c9e28bnQDoS+/NouZ
IfM7HU78rRGhPQaa5+HTsmnYqZlfj/1Ku8caaCaHf3eRjqn7gmEoXewMXaOcggMHUOkFlcTaoRX8
cC8gQRQ7ABVoX4ZkWdTVrnPg90ztkRm04DNKQxyKUmQBN2rksBc7zAC0P18Bf0xnSHmKVN7c9xGX
1y0xVR7LRG5oSJ7o8SKA6ZgdMXnJiSoqw08w81NSdQprHu09AcS57ltT3fSkb3BulhRhnqjqFuTl
FpA1CFgGHn/q5RG55jGxj/0FCQsTr4pfxvLJKeIUYSC3rRcuGB0tvqF9+TzIDOoRDTMRAC+74jbU
Y8XokuMl6SIMeT+eAJuoN2EYYtKOSnurr85I/RE6qvpifcI0+0eyGORg7v9L38U0zQjRBGcMh4LJ
foCiSmjP0hzeZRIpbFHdcrvhX6D1Cwsf8HFXHhpYSG9+0t99tvSrbnkNJ1nfuXLBv/S2abslIoTv
yh9QhQ0SrFgCrbpkpW7r5nnI53ytCHg5FdXV3iC/xIEcFSOhpaz+gjxggsz0W06QC2ulq4+u9wpZ
UWlgS+XnuJhQ7LLZ0q994KlQ7ZTQOJmbx1Xcdvkf8gl+N9A+sXFjhAPUHhO1f1Z1IHc/eEVM84Tk
QXDVq+4NSx2PV9lF15JJo9sy5kkmI6rHP/jN1O3AEEoYgj78GK3Y2A6+D8/TzsFeHKHsnUNt5A9M
zK/Bcdzr0qG/1B8ye3lMeYR9xXCqvv0CyAp7gyGuAe43OHRP9puCgE1VJxrYIoPumTUAkhScwFi3
EZGdLzjFeQ4dSiWql07GoT54m0w/fl4DaG0R30E+uXKSlUjfNe+nvNtrHOpaiJnwrZcl60UNHEDT
jMKDPQCSJBm+SiUwyefSw4vgP4+VN9oQccUdQYlc+wqckrNfkGW+VjCnx5gRKT9Zlj6dvW/SaKDK
pfP7xOB4zRVcRYeU4YW6mpWeyYZPK3OzlOUHRD3/XjOB/6wmeVHs9crbK0/zVB4n3EPlKzhM+3/w
3DqPqeRB7GCWfKVxxzIX40IDN7nLk+GqR3rdjw+4sYhhmsOBsES+1GtviV86wWif1MemaRA0uxPq
fF7FNVrt9XT6KYFiAF8PW4r/CeUNYkwGzvbu8FM54tKrNyuFCxvViBvqsIDU/vtXKom3/4j1OvSm
DKF6EO5Pv7X/vbdtBurMmIDPszAYNFk26R6sm0HaxZU7Tu82XzLnkQiqfhMM8GKGPoW5/AuFfjIs
TVF3sxE+21balZ+p96nqpdyRbX6ro/q5+oHMgXhbuwnUcdpJs9Oe1iWUmro7crcpP6i/B8iLosCi
hN2Taqo/JYwrma7xW+OwnaSTNhGrKKPZA2oakAKz0rQqJvMEfaRDDSErl36f66zDdYeTd9U2jxOd
1ov+iMlNa3By0hF4Q8WKxp3akt7Qf2mh6uAHAktCUjOAgFXGsB7S46gB3bWaKAprn/RcBDuhBmhH
zr7ISOtXJzdcXeio1vvpoN1tUWCHZsDPfg/z0tDIcKu0uk3KtVW4/2QU0halZNXcBr7oo+eleUnb
7BxUHwNpjFwuTBZmfSCYVKSFTZJLkAQrKfgsuW9GPHzH8S62m05l7cslUU1EFXoVRL6lbbE+JjFU
hPUvI+UbWhYa87mGhq2qDRE6eWU53i2l5XwoqRd3nSHbkTXoV83Suescu+TPcNDq6aZF7jVHPAF0
6iIl8DM7g/YD+KjUU7sL2+UCNf66EJG1myY8JKvKqpt/pQZX+xnTnjfdaUQMO6/wS5ChWFk1Zu+m
DtHLpmg1/d/GkxFGDN0WDadv3+P5kZQdwv8PBSnvKPwz/sUVq5mbBJgHp0eq1ihVQPcQ3XO1WHaP
PyXRnBmDiaf3dTY50HOpfKCS8npPz1LyD7EKdx5sGy1VX2Gea/uDvEXFB7TgNkccMutOX70OPQ/V
bWi8YRJD6hWc1mnxtNzpNtb4xM0JL16XlkzTWlz5t6OGEoVLmSvM8iLS89TKZoNfJeuJ9+y6Mh5R
UkZnYy3TbnTrB9bOX16UqnmZqrhaFEOEKQi+BmMNLg/cR/FRw5/xt2qUnmzd8VoxFavYYgayAbVo
vogpEkdK+Az2lg6VtH95pG0ZB8DMSZPWV+GZ4rS3t2zh2S5OxVAwvDBjhT3RUZO4nDqdo5GwIkUF
BUm79/PFsvgB2HqKY/zZQ2MkeRLmnUcqGzTazcFM58Yq9v2JkUTtpmxZhAVxyjCeK5SVF1MrBEwJ
E8o9lLLSfRDAV4xjmBXbJCxIHmcZgSt6y783Cs/20sZLYwiAQZjIIUmTyv4cPET7jZgax1HReLyW
sXaXPylyazpSQbceaQ4ff3POWT9pfZ1HRmHB5cQzw/YCnZN6B/0mWswa60P9QWtw43DU7Y0Q0MTB
Nd6YzyLSoYmsyn+0hSt8PvNT0DeXJB0dyv+AMnzLa7oxcxIMPm2dXctHXx3KZ7jYM4VGzUznzjvj
CCuJojT9+4lLtJA2R3fQxXBYE6VoBsGtQpsfbK73wTAfYejDlE6EuEeshUpIemDj6hIO1srYlLTQ
CTqhovK1dpM+0Iydfdwtb2Mp2C9yKr/WUZreCwo7WChk32DTox8MF9l+KDNtPcXieTfh60XHv1fU
DLyhVnzyrFx7YlA6K8Du4rnJmli14laP8y4diJwALmUt7qdaq98YDUB71PPAhBqGQOLDhfOmseng
aHYTs6Fx49/exNsRnF6A55QHgKEjhJqaUFhDsLwXClZHEN7wAr90DWN5mYLAeFT/B7vmLsqB0THJ
OCEjVOHo7EoDG5U/oudepyBy0uWZmUmkpkH2Dj4N6aORj6h0jcFqxbap7Zo7uDYwUJLYHKpG5K90
uATnC3O7NrIrXPQwkCO/Lsywdmn2G3zqje+AqM5UYTQvskx0SvE2qe+CpLAnuzmOs2k02OEwD2D5
yuhmMP8QZuGo86H5nkFKLG5Um+OfRdogZ9qc6WguEdtEbBVaTGL8L3WIBoUSTs2DXbFaUoSqY7ZU
hvCZDc/M1spjVVV/vGW51WVGlJLsJ01J8qMHUNdRYjOe8Y2zhYeeIjyuD8TCpfhSUTGe6uTeNdjB
sCVpqXOmTYdMKNLWjOVky7Ik9kNwvozpyM/CyAvcWeGe8DOIWZp56n51HiK+YvTzmQ0N/vAebhpm
3dxrmUhQ8udDZ8nTWoOzrR+W58c6XnLIVMX3DFm7iNCveLjZ0v931B1TDFCUDYVPqNV0icfDfmlI
ZzT9ph8fqSxuPFSsBqfsnqUVIjaxVQ6hC5xGR9giskZ9/upA1e+GjznOnqee1tHTVQXDUmQQO43V
Aicxo1o/lv1zeauVpdmOfRsZZQZ4mwN5SS9cVHtTihZNONJAOl1HQmT76AJMyrbFABAMI7CUu0tl
3xexJgqoF/v55Sphmpn62hBCrGzsbYAG2kD+lnE5+tR71CI1eD5xu3fwxdsprEa9PCztuL9dURMK
ILs+G5GDl4cpmwFa/b6W7WCJYDHfv8hj2AD/HkOEWxEUs0QInWYImGP2DR46K5d6yroL/yS+Ua68
XBl5RGR2KLUtRuu03Svt9Yt/vQrSFB4tw6Ga/xuYqQhdf7eSJ6adBliHOGFvmO/VGXqb2Ss0Grqo
dCr/d7Q92uHbsJX/1zYMcvmWa3+MsmJboZnwdDBs99t3IhIVO5fpwL5XXO3T5vRmVUqa+YsPhrK0
EqC4TtLXMLL+xNH2rnR0D3nakAHaqOOF0GqQbWO+wDYPnYtAxZxIz1sD45xbkI8bbn+mH/Se4mp6
6z1QVeVANMK5m72VsK7On2Gyc+lhpggR0OEaaVfGfGn+vHIvTbsYP8v77rzHrJLBeYOlfSFwFnw9
ZnQCVhHUSD3roqGX1M/UsZ00DS713J2cPzTUdZuHb3jTK9uHwNWretFOzfYFMBhtP60qyy3B8WVK
PsDHYj9ghj7YinO6YIaI6iRpRNcwxH16nzuztxQrbCY7DIO1Tie7O1KeKGOGmamekY4lX69fcmpP
h0JTqhJFWTs69Av1Ek5HCeNuNou+HL9Z4AiUHCdeLP38k/+jyp3gGgci2wIC2bn2zbFnk0lQF/W/
JW3G7WdAWwaKpwXGZ1x21blMOsREiMrfBX47nYwutOaVJuBMwxyTNZlkSaHf24SvjiYoZ7GNkVKc
TVYvWwVHE+kJgDdRkUDOrgkq4DeTrbt1KxjuHGmY+SvrT13OgBk8UHVkNhrCI7eBmQVaJvapGw3g
fqeHWakElz4+pWMLFA5ogneLbKqVCJ51uNwlr8zV1aBsigyjh1JpV0X9L40kIDbowqfptWmnUYvO
ynRi1OqGBUFH+Q0BCbBZHAtwSeqgnYtwJPTYy2BrS2saoH0A9dL7JOMibbVZubxYa9T4TODnwcff
sRt33Beb1ij0Cr8luSUmIKfFdx+RW6ElZaCl8YV3bqZfU/N4RjyGQCfRcjxYqKY2GPnD8T0FLK5y
EEPzEngwBaaNk1lsKuB77uaiRgh81PjFPMNRV9g8NlQxRU4BAOzN7zC+YW4zyM8wKBC0rdkF86Pv
DAFCL1LBl72e8GvQRHa7PFx8KD7shOHQOtJWW0ViatAv2z96U1EAqHto6PxpE48b3e8Ufbi93k7T
M43b7m9yYLFib0ATXWPKATulvcyDKmVzL7oYaoT9Dc/ty4XUDVZ0y9Uoc+jlRUVlER367DgdwZbG
sDi1aCSvwnTutghiFWpGmphWAVMHkYFKRTqIbmgFg9rYPvIQzBccZEMyGK2KWODCOY1S3worcbeN
pniUjK+Xl598LW/rvLE4dShe1/ZUSK12sQm3oK1t5M2cSzBQTVyTzV2CbGnbXUrG5y5xF79Lke7/
zqhBC4AeebEVv1CGAavvxAMiZjEYXvmZchzWpMEilhkTr/eqMmpAMXhHtLnn45P5LKVSoRwDLFmS
fBpYv+rKQ8QPrQ8mtFMcULmHFHJarAFEv6w+Q/ogOQGwhkpUTqJVKb5u+aWASFlIEgBnT3XCBgzT
78PBeEf4chk+0ym9Vgqxt5hQwey1vAhQn3qsHrlPyspgHiBiLbLF3UtSnXbtRSd6zpSNPO4xqVsA
ewBQvhiTpzTEbJDCBz3doiJVB9cVMohYRH7/IkMrwP/rN/esjUY7jNtUcjvzUxlI3xfqYa6y+D1i
4KV1GBRo+erme09AB9LAN+PsmJ+KTAMLXEjFkTIQtsgPXdj6n7+Jvmen3QDA+tVvK/7j4PKs7uqz
40aX2E+Ie9bHSHYiDh1SHdjG1Or11n/cz42HO1Kc2wNSinPZ/kEhSHFbCSCXutRXjWe2fhNGrF5V
LunrvJqjdt74bh2Q1fcGqTT8ytmSMi8IK0tp0BwDZc01hNZh6xYOLaJVyU+e7mq/VZy+T2PBjd+V
M/UeronoVgwrcI6Pz2+91MhwTE8acbt4ECpGQXJWBq8l6UfLMoQcz/Y7p83z0HiIx6FQFf8V3oyX
BpTLpsW18Zumwbi2f3jox1H2s6zdI6wmeuAFuWr3V9Pa7+3o881C2v87oHl7GYwzJtagp6b3L+Bi
4pN0w0jk0UDXO0SY7pA06F4QzobaDmPmRQ+rP5dvzwKybeGRWaNh79F3wky5Jf2xH7y3v/zggWIs
RuplLz75ndFaAid4lTV3DnPVMXfyJWsl0NvkEK9uHRU4CxwLStCK4g1P4Df1fw8iX9rOXq9HRapn
oDWmu/TQHAK8VkwNspyuevt5khM44EnEhpWogakKgmUYJJ5uSlBpxsMPa30j4NzJpG4NBUhZsvRS
pAJeoXJiCneqaq8GKY2HOKy4e9R9kuZffYUyMqiTIYsUX8GzgRrAPta1/5SZzXuRQIPTDgsJ5Cmk
39WxkaSl6lhB74e2EL8vo5snKOQcezXR4cP50NLyXXeLfJI5yFw6K+4e3gHq+0arCetl4guaiUzG
tPZPT16ACGKVSW7nOgWBIVBn+AP6vuAmSu6Z8ngDmjOsz/5VnHQcUrX2RGOxEM9z0LRb/HkiFEqV
azQT+0k9ollhOiYhTv9yDMMCj7D2nGwZcKsxrMfX6/hVwfqamEUJgmSzsIemCwg3Iojo2BTKxhQs
4KBHbLGCxxjPLw0489gmeCskV5FTVe/2FNdji7gWXRM1wKKZX4LpUlg53m7zsqJHO5mGmiUiYcJo
gGmBYd7Yb+VhNGGTfWs5t7azrAv4yiCrs7sRQY7zms3QPt7aVLfQu+5kOy3WbBBjte/PHWVOZ7VC
Blvs57rBSqyrtLD6L3fY1KnNg64GrwAUEtLx8RklQgZb0o3PrOcb8p2tGlgjFimQ8OE/npOqX91t
HWElffao01KV260FS9sJpsrsfRKHwuM6jBOJBe60NVeAAkIz+Rf9qy6zvzXeDeGADkQdR00QUH1K
l7XIL3vBmMw2oVkvZbXyl38nM8izQBL3Q7k1SrTdjFgwJ7doUo93Qb4BFCsIk9jxAUWsUtcKVALU
kNnJ6zUktT48w6kAT1X8OTk3x11dMRiDEuKSyAPYtVHC4Vh6EC8avo4C4kOcC7hoh+IWHcC4nKx5
iN1SESgLczlxTua9QNoNSVknQkPm+o+7JYTMlXcXRBtNNqFmpDNI+DROvXLVzdu61wFPD/spEm8Z
WS63ippxZdk93fCFQRAB0AaweB1n9eTfKAEvjUTnognPGCibhsCrkju5oDm9Q49ABeOseXurfRZU
UjfKIuaPuU0sJjT7/91odCH4hBDIBdnk9aGbd7qH0vFszerBUM2TtjdE7IYE+q+QKLTQXGLGZipG
wc+xJ3WVQIeXC6ZlAlVgGN0wLw/TGKZl3SU4urRLU3SkUVT1fNdzjzPYvgDHkHAbuYGWxKlonU2v
Z7N4rixKNrmFUff4BX3FzcIA2C3AsgGDkiyHSphJsjkmfwkFOa0fV33Zid4rRN8/XTUcaPxQKW+p
MEYakdSJR/HCTdl2dsUmJQV1Q/OsApoBQyQlNV9JpvfBbTiYz6zbKDO52wCgFK5sA+13pSaM7PKT
0mJRUB/5gyj44wyt09aH9gLTl8jUZl0kXZZNIVN/pPDOkGWYE93/2sqMRrIOUS5KKfLVQTIwvqEe
x26tWCzfPtTXHILipe2RDGwNELUeCB3DdNLu2tAsZIXesgyCLcAevar5QBYuNqunReFWbc1L0NVU
puE9gab8A2x0aZvdq8xkA72auFkfMIlnsMSZqEeHPjKY/5Ojj5C467TbaCA6aM3ZXKbgJ12IEVv4
aqvprxe+Om+0+CboWYLvmsrZbKFTMQztT1DCAQElC7SzoVM/FHHNBwZU0o5nKqEzmzdgtJLIdRGs
RYdnQgGQMUDpkwu8GmVKnua2wRqC+Czzmjrf3Ah0cklc7Hi6jSuXM8VcBeE7yJ6ophkZPMwJH2cK
LaVywXCVMr+BzoZDZxH07v+R2QdXVySGA+9tUoKnUqp3GwBewp3lrKWj2mV1r2XPSOZ8XqQUNbNU
wiylRA8dD05/jLucMzVigzzuI4Uq73TO/kIoJOOLYcQIbgZWYlz+u8c8XtVEZgYPGc16KMmomb+a
Lrg7DxZloRT8zXaGNMTWftOHoAXxS914iOGlbHAo0pN7eP1It1I758twJd7AkoPRdic6EfLFOKej
w3lrXrFyJWqDkcpkZocOWUsGEHntYzzlz1O2/x4sULyQKUsuyGcE8vLwYFg28rC6HVGiOmnG/j/3
y6276rznNofJlv++N+MRMqKt3X7rhTuktw3tJBquKHiCamQfaae7UX36u1mhcRFwGqJUF/Sp+Ket
GmJrLpVqsyxcZngDeW5FUO8BQCG+fNXKVH4nOna9tDoC/UKYeb0Q0jsJE3gHz3ypLNJ/dInhGir5
1ya7vTKFn21W+Mmj5JDDTFlgXp3tKwkVOfCHD28X1el2F/h1+86r/mQQdZjYpVWq9bV81GcP3zRe
oR4OBwCS5QMbjkVRGdNsdFzR7eYeWGTqr+hyGh/mxuynWLLk4bwctfbKd9InUvG0v8BBoqZSzHNG
gDvCio3f4lta01lKcbwd3RIEy5/tf9Qw7r8ZDZ50SkTrHF+o7ZY9o//IOEBb/OOsKlBk5YKWdH68
WgGkbtRtKOEswB4Ng60UYyw/YBCyWgUvB2zq8NOPqje5xnig+qSpUAx3qGchoQ9Fx5wOuWUA4d1w
IL3e+tTwngHLpp4OJKGVCiWenlwXODyoq9d96UEmlINk4bCr8qzzGVRkV6f4GhEzhmtcwDfmixbz
0gzW5yGQuwClV6CXtQZN9AEDc/HO9YuleOaQpeRomF14cWeLINq8SbjXoDz1c6eiClEvrh1yYolS
UYPZRrnKTrjqIONItbdGcLh4Cve1qqHr7kBMbuanJuwg1bSDqyMA41mSibR+1tRuuUrGmy7SXNGa
OggGV9a2Cw0UvDzFalL3gHzEUgdmav6V2AwoBUPxwR5ZeAxXRP/3JqwRWD5UKQnb74+V8E/rfkXQ
2ablOiBRHlqyWC09xncLKxdBPxu9DwblW+pSkqWK+y029Ai4A3ILdGw0AxlsMRyGDA88JcgAsqYq
5r0QO7XHNlSSgxljs4lf6K971D3SXFHm4G69eE0BA/0wILBgc/oH3vnG26w45Jlu39Ij5ovMwuRm
iyLdUFBIT6LmERD1cesRTkJA9D9mpIO/WuoKrJQFrCxagDTpCOo/7JuZ9XTeR4kozXIBUDnoBHxR
g2vOtIM7rQQ2eQBvxUc5c1GMQHP/2f6vO41IKwBgvRX+xr32ulEVWF8E/Q34tiPs6u+59n6syoad
4LTuaIpWWMkKsKRIlMfHH+vcFSyWSx0XSfENtZJnWOjIUueH3V5Lc1EGtIo3N7Pno7y6KN2UV+Wx
v7i/Vfsz+cIyQLFi32MVDOvE59lNQR30mqD8UByEwuqqTtxqfd700nop1Ib3/p6fbQCVKuStuH8F
5Oi2ifrb+aHMZ0x7nQe3oQ7N0xpdYQML1HBGFdoL/QX3qi7X0wtS/Zy6FSeQg5bxEGpvwXCwqFtt
0g2VleaHNEqoei5X2jTmEIKNEk8t9kQRjmVBVcZajn6b2bB1fPbwC1ahrcnsVrEFZ0pQdoM9JjPQ
gGWW6aEOsTWndqzIPpMd6Y7dOpk3JiTRx/dl84uchPdEbNLVKwmDiGeuAdrcM+RMenwqpwKvpyAF
qJmWHDemqhMb9BVrT9w/3hzod0kjXqiSum3yzKgELynONlKHMzehv9hzdVnbW8Y5pi+af+zOEopk
pexsRS/ieYg1hOa1m2QkT2VrPiczSxUzPSg766eT2A7ZGsDOAhze6ynWb4Y3oV/xXsYieya8Zbbo
F8ChDZbpfZIndpY4w500L2TK67R/MuULHG5c2wgSQEZiVpFHJb7B2YuXyugbpQyC0HRl2G3w062w
LHQdFXaAc5+cd+xc6FrHBbLKIlAP1c62jxpqxRoHTM18PosV0mZd3KjelnSzkYj5yX60KZ4T66ju
FHkrIVVGcC1sqsQq28cxDMBGYt5sD1GK/icCGMi+WL5tEbWGWxdwhF758U/ddyHv4LzOzgJHypHd
SlePET08MOMi68JIVKP7v7bQDNqSNvh8Vvht6jRXR/rOLAGKA0uIRc14suy3vmSNPwZIvh606knU
MT6OTjvk6465WY7RUCD6x8fZNSLVY9eW60eYblmMKncRVBbCAmR+0037Iwn3/X1nGDUFeaztRGsl
cz8o7OOI+g5QHK9ozs2wOTx/f+7d39dy4DuA1K1a2k9/S1L0IBF3P3yEQf04AUk9kfiMWDxjplG0
vPKADCBeFTolmyo9F1p05r3YHpPlBa3Be8dhesZ1RLiNl2rp0UMN6ctHJnOCYQ+zDuLKgDfmCGRX
Woluhyj7PqqIfZ2WGZgQbIJRY/MpC83/5W/+A7/GL05wCevA4KGf7/S5H1wBlrWrz5t71VkzyTQT
idxikGzvfifrgMVVHT906evZgG2VELUqmpgUy/CmmTiGaNjAbSAeT1khx/nkPLBjnjWuRsAspc8s
hhTcv0zm84KI35GTNe1gB0R3fCZX3VeZX4Wf7koHs70XZQMWdb3aqt/tRCuPTMwtZPEeWw58Bhyy
S/Ywsx9GmhbPD48syP6DwYwEKBQQSndexZGF+UuAlPHli2BgYwN3owRnWbQQsVQz+w/XvFRpcDNm
YNwMfP2a2WO9XLNrgkBSHbetzlvaBnjyr1IcZdKsCqYGZTJwkWwj3phcj5mtMaosqUUqsa74/Nzv
MblZUzRari5Vs/7qMHLq8VA6DqFNyru07hejZWc42iILCFihs2BO4RuLci56YE/UKuscz+be4mcg
5GakDaA3F1KkifgsZhaglS4Asm3Ye11kip3PRF8uYyVweRE3EXVTnf80l7p/nv92MJJXWhb+Rzb/
cLVQJ7HfBBwbMzE4pjrW9+nTXqhV8Gki7yNAvWZpN9utrJzpBxzVnEyVwiB3cBNqMYWNYIm7iFjI
BfU04FVoG3JZnci/cR3794QMS63/ASZl7aBC3IgcTsQePASsVThpP6EUOXSdJjkiqEweK+fMbWg9
I4BWigg87GY0XawprNB4v2UPeL6Zah1wocgJTFtMJzRE0XOzDTujE0nCwUXE1gksPYb1FbzIAjSD
LpTN8JKJ6rkY12suqMRr0k0fG3XAJBFAMIxxJx2H2QSUMCk6tzZUOSd4ieaczg/J53WKehUQHtPo
V89RwGCeMGlh4r1V1wl/LHveYFvi0WyCFpl7006a9LPvemiaIdiZnZzIEdmMmGXLkqiS6WDDKI+2
rmLfj7GHEh92HvUatpAamcbSsyiPUJCxFIgouT52Hd8L8M3Br0PIk3KfyJ1gNc5UFZ5XSXQ/gMfl
e6mHNaRpEeIouIbUp1Go9AWQU8cbSbnpUPh4XHpNhGyKIzzfJvKvCX1aIJPK/yWoZnlDziP4JWSN
xyzdhzGZg6Yi0pwq86fvBjCCI9QDyaI/jiLvRCu7n/+mZ1/iRcjGYAn5OqTqET8R/neYeNgnmQDc
K6UB2OO1XL8VanooWlSoxHaG9fFoQGXRz9rsvG6lUfYHpPt2kLRbnqOtCioSrkHoLj9d4mDlvUH6
S0TgdkA2kPp84kGh2DSLEWuaGlgPjPC12eSj39pQ7fPml1cYkv8bEQfFU5NsipLi50fD6wxUH2zG
z6oCRT9MAqlClIc7bBjV6WCrUiz5Wo5gS7RmTNk8wg1PZ1EAvxx47DlkgrXQK5J+837A5rOVe1Kj
th/2BjHrUH3rMbxVth8FF9cv7P5ePl7s+IMLL6nuLMZdybUU7SpyvL1z3hz3E823QTbnnuqgdHSL
JIjdhZwxSr5R+quUjk54vWW3h7XDUlBK4KJwUdCUvYfXPY5QoCDFfWe2fsGqkgKj6iaug2sj/OEE
C+YveN0QRvq9DdcAjfgCmit/ZHO1Ez5+ngDxlTxNMqQ7wEGwUCHynkEpErrzDTrE8p/Ma/pUMcmD
JGtvq+z+H7U9N1Mfp2RBLrqDtOJvAMSpkMMT1ihEAlgXtUIAWEoR6Jzl8wXJPewYVV9KT3+/pVW0
PpePbfNId+DIULjaYK0TppIXL0vMlaf/nlvh5bp6GQn8CoCRYNYy9RcYR/G79VJTiAzZc0EG0q4/
m/nUvdW/iZIC86yNKWkR6vRoJlGiEchQqPsTbWdKeIK7IEApM1QmenNgcVGPtTYPmrHX0zH7PUjX
GvDNlGHGB0tl9SCN0fjzpIa3KMQtyW41JLC0/5oAfj6tbBt+n5FkdmRlIMd9/NMI1XcMyq318/0J
b3cslR4OG9lJsu6BZejcKJqP9mQ8eyh+bLb3/REG1k3RdOpKh2UUdT9MAgqeHEkmlaeiSrV2X7b7
/buiNqOMQmYGa7iwlcOM2K6670jvAAwjTwXqDj3PY9Ujr9/1ePV1Kk5SosdkEdvcDRAbBV9uR8fZ
na5eCB9aXJKw//VMy4RELM2F5dgTBbOyZvMEAzi/dhxYVbN6XwhhwIdTdvbZKUwqcGdyHFja1nd1
8lXoOsuzlXoc1LISbsKNeMJuhersWJWG4hkiGBZJdC0bscpLN2iyfbx4MtUM5hcY8JMeHON0L343
m/sCKCqqdX5ZAAv8maGycegAL9kZu4cxiHdGVNGHEnJynttH0ZZHJi3nlBOqOMd0cr8ZkNfUSZHy
qJ2EWYovltcr0l1iKDyMVtq8ngEP7tZXekoL0Viv0dHkmPlXDQmnb8iP2G0uqyJp4zFqDp4Wq3la
0+F3h+NZng49ItqReGX5Tm7tqQDSwYxdPG+1Ql9b6nlRSZa59B3qwmQPmc24bhW5bP8kTBXJLopl
M6lUG8cTtuHlCfXX3Z92LeoENLTYE3nf1jHx1xANrqEHafem+DkpdIldacrRLattRkL1qDGc1wti
d2WObwLn2SUzxLXJ5OhITbU7kSNgfI1E7C/rgyMbMrexXo4qx0R2FcKgAY+U+mTzDr7tsXU38Yop
utUdqnkTeNutibKM40gjgHaT+PNVDoi8sk1t6G3CgcNvrdCFUDAzin983F2nJcGhen3TmhWUXNcv
3oBdf7r1fOFIHahao+bKY/k/kEK4gKVCkYhbiPJPcCgJ2lop7ud5Kx/m2oSvMIn1KUnY1OBe7cwG
Fy3z/UuKjS0lfWiliEzsNnI824Cg2JxmvgZaMOuPsgOZkPVeiqYz9k2iZWinnS04yYVFTZRwWbcF
CN1cOAhvBLBNZrIenoH+gYqUc6VlY6OJkX3A1QapdOX9eCGii2LfGvH6ES8paQ/Hk9Y1w5V+xtBS
n8Yzbdwze0IrHdSokeRjzoqn/jICaFN//V07bm48Snd3z6FPrrCvzqLnjoEe3HfNkTmZYNZ4acoy
XMKqJGDov5wDnk0Ic43VaJmU1xpDo9uZKXKNOAtY0AAOeMIG3Hfv/r+40ScznjwpE1W75AbccZz2
A92VK/SGcuTKyABuGcYyFtMndkPZdBZL2M620EzJqVIXpARdVaf+GSKh6zRe2P9sL0zFbBoa+a11
TQ2JEqQtqtqIoNgdgS1x4WvTi9xIQHUEqsawqtuZmv4w+pUB+Mpvxnl4L3Z+gHtcBOR5LtGcPUD8
FxVrpinG//P/q4lKJrDqIBIXFkciImUJn/y8SURpP035t/ojcjb1+3Z+UU/H5m1kif7o9jG/fkH6
2Ng3Y6APy34l2sw8fqD3khTQsJj6E1At5FAJYbZt5adHDC3JAT+1Wlq9tCKBdsNkJr48MOrlL3s7
p09uvj5fEJ6EGGbP0qI/S1PL9mekolixeOgPl9ii0uCq17s3lq0r5aMsndNlSd6syYGWka6m/5XS
uWvtb8hYZjcMLsnAALWzf5Ta9LkUrUwvVHfyV03zgNP6PCTUOu4TsrXd38pyY1PCpL0LmfsOZ5I5
g8EcDqfpJtnmxZXKn6inOe/U6NozCEf94qMd7qabO5mU87/Czxz9KuY+RjbOIlNZ/IBZcNUC/zJc
8TN4bSw0oV/evM+I5MpuhH+1D9fQsrLR03RKKtVxHBPjpJPJMQQNs7jOCkMXRdFuPQXNz4yA9fVL
Jzfoe6d1LeWWpzwzfQcbjDwEY7gXGToTeqqB7MoQqPs6Ph1RooKZwqkkk7ud88AcaKeNIKn67sVN
gbF8Yx4qtgrx0yTH+tFPUtMpYCcSUrSuP9Fg9Cy9V7yYnSwRtSBGwJM/71ENMvm1wKchOVcOZph3
8cHpGfiXXoyww3cMXbE+uEgC5K6+xLYRHkhFsJB/RNKrclSXX5Lx5tf+qMi45tKqBJnsh4RUqry8
cMmnzF9351lPkJLQoul77VQ5afGvebfNAnrowfExxcK/9sFkPSY6l3v5Ufl9yjVvlTUuMiqKjrGS
/WAYIEt4Mrg1f4bD9WUYS5/tTx16TjCd0eJKJEI9qhCr9Ok2Wi8qwjbPjfBJcGDNpTZv/FYBCA0b
MZdLtNs0bNUzqWIn316p+3oOpGkotOdD3Yqk9wDFuuHgQE6qThFrmbko5BQeW4tOAueAATWXSM1j
GZPO2OihunSQbsd2LQyfZtN0gT44HVJlPuwI4U4fEApWiAJipHBWzttdz8hqOqrVUwDLCmIrnLHg
VXndf/lc282K7uanwpPwJO7LApKV3ho9iaA5pQ3Syox/Q1hZkJwxr8jqBVVOpqQYYKMKs7QpxiIu
lGznl8sXpvpuGVIY2hjLdCq/OWuH+PFvWIpOcQKUj6CyhIoLxD0iul0XvWwgra+eLGXyroyy5FuD
zRmyaR6dT3p9AZGNXgTme99wY97cxzhpeQ7wh4b9YaxQrOU1TOrE1E1Te0fuKVj0KY+BC4uR9/Z/
1gxP3KgPDb3xSnZ1z6IMH+0Jp1tlXbCXe1jKr4ZYsanG4zwBfec7bIzcY6qwKKg0hxnFWo/ClTKb
fxpiGX+VvNWbUseRabTiaLcBwToToTvVwCoyIhC2GjaY4bSkcQZi6Vhuyo27C/E1OizfsBDGfLQp
vBzHWfk7NNUjqxXstwJZIMZd5+I4GbyeWcR7NkcHgZ1aRXOZrQYUjy1FojtuHio/2XiN3nQ7yxPm
VyqIy2AsTA6giB1nJgf88SXTokXk3cLSRsNpg6Uy1bJ47wbRABm6Lrhm6QmgvY+fldCaBj9YIj+n
HerwNcOuVKHh4HWuB1HoIVqgXEN40gFG/uuhT/uD6byrc2z8cCsee/sEYjmUS98mRewIifHBPdFh
7m4NHFJnKDbOxchGHHt+necpymrjOtSCPkgEoOk9TiscSCdaK4bp+UCoymnu4lud7Wb3HY7trMMX
e2qyp53CIz3qQALp0d2T2aM4INc7pKLsOOFYJvK05OsA5ZAt0jLu86A+V943oSkaC0WzNxyIBbcM
jn17jBL0utU+lgeu0Tzks83TPFB4kSySne2PfUPk9+PswjIObGaBjAu+hX0VyT1mkOUK4pd+KHcp
ZYrEwfil3lmIOOUP7g06DbjH1AW1f220x7Xmel2j4u76gem7OzrichDpNKR6G/nnKk+jJHWTkn2i
OrhDm99NhrtBZXZqNqnXa6EkOgi9VcFuTkcMAgf5hF+oIfXm6BbnCxF3nMlEAbQpARW90dkFz/XR
y0V9y3leth5wFcJmPpaKmwe4YKSUSWyrU9ku6LUfGB2T+4iR/kg+iI7NrLh5A8KiMPaIbay5ZYlf
cimOQlu1hbDPuaIYNe5px6s2Nqq3UFUfeoZqEKO3Ad+XMhSOtaFQ8CGPHH1RlAaOYFzstvukR6sy
KkaI3tAwltnJevp2Jc9C4hNOkJ34k2j2tMgggXMUjBYqOyIk6dj6lpd8vR1vyOeUiWY7ksUySUUF
1HEjd7neaGh9XmgI1cxmzpETWoON8ZWhxW7Hmjju8tXmU4Ox1pTp2eUtIDAT8+APYGUKMdhbZEjS
NSZBqPUMpU7/aMTYrSPZJ26O0pHuXaOtHtWFUeA8enOB1Rc8Ikc1ksrW1V12AHsfiQ73KHqGcrVf
vsY9f6BDtHfAhJt1iVBrRZ62ofSXTTvLfMTxmQdBhqZo+r298VB5q0AF9/AfiFDv51vhaX/DQUua
gb39c2iHngqXUyh/XXUs4wNzOTZOP9kfC6CyOU3Yx/wYIUfimZ5OiUxhpn6ihFXUiTNoOzBnygbM
K5x1RnEWBzLv+73H50XUyxguSu9m1T7Fy8OyK1ZYxsxpppkxq+UJQ4Xwbm41V0dp8w5Ffe5dq/A2
GHqGluQ7q6/s8gL42Vaa/FtGFgWDGaoPw25kFCtn6sh9KNAcA1i1ydse/tfiaCt07VIMoQvWMweb
3T1BkZleldFUAj8Fa/hCGuIvXreZKcpHF+SIjIPLf5itowcm5MLO+93hOWarLA8aEPo8sXkAiYpN
5yBL9Xgm8iT2r9E2s3BKbjNXWnJMVl9uNjoPW7zmJOJ5M88RISOJ8ngsg3W/H/M0DuJhSkM9py73
2AMp5DNWdAXM9TNj1alqV70AhcFIPO61jmJwj28xkYxdPF3dLfUWgfXD0SU3IiLuh6/c95mKEfZd
FbysySfAgFeiRsHd2+W+Ir/GfsaSOA81T75neVG/fM0Pv6nvgWkM5WW3LaeuuI2xm6J6USeA6eDr
Tupkutr/L9PHzzlipdX4n5M1Y/YYqTYZiKcDPU9V1MBjwlRIp7vG+Kg+jfK8pNbr54gcwkjItezk
Jias8OEl0RBNrPx5bYKEx+EnlOshhO9HIrMABUeYwSgIDnLgMX/gQC/9aEMyBGr+1siFYrgD7IiH
wSlYFqubK6/h7DgX6l0uFlUE5PZXwUk3/tCmQEjV4SmWeJJXjdQXTNdCdoUYETr2+2/suDLaXUzZ
/0yziLDTGg8sGLOVdhlSbM8SFA30xZVQ7Lbe61qygULsLnqf6KPJQIqPdLWawGRpvcezkckZjoym
qqQFzECDbkJ1qdx+4j+mghSVo9GYtLlQkUtR2Tk+Xh9tyn2h8YAXPRpVepnbYFSo8OuX9NEh/V2+
G0aYoLfjzeFYbo5A6vObyy/MCULex5Uw6KZ5huUqaoQ8YCW/hus26g6A5Gp77mSOe3A3XynG2vBy
xDq4YCmG0Y0SJkNMWoCYQtcj1EQwdQ/PDubIbYIOLL9IULSZ1IdjpahsjPTrRrj5ce01fker6Uip
JraaDXMKIxnvgmeuUPXMP+aPRnlVh6zwO2nS4Q3sqv+oI70a1H5b0AeYSpJvMkfqrK4VTjiCJVF0
C2h8w+1hnhnzPkR4163YTHiOt7FqaZiLEG/DHrV2N3VEvEF0KygVPR7UhCnlkv4D5Z1tP1MKCGSA
K/Q8IW4M/+6tLvffh29xFXioRaVdNEWxoq8IVRyfta5PDTWkbU37wmK24LgD9wUBaBu4rRFL00M8
W03x2Nvq38JiyBHIKU2twMDA+5pTvPlQtWaboMAGnTKPttVjWgmu00os+wiyMUZc1iG79w7LL7wO
/7LrHvaFFIGbCQWGx0O/94N5oNu9wPV1VVMQJueRPG/ZbaV9B3pghaxRYTClRiuWv8df4ivctdp8
kIX3lYUSq+aH2dS6/Ef+/EQ/aBWIWrvwsww2Gh/K7vWDLb8OKfC6VIurD2tX8ZVAuUal2f1dy3K7
OrPnpySw3JGP8uN6MxfuRLZZtwqvHHAT1RuDSeBlbpByBBR13NigxZbNug6JEvfZOkNHzlsYsFPG
03Go2iRSHBpxslF6w8XfxXe9cWuJv5MT1I8WeIunuPSZvVluJfE9EACkFZxIJfiTnqCIcs5pi8Vx
Vilw3KUdLkhYnKUzvEGhpEq38+E0ovpt8A1qTiGLYXQaRTVaFUON/ok9Piz7FJ0eWd2yh5ZeBHhP
64C4b/y/0TUBH/Zykk3N/np4N5iFrPMUofbPYS8kX34pAWcCJsq6oE4NvHzjwFh6ZadtRn7qVUMs
K01rVktliLajhX6z+dPZof45EAGSjDpK8tR4UacEIicQuKvqiHlt7eznN2jpbdPRkVsidcqk95ha
PjrFyZ1sYswKGCREglaJalCZo1cgmXhQ7sxDnbXYmJgmyeE+eb6HitEsHwCAHMy03fzVNZkaxekn
NR2nl8yV+1HGFbL6iFkMcXTQyqR+Hz7vhXhaSJu951R1vR8gfniCSnE1MapmLuWk8B2jaaRt9nUE
+ZB5ULTAK7/vE2A8ZiFeyadh2qra/bOTsJPP73imopsFEsShGsuw6rO+yPsnh8lB1hMjKN7zPTfN
VbDo1CZy/CSJ4J4lA+MVddnwTSzW4WBNWHeZ5yC/B0bXYRlcfmAGZLQFcT58HqXGIprriZdA5aJn
S02rbg+8mrUYSjRH3kMjLrWx6ZhRLtA6vv3fq34Hz73HAhDkNdhhRVDfI1oLGG1xjqJV7nvLCnWz
ahPlDvdlgXbFQXgYo90lGmU7qyzdtRv09YZ8O5iKC73uuDahvk+I6vMECUEtlYzQLFQjvU0CI38s
z2WPH7kdlHr+sFJzdjOnr5C+KgMiOt6Q9rVu3Rp9QUkclmriq7FeSNWgCpQ2AXbrhIiC4/1XZmle
y5F+SzALnOSLAhFBmkc2bTB6K7fkhhv6jefYoziu/UHBA3gXD2xMO48EG+W4ZHgTvOkSCPulzLri
pL76YZlIu/VsWv6TPZ7XSiBIEKmNW+dXDdEvA5HVDw9Iwti7vf8oHL6/OEEWdMm7LdsWrQ3jnZqH
0Ryj8vZPbfIXlD1TwT+EmpMT05vM8nANchbvqle+BDdwCApUkMhusmBqkG2c/36S2Jg3sJC2pB8K
J70Y2FIC2kzPK/HY4gpFug7Wf3+2fxOoB7AyutZsWFFwC+IKKP1LRibkzjYctzB4iM0BT0/CAsje
kvsTOUCbw1eDszFh7UIhYdgwGuezzrPXwoJrFdmlO4CGX6S5vb7SGabos9RF1VhpB8TwBuSyfLm1
tjYhHXFYiPfcCi/mx8Xd1vEdokwV1gH+8syhKutP+yObdhyJ9ZbNpEFL2QV36whY12hf0GnJY0FZ
XDZ7L5qqk0akui8T0HYBheOFCt1XW+e9DFk5fSfalC8X7/gm+oYb23qG9ZadatJDb+xznsi5LhrL
HQi0CXSaMc7RW13chB13NAur63wfb3NCycBIibW88+HKFctErQxWLMa3peSRlSohfHSXLrZO5vGb
dgk9mIk7Z0dW2EPXpPkEPLwX2EDq0hNr0IwI0i6yENJT7P9qBSKpo7XwrecKpfvxHxfNYu3fc+pb
5uQieDAVnpV+p4PSPvT54C1SAdWbD2NZitYiujbPnXA5pe/nMRHvAp/k0GFOb4I1jha24fiT8dqo
RqSvYS8UuxG5/Dp7ZWuUruIpETjqgJmO9eknlzufXoibvsHzDQvAoOSl1thn0TI2QEuR/L4H0znm
XgGMHKAOfuP4amcOoc0Uvt3M15m6xz3v6/UGWf1zWzPSAkw4T4W6xdOwY9w8RapI3UPJHx+z7klw
oKQ+frJAaj2w5GcqCd5zQzMSVmERtD0+XuaA8SyYWY22tbPIe4fJKeaUTtDURFpDC7ghxGm3a+z4
qAl/Yngfq2P+ewOJll0BXjA5XZ2CEw8xakNSOqFhnaD4OzSeAuW/HppSNCpjKFCxFVkkRhIArsBk
afFltxfmxuUxofJvAubHzvzO+Qm2czfMHJbDHw5vFjjInU+1vS2Ep7D2VQjbqdFAfT4RbgKmoymY
lxQVmIQ2kmI4RfnKH6QA23UgHbuV5qMIzN6GhWLlpZQV28JWLwsDOBSG95s5UXRBlHrSayolDR7Z
Vw+LgBe6TEXtOqdZLtTKgqaSp/Dn/M/KjEesxOSkmEUceQ8mpOf7m/WpRFRX6g5bvzykNIUb82sJ
xyHQ+zo3oANLGjYAgvBIhrZtiE5e81op9odwwa1LxWYc8+yTe96txsj6SEQmS2EX/WpdTYj1VkjP
B9UDcwzlNZ/ltho8zlPYt5OhkXbCcBQzR3IVxCVkyDff7hZezCP1xOqrez7e+xGL0UCJMsBKP3bC
2gslCQlLv7ctZFs4fWhi8nwNkCnCe76LzO7gqSvszqRgzSSAbKu79BOnU9fTLxivWS2V3hYsc2FN
Y+f22L9adjYIAZ/o8zovc/lwhEyRRNGnu4L/3owWjLnLEjoXtGNGiw3DyV0USlbVrYGIgi3qxP9y
KVAtZfia4XluDtXuCOFqaYkzYETbl+34qZuMiJDxYp7V/3830RIDb+4FezimgpOoa6gmkHeWtcpM
rtw8Hr+IQHxawV/rJ12oApEc7v+uA8EbLKCJdvu7HYNUxcGu7uvrbBzb+pZRXY6Qcmb0EXhUYXJp
7bNKp94P9lQLSUUeu/BMPYyFmMeexhgwe2cbOFjhVF5DWVisttUMD1SCyaJUnFmHGAo66HYVMmOT
/abGDhfNkd2qXQ5wLFpy60jqZzgJtzLnZzbG9+FAF52KHFuTynneygc0t5IKcUK8Zq909R2lZ8S4
XJT6ZXfXkuubFq7r2wy+KgE0JPlrkje4S0xHkA9h3nzYYqgU9PQQ6c0Tltx/AiKsBZ+h4CCVHgq1
IdOM+IMQcw5qqTmDsqGK4RK+XR9oJNt8DRCMnPTH3OoquJ+uepvIiWbUbj5KJq8Krykg8F/mG9Su
fEdaicNAye4W4mPP4eIt86anKoKPAssXMlrulE4ajuAj+wd6zDjxE8jOq1bpiaOkX96JFJLEgCH8
9mwdI2L6cPaUgtdK7lG0uQmD/3r8u2UuiCH5wiZriwaK1G5sskAY27wYlhpj0OvBLSJzzZnsrVSz
aOUS06uiEvJ5kBSjSQASPRmwoB88L5G2MhrlJwage3nN4ucFwYEdRI9wEnGfKx+h2WaauGwP1MR4
JuLSyaYowQNpuOro3VlYNULu/3DNYMGV5Jfi1GWFziDP0z21Yn1sUaNUO2vmf5TU8eUMp8gkoLee
+RdxIpkZXg9Njj28ASq0QmjoYMwnlXHUt5wYv14ahwD/W+yIVOtkQ7PMii7q3FPL7pdiSWnAe1X2
3jzPNUmd6KH7+sTwiHiMFEXvOrifMSPq81ae0TbsxHPAXEGe5pECj038B2tehBb6zD8HauAIhCDh
s4Ol/O6/cbMxRT+u7DaL6tAljDc9/5L0lviCKQDMe4is2qK6tlr+ES4gjaXVof0ek/DympqgvYo6
1d5DDaSpk2QHLl8DkvCzlAkoVwDLBRhglX621nXu/kZcnnZCAbot/Mo28LAOI2ULuqenpKZ1Z1+y
owXnlH1DF4KHe8m2BtVrncbfB67QJt+HS1HAJwmUAtp37MzAMjb8bpQwfmCzQta8LS/JjMpBMb6Z
e/9AGxb2Q0VfLBMTwwKyZNQnKIQVCJj+W67Au4Ss3L2zXVktVKV9+XplutgXKaXhkaDT62ss9C+0
iovLwilDt24hPTHUjnxLnjXnwkdluLDdEJs+8EtO3GFOP55Xj+qO4h/UwZBaHNhRCRLzhcrBwitn
xrc6v+Dl/alNRvKLecPfqodsyuBlsBCPVdZ6k+O5A745iKqXtkGaG057Qq4UCVjMzSfldStsEoMH
f6nXmKbOr/hskEiGcAbJzD2ISN8k0jCUnb1uj2m1vNtj2LnMG6zZ9nbkkT40yrHcPw9W27eBkE4v
9GiH4SoVRVpmnoh4WzSZlL46z8eH72XfOK5m0SkhbsYpbSTUVrSe4QGLbwwx7rxUuzQxMjnwbFGD
Pxe8+oCtKX8IOJZjhjtLYJ0AgLeddwkfhJIfg7DHn5dI/d6ta6avPmoo2N+YM91EnBzAw/BWlgV9
YYahz5Q/8adcPMsDyx2c3KkUX5N3SOhxhotsJFeyxhE6dL1nsdeGFeAh4oEhdQnRSOKjMWtSnnkw
NqdzfWRjbg9krad3K5YOgVXX2fvOV5xpzDSLgvviX0uAn675QHyrdIhqE7gb1adNasN0hGwJeoi+
41HfLh2xthPSqqlEouCaMX1sh/P+qwDEmG0ryscjvCwYUupbV/xTK8dFopeNPKxKPNj7tSLfWhrJ
fOWJ6BebQ+aDGirVKgkTNt3Zy+H/Hifm8wquKnOSB4TY3ToRyf585t5evMco+Yke431YXh/BnYQn
RHEBW+R6VZjw931ZXwxDgH76BOUfX4grGC8iiZPAyrCvUgRMTuaawPhnMuP8eZ0bx9DF8GTucK5h
8q7ntYmycWz8SSzOJF2RhWGGJnnrkl8QVO/u5y+/OWBTPF2l3bQ2ZK+q+0ABCUha8IxQIGIBkmkS
1GfpSTdOU2nKIEGcwr3VruwhrpTbWTLaX6Y447ffcqTxDUb/dj2pgk2XfDDBLBLEM4s9sBIcV8op
TmUoF24dBLac7g9ABAGTrotP4kwXi/luWKCVxh1be3GiWuHC+Y7Vu9BCDKluQOktxdGtsuuzi8Xm
P7UeSvLVRSzW0NYNG5D9hI3P+rOAuMYGcRzYSVsKwUBd0t5FifATFX6AE8+FaD4w5wPY/+m/+iQZ
A/tpbni2n9I+j3DXtl0xRMnJqt4TVqshKFHIOKz6VtRWdDu4zppR/1T7YAodRCl9i+a4OxswOfxq
q5y7B91ldZnfRZpyAoxK69F/uy32oESzwQv6ugD2a5OdY0GB40ib5uUxahjZULJ/FsD18szfLraN
wdgg93iY5NgnClDwzcp3FmIN5qE6Fwjvyf/dUVs/OzyAbihmzX4WSFFNMp+3gMyC44UF5Wfwqbdi
n7Pq48rJbu0Y4LwOZsQGCt+XnhW7lhGOBDlNpo3ElvogixBgX/ikXvRUb7v8jMPLFiaNf+PK9AF7
or6zrxN9aLLADdbsct//hSBO3kU/Idqlzwj2XGo6yvN0dJdXtoFd0euC0lo4/A/y4xWn0rIl9w+c
T+Q9iBEtjg7uc/OhDxMKwkFuOgkgfDyKbh/LUVoxls9fS6khdEs1NOjFeRY32wfhAqQfgLv0aHS9
xZWv3akB4mHT15Fx1ONgfqkaG5Ex7flHUfEdmWE+GiUTxVqpuPjEeDfIJho52kCk/eGyc6dM74B2
p7sBijZJcd/9Nwo2UjZzmCjxA4RekUTyMSseHO61VhDgmzvpAKxbIFNnuSnjRQhYZC4t+//9aR+C
581laRKzMhIc/Ag4k4uVYhYJXjobIpQM8LW2G+ogOf0Uiz27YzuMuznv6pUYB0FTzx6m3KwrU3OX
dwcHVaLB5Ki79cVHG9vPzqdXGbKZil38CLxInp9ReXSmsADv7MiBPNq59U/6Gs/NNg8Y3iDwzXmg
C7HhBFvcSq338146Rzm6gRFY8bD7NjtLhunpV5u/PBAs5wiCG+PmLpfkvOUwwYyvqY2XVQkn8Ojz
Zh3pTxx3S9S5eFGx4mUNht017xIfG2NR9W+0/a0drk3q6JyeLwAG9hx/6PUG/9f5Ms6wxVm920Ma
/1gjXROLvHzVdIv+mS01e3QuyCQ6HVhUuXeAWovUnkejiIFWNb7N3vb78Gm9JtCBK5fZdT3tKy8R
rK28iTRTFh5MaGMjvULdar+KMqaxMW4zmcR0Jz5EoxDOtIz4a5ZSF94K1X6VYtK9ePXNMZPCy/9T
J/Ja4izsHVE2yOR6zNEbWq7LIEYfHSm/WFY56Q6321ru9KpQpf0uOw37gArGW/vM69rBhR4SiTyN
K5aiXUJRo2gcHKUNcxU0EDQDx7pMqvhbMckNJp51zGAxU0FMNYAAj+69PMfpJ6czxrU2rrI5aKf2
PiZy1TYi1sC6oIWU0rsmn65Q8q6s7pr7iC0BqOIlzzUbchxonr/a462DPgX3OXm8WCWUDWKhxxoG
9dj0y8SDtAmIGvyOKCzF6x70pWHa92xeD6NuFdOvuJibieUuZyH8awSBySTdpCxPQL/WPOV8zNep
6VajxYMU5bAQR9dUE15EkJdOFDARSuqvHITj+nGtoWB0h6xmGLplaS75hAr4Bjz0+3AHDNizkWXb
fOMrgHd/ar+5M3j9NlSKrQd74V5TEqhx/xOkQw6k0zpZ7zD3Yrf1TiYgbiWu4kiX428Sjzmxp+Qf
1FvcHGP3STA1p7zlkNcCizuD/6TGmhyqbHvVqM00277dkBU/2Y3CSWhTZLvHvj8EqdImd1eEAET7
LuVyrrfCQL1mhTOSIey5wQhBOrCR15NCa4ALjkUgasuJpMixXiViC32tUMKmLXgHJQeAO5LHxLHP
h+z3T46b6IrkdOcWYKHJBSQzbHqMpLroZ64eetK2hMgsRpk0UcDf0VGTr5BbXg1nKwJHkiQhW2/m
USDTcoEbusIZ8MfFdbTbPfPL7j7lRRrjn6Q4W1wFfu7ooVusDt20puJ+mxPu1jc2GA48quYiSV5b
D2Snvnoh4ASc+btFzyOyZH4AbMt4KtF4DYPLkOomlJD1RRKlA9kQUgYHZoyhmmTbdSriNv82VrHz
Dmajhh7aD8uM//aSwnc+f9nzZa7y8DExqdN0rT5sjyTyM0gAfWs6t7cbcDeMn2FV+XTnZ0Q+Hu4v
6jxGlUDIfZ5gvFVG5vxqyez/ase9tZCfcXfiYUhjS4T23IkXf5eoxjEjrl7p//RIjX2ajma5o8bJ
dCS/lUT22yvjNHiVcHp49cuQ1XT5fIK8aRNOoqUn/qFAxTNVcdw+njhERDtca0XevlrKNv0si7zG
61sLTkITOyMoV5iCLC7FrUwo/HzbjvyvQVpT2+w5GeC5NDlL+K1W1n9hkScAj5jKykS+ax3aoGcJ
gQ/1eJudU78KLejTburiaabK2Gz97T15JBY/oAVwQMipoWEB/GETDHJOmsP35Pj+yi+gOmVFVtZn
xEXjX4pOh1mlPnF+31MVTBsDbI6V7wsxd9oGTNJwkBvwmfxv1ki50XtNW2aP/Pl1zF8gjBFeCjZb
3H3r4cEulZxlVpcOMuWRVF/5wpnpji7bjRcPmka8szoTWI8Mby7NkkGahWe3IbVH1foT+AS1AArp
l9jUje544U8cP1NrT46q4DTqKkd9I4W1o5f+PBSXNgkUplD19K3yQ9kqSStnNEhzA+Dxtmqfozpd
3gp80th2WLwoVOtS5bb+CrUO0NJIx9OXNarYa870EzrB4MrwocGwdNzhCOAPbafFEkzO0TcLzFp+
sleV5J5vefsNPmbJDx2LabfWf7ZR2CmfbIjBtZFnht1Vn/xXyJtHNowdfwqWmUwwYlLOQeVXZ0c8
Z0ywpcgrkZfdhf17TGSqAOggG7WFHftFOsT/yx5LJIZPLLdSLTrOLG05/062l8hD20gv+J7Ye1PV
FWZ/iLCgpyL3J+DJr3CIw/ty85C8lYkmEDFMlgaxT808B1Vs+pLlCfny3FJKsekTHBWUeVQ51LFX
p1uiDir6uBUrgDv+BVbDlMUp9sQI4+5gO7YFfg4883MESsjvPWo8LlHkZVEfMb+b97gHYXdKRkUq
UMFw1nO9oFVNMBjoNCh0FV/YNu3km21pR0cvda2n5grarYDc+9g5Wh9MHbRueeNq8EKMIqRpcaiG
90qwsMvAYkX8G6pfGkT3okH/uacHR59PNYEvzJo5iA+sgJyCAKmfSUN9VmApIoUXdGYaRL5CHIL9
XUgQHhiiIo0e7HwDHdyYa5QOVKD7HNw+rIt9rRXL0FLKIgiFDEMbn2Bl6dT376yUmfuXGFoGTgMu
nN/1HiBmxCouQjZ5USrIA+OuKGx8DSj6sHZoWSjE8yEVEBkFV/I+dVMInmzhOYQCHaF3l+ybRJw/
MAU50lVszm6Ba8Uk+0UqC71AxXKarNcOOqtuOxWwe6FyMoe9PcwIuom4ACtfXxdpe5nVOLdSXDih
G3PY+r6yRqqQufv+PJXBvMvvD6UVaGTesPQJASd0VPsTG+RuqM4GNVAbqrSOePYNy/WeI/DbQU1F
BlOW/NXEBnwtCSLdYUIXPE2HnPfG29azVxKKAAR1a/KD58WW4rjCmdA06wOd+dRFWh2qeLvD1lnC
1yFV+QMiDBeokdIJduPC3/niDriW/KNzALhDnvvX5ZE/Es6UooodnHxZo+ZBh9Fn8SJ0tvMw0ZSs
OOToYnBvfuigH2vYnj5pyJPSRy1KZYQ+LEgq3D5VRXmErlkCnn4CsPXELatxzJelc3YFZiBzZIAu
wSaJaBTpynxfeGgZ4YrLMr26VNFAry8OfZfbD90FQSWz/LU/jAeT81ixuotIkgDNbsvT/+BuNhJK
+jZlEBqW9yyp/YndfdLYNydXNnOtwedeJ4JD+tLFD3Y7RP46sqOLitWz8PePAnphprs23KkKGVHM
Bjw1E/zgB6aoVSgfDIgXWzJqmXT8WnHCfck57epIoDXMUVCNQZejsbdBD+hm+mn166tFZt6Pku+1
5TCGzWx83ENDhpUPrRm43LEgkWPq380kZEL5aU6IWMpaXCEEmphzfLOB9cXrywga0BgJGNcWlGDE
OcjNwHo+DVX0PXfZUQwNrXmjefHDFY5s7PqB86i33372TgOBIOwLyrH2ZWhdBI+H6J8QGtm7EF2T
cVm0UeMtOtzxIGGYqRp97wbo9FS/j0VkrAFO84+4bAtJK66XxN4E4K1W0IGeLRtc2c2hRdaWE7DV
Aso+wRjSam91jSh+jvcy1pOSXMLdgBTKcatIPOSitR1qfnwUaWWD6yt1pV2lefH8kw7z2QzSx1cM
zYPSuWypSfElIWpdz+bMzX1ZU9fbSzbaS4stGkqBGToAgQWcSfWHLDgjOpj7qkUhT4Iz/TSVBasA
G0Ju2kQ+g6z6ewPhYHB7EP1t88qPDdnDzKMjJ9AKxh27XeNQy/JXu0o0MpOvoXSiviz494QyVaES
0/J0hCFZ/zfM4FAW+4t0Xbr+NAEYyhCBMjVhlWJdEPPobVcrjoz2kZ1yFOXxlzjVHR8+ITSPEI6h
0iBUD9/1EKggZC77xBCcTlLPlXBBD5r/pB5cRF09+FGDnYpGsGCwldxUxCfyDwTkYUtFb6gHTAgw
PMwe51/OtjAaJZ2MU0zcrIpHS5kZLSgUfS/gj5R5QX12whEgeZ2omtaSVEdZlaO6FEyChqyr7fhq
QgH0Qm03KM7BsIOomrbOBDaGTZNBynV3BiP43S9VLqlw1hlz9cIoJMEfXBLesF2+9NULcTswXdBL
srLDh70WuP2KKoSuz/hCyn2CezR40CVY3KmVueE+WMdqQEwovfoWtqcIrc3EbZMO9v21+9bryl7R
+Fv5M2Br/5xJg6ZMyMMgIlY0dGfVh89rmz0Wlede7tFwHRfUuJUVhHem5kJcGbQQZz/BQ+i56DGO
YUbomvivX65NUSYEK1PcUa0O4Pq50k6LXMQTU97O5ss+5sYx83kC9j7agX4/WPAorvwd31hSFqXj
/XkHdlZa7TVrlwkuM5YMrREu2b9cX9NLJqJ7hJgSwqimOjd1Ko/YdMQPW7lhpVgAUBHHnyDoKXYU
14Bkd6MAxiXd1nth+Myb2fU9hiD556lpxX8KONw2kvpGjT1zFcZCe1ik3qTfDNPGbKXRxg4WbANP
SYF1C7YiXMeJzuR05vEMU2lGe7qxEUj2/g30m+HQd2h/FX3Rot4JZG7qto/1AFDsXvm6qbulOJOf
0RlF/CCL8gcYGhf6OKPdgVDidGFq8MiLvEG4ISsHIddS0cMBHtOzTBfexUqpqSB6eISE+6e5wJwM
YkZ4GYJh4KcdZIlkkk4g7sYrbruXSDtde5z2L67W5aEJY7JcjT4Psq2xzEi4LIr5EB3p3Xf/00Xr
1iIBPFImHiELeilbIp5KN4tzm4tmUZya2+EZBR778CuMXd3w8F2iPYEkNFKsN2hKulWUngThTXtR
EhLTu7waTdnXoEb6QhKha0imYEOtSd28lffN+aU2Wc9LrQe2HQRWkaU4EXYJf+q9E9k60jouezBA
pSi+OTTcP0mgwqEk+/ka/+JXxiozR9QcY+xUloXU83s5KsJfEWpZJYXWM9IzL8EUT7D372eNdg38
JOrP7zNnIgN0nFO8oip7rXkwNh9HPkW2VPyZKRnx1RBk8rNF1lBX6lDaBbVIDp496OM2sufvyWge
RBkzGzofD10koYdkSpuSGbkwVCzPWRP/VCML1bto6cub6uOiahlKiDScsMl6eEtEAO4O7u8Y0Vet
m3esxdfcHxmkyx9ztqJAL+iVyMxQvx5mCOOCA5csIc9AmN8BSdmif8OvMWEJO3DzObik1Slain+4
y0e/z78BIMqyhnqSrKs+qAQgnN+xHa4viWGUWKU0ZHUc53McxeQ0/zIwhX3kCdrHKwvs+3AqphOC
vvMCcxNAWydf34JOVln1HVDAaiFAX4u0+lediJMsoYwUA5OEN+bWRHBUeLxeJ9zSfogd383wW2AI
FPZi16Gg+rPrc6/cWFnz44XXcsp2nY9wiwUFot8W7RcI0/0aoZChc83XPHGd7uGM08OnO9FCPshT
vAZqYPFl7JILsJ6/FPXMr4WhmHZPzyRwJhPqcVihWP4b9PMxMM3GqTjBjv46yzpc+6dOqxg3z6FZ
eXeBxj5IsQStBeBhCen6kSCwt9yAQxKjXFBJfK4bcz9Lf5N65kiQqzblku/CBBSc2nLuqKHmORQZ
AcS3Xavtb+FNBswRwic9rCZtPVpOA1CP5QBbxqgsKWr6vRP3gwqpVf2807DFs+b/AHZFooxV1nsW
x65UhpaOD3V7pbgyNhW0se/0yXm/zm/bjzjv0rYjMhAOmn8jSM+lYVwp9NXpzlUjCrXK5n5bzdKH
A5KxkcQpuoPglxmk1cR93ixWeDMMRW3kS5vqHkM2pLl2w+XRey/ZEZJqaCJos9BypwcLiCnSuqTF
/i1nHa6Uc63Xwk1iMpvIApX7kZexQ7Dne6ay1X2eUUGy9hQKs/diG4eUJMdhqzXlrycKCsN3Cpew
BdYWNynI2hhWYTMmzWzhjZivW7PyZtmwkSfJ2PYjntS4aZYgqlHEAIJqxpN+O9RrY4q2mi/S1LMH
ENXP0l5S6PiGTSVQIhK4HZu5B98OARc6VYNWe/cd6umslAiYA46g/MqmyUTHunRQrYlhBfPxe1Dr
qlIUFBU90GtRbTNzkhYLV2kXBBKZcEqesYlPSrwpw3jHI0ksgcz99xfX/XsiVnYan2ISThPzYVP8
IndH90LD3n5AE5ENtZefCM92lVjgkV0QfDVmwaag4xl6+bL6vraoAVAKsHKee2tPlWTaFQlu6Fyn
iWaYtlyAu4EqiPNKkJicuvbYUqzFvOihmPYM6TuSEL34bYqekhIeTpk0CBu3tZFyd8PRNjoAjSRJ
IiC4VmwPOMXgUBawJ2M7QNJwP6pPGCBbVDbhIriaWgMjjfEa11kcLp8zn/voTlrvCCa9vV3rYG7T
hTzFEfLic3u3O7AmTKliIWQwVdCLQPQPiVckcwTqZ0dNk7djj2/LhYmYaQHVxRxGzHoUdJr9qYdT
nLxE50ips+C6j00OoZpCLcoVbBzMJCwDwrpq1z5JY8ylwLxZyeN1OYa4EoACdz07QQoV2bH3zc1U
9XQfWHNudxTPHsvg3jouzRBn81YP27L2vLn6ofwhRSbJOpVFy0EtzgOxUEj3T5hvcWCbFEwIAEWy
MJbzM1rA5uNl5qUJcvP3EVXSqtGpHBO5xXGqDf8TRb5aSj0XFTJoC/85FxH992HhI1VUmS3ouTCS
4CBXqpyZNRSvAUeippFk8kPJKVW6EEJtZu3s4chICF/+HEnNZ/p4H5eqoWuB0RPna/WqAyGCZe0s
QYdD6u3oN890t4Ra7bUhvV+z9I2I8+ZL/wY86nwoxzdvWraUfOeWaVyP4fCmZJsvvBG13mxQO8I6
A78PDZK3t+licPNUhRAHsszVuoQZ79Q31Zo52qRiwthaVwcx1vSYDYZwRZ4mXNig0Zdsck7JMYJq
Ei/blwjmXtdhSaYInqS1lscPHn5LQVfvqEjgpMAvEnML5tSm5PeOQhq97pHsoJmahsuZR2oDeDS+
n0g83Maj0KpEnkMnESQaoeJsD6kM1kGXcuPS4m4ZU/EW/PVg9o1PmD8M7yiBQawKD5UWT+4UMK/G
NvCOrv7MDHcJG85IaoHTyo6hN7r/+mlhk11bWSM3zK4FPmxT20NIUeqE4XW8dyAClk3v3ypg3cyP
j3Kn2xdtnLVWf4vxuv24CoB55U61nA4dvFBlqlHG620sYvmDLEjiTwnYsHFAnm0ah5773FhwHe7j
oUG/tQZXmLFaokVh54O/VJGWnf0kXGKcBmMyJZ9woUKuxiF6xz7pAOd2N9MizD7YBdeboMzIkRSN
A7UgKpcY74wmSrqnWkIhXoCuYIii9XlAP6GcPCk1f2CCohz9KTg3cXBrCEi0GDPxNp5AwWRssZWu
y1dDKprQon87Vdcf2dUaOl4BXmoqjyuyAmw92wI42DU0tzuoHMZVOvUA9puKKbAlFJisg8sJ/wAV
5ZDqTvcXxdIXDK+vq6qBZVhFtkp6nTr/YpH07uCBQjF+3AmM5w7kmyIbZsMhwmoJJ+b3djsmgXcg
7OsU43zBppej1wtw4HtuMVd7IfA2kBGUa8XYTo+wlZ6CdmmwjFi6TicOAHm9ISzNHam0lqspCLPn
MH/Z/257KJx8tx1o2xHMZMpvMMKLUUZWADSy1X2ncYYiMOvzOjhKnG4WniawR+/SrL6W/3H+ilJH
vZfg083war0F/Hcrfme6W4JxPM7IwuRQV13Y6IvDfj9UuoPvGgdVRwybX7okb57nbMkRIntTZbZh
XKg9XKxkShDt47W2cPNT/TdZDEf1i6GjtB2t/iiRQzrjaE8Af4hkGQXc7w25aAdof7wOxGPEm417
ebPwQzvadDypHNNrchnAWAbXAJncRKRMl0cx0vlmX51QzYDTkVOwG3IzYx6/nFUfIcuHKGn86S1V
RHud6Fq0bU4rb55v5eBInNJT3Y38lNXLvDEf2yCG4MH/kMKqGFoO2+BTnKhdxfOKWXc2mjmrceHF
FmwFJ5h8nDx1+fhEVNn3VY6McJR0Zh8xugPQle/3qZuTDJCOGRJz37XrESAW3jv6KwAbEp77gaVa
tmUYUMmBQT6EV5YZu9Dfs2yrxvhjOSAi203zy4hw/9fL0PY8+EyWxg+Y1IzwUw+7YblOglk2tUNe
qpFwaU46U8LewLmyIjVX/3AW1FJZ7HhZYBEEbEhdkcte6djVWXwQGPMrrCFQ4HF5LSfo1KfvYiug
nzuNRwOkAN+whXk+c26cgOtgFIXwGtxvRBi0STaKMC6I6NMiOS7WNGd3YJCKpUlhD0L31ru8M2A5
YYAyT5Dmxmw1TeuJrh8IZFjptsXq+NHAjGXwg3ec7Cgj4zSzRFa/BLDdZMaHjvHnQhokX24rvz1J
Jjgs9Kk3AHJzLnuLmgQlBIFRE/Gns1Ww60EWGKxAHo8qEdhrehG3l8ua30JG92dFWJyxxtGvDuJY
/4ugD/sjCuxlm7OmH+bt6FueE8L9zqJfEx5vgMssAtx6EVQJd3bO90C76mMdtp6SWOaI9jPK/Qkh
uacqwz3qFWlQ+/jbCPrf/bWouEfzbImDJvDLL+vqlgSkY4B0eYhOVUb7EWxHQabo9+TWLiWRK2CW
o1sO+MzQu60Igw9OAkz/nuM84RqB/wW397/UdoO/u02HibNMdC+Bk5kCDO40YUMmIuiomFQyLQ0v
iGh/af1Y8ilhlfYdtltTpS0CQsOeyPIIxOOBS8cpxx+7q0LClEVYG7dHpCv4utp0c4ENe2oNK529
Dezflp7a2tpYXkd6q0H9anA1SDmHUzMMdYqCF/P54Spf8rR8hpP/sPWSSJKdr8lUPZ0PM56N6lJ4
VaQqbMuA+tD5xz/A7aM2M1ATu+TUrL9TZS//zLV3l3+haOlHlIMhasQxGR4GQY06JhPB/xk97W89
Lv8iQAmwgG9RGIu9e5OyNiqN/v9WdSGbKewZ7k1YGNO4KnGcT0O41BVSOmHBqplDGiNuEmU3ZXiT
Zopdre8WKiK9sKEj/c5Ls18BZVPNs911XbZOQbWCo2u3kyYHtBIl7XgGVhODHQBpw6Lcy3jGhHGC
pC7JYrtse2z8rFuMnsGikGYKIzZGJ06J/UvwbgYe5cVL75Vo23rRISAcb26K5DDpNi6j4tTN4oGP
Lry1V1Tr2bpWoRmR2ejUneWqrIHl12yw6t3JKoPdh9AdFB0hZxwTUe+xlQTM94PUkDHrO2jqo5Dm
y2pnNDI5Ee1SWjgm8j+sK0St4iE9UlDA2WGpAfoT3uJNzA858xIR1Sw3gO5XAIZ74lsUQa7iYQFy
7sliA7wS91zm7ZF7mZB3E71+h44uUHNA20V85ccV2CaEaxCpkaC00rmIhorfF72ACPv9CQb4DFIY
N4xErf0L/WJqIiccpCLK9OqVScGC60G4HTeGX8uJRok8kGlHWGsOmwYRXvadhd9P5+iCI3fzrhfI
kgwZzNLrrIJL8BcJTW34Ne7VfnxzQRhpimIKYfA4hq5/C2z5tVrBq/60j2oKpzLxnmfSo/3ajtzb
2uZvem39scQtCX+ueOh5WW0X00wX9Ct0li599c3FjyG+SI40soK5sw+TF/5ie7dUwVYbJ9uVJIny
P9l8szQGfPuJRAowOm5IvWCDGriz2hIl9jgCjNgHPGciE0ftNCofSadGZkUUHPqAYdvw7+I/g2PZ
D3unTU0ef5Q0LD8WM12F1gW70fT/bz8Ia5BJuBUz8SrUeeaX3lHZvkH5EkUcP1gLCyBj1kn+XrKZ
x3Px7+q13FYXe2cWA/N8MgTtladAw7DzR5mWmfDx2ytz1vgks+pKqzoeoy/HyO5Y8r70HLBurg1f
iN+zXtv/3bM8NudW93mNCSCSgRgs6Q/V8dpCS5Yq7q0445KesEOmhnKnqayGt303uftRbbf2/9uI
KVKA/fN7Bxsct/fc3AnFyFTz9GvD+jt+F4Jngi6f8v1mjfytLSgSsZtXZC6Iu6GHJb7OcHwHjjB4
fjenfv+/ofoc9ftIMAH/lg2qoyASm2m5ie8zcvE+gwM/boAyfAPlBss9eVR1xdfZ6+J51xuyyZFH
PcE9wM/CrWoA3v6bmpAqkeuJ86FfFBltB4gduSaCnTLS6HD5qjKFeCRTwclw0CZhrHxfAGWxO+V8
82a1JQVmoBYJWk8WGquN66lOjSnBmPSJ5q+emNHJ7S29bRe5t1qBYP6CgQBJIJ6td1fFeKI4FbwX
9l8G77SiXK34SJPoslJA3fgXVyttv6oRQinSQhVM+G/uggwo+rckaQxC21r6SWnrZh9LiW9yMdx5
KUCElaPyzwfWYDUq0qx2V0zUoBCV53dE57pZf2FthzPP+KPi3cCoGT97mKyLtZdQH6VFxHVD0snX
uLg3p4wVyYHS7ADVAV8hFokYKDRr0GqD/gKARlqpC8r9xVcqe1P7cReo7KrPRZT+/an+9KxoGO0S
cq8D+gOBntZ0L0hNuizSjf9MmzbiCdWZLmcqL2YegsbtbtZ2Y/4AUXp0wzdnRIkkprJDsJb7DTNZ
j956gnvuLeFTQLiGUHbK0J5i9hMdBl83hbBT8Waj4BZMR+AI2/4uLgWQ6KH6kNmfK8KnVKcSDbmA
kUUwEDEqoEyVy6OfsqpBN8wA+DsDI8F2OUlj6IolpS3yBk2+fyKY4D9aBjpxdOAH7LUqswkennR3
qDgvSKyZHPeJE1L6rip9oiLGu5QlDFeDdxFXdsqMuSWXZYeNtC4Ws+i/jjRf426Ipxkqq8PMQzqA
XmyL0e/tcxgUJRAFiNLxHRn5+AH1wrTeX8meAZouVrvSGPULsv2I7Mz2mG+wqk01BkqZVQo+uVK4
LviW3tTIu8SY/pAUnGL88SYT0SZPbZRzIKciFstfNVqpFFXHXnMuyegfL2wX6WW1oBJNjWg/N5QE
Ee/heOIuj7lGHbn+2INLBs5dvRz3cTktcd7ePH/IwMWPEBJjJe0L4eFrva+Qtq6qKrXr2aPNBXpB
+TG+KFhfNo2DXQOXVfpBpYfGUvoVx6HueMbHPrqRHf02UQZoVKNjL88TTBCs2yP8IE37nv/IIutQ
sq0Z14ccDYBWBVCSds9sGflo0yP34pGI1i6LwRg96iE3338UaIhbcm6LR5oFL1qSxIA8oFkPza7u
t+Gkw5FjdfnLMAXSNzk5rYKlcdxL72FsqmPGJULbdfqUt7eQ3AmmsNxA7URRf2CpSyDMNwW/AFPL
48ps5YXch5A5RVmBXxWEm3Yg/F368/kUM9QPwvhBO6SkdUPDNB64Bids8KAg9oKHs7Y2Si2b0/dc
BurDrmBZGJrXSCdX3VWl5zH7h0++2iJKzws0T5iCG2NPPzmoZ2ZBq5ivlUJwS4w1Zf1IGHmD8nX5
dmcWQeHnDeBKGs0UCAPMuTVisLnjBvscWZ1BkPH9IuDg/FcNnZr7l7HiSUZTT6rIh9dRIRevoTRi
/ZkbKIcUgVOTzOswg1ki0UiqwvyyKTJSD20IS/yWq3oHzvgslkoJMRckyu1mbYP/BzriNd15FDGR
oSt4Dfeg9AAVfUwXxY4FAmCT8lTUXNc+dIcYkLP/RxjwxOZD/bbUvhrA90UaKFIOChbvzxp7SOGj
T7+9ODuYY+56hNpmxLf7EXw3exk8ieX7sZL+y3uWux0O8rGt0YhjP4T3VrM+wvMsgyTET4LP6VHd
Tjx5/xvexBLV5Be+lppZkZQ9ts1Emhk+BNmUuks8ezkptcZa9wR3sKOESoRGv2GTL7kra6Su002N
ZMDuCUMgohKMP62h8ZmZwx5s4165XzzppBcJg39eGsYK5G3ZkqqrsaCNqdWjqoCrHuMxJTN0OQPy
4bfbtiMdcz52LKX3OZrrABoAuR2EnvKyUyWrWTvwYTZOz6H8Vg9u/kpswWh1Ko7B9TZ4huLMvltT
jncbY1ik9nkbqZAI1hhJ+Wzj0/Bqo3XpgUKJx47LCYpO0YAkXyw327+y11K9/pcsQlu9InFa3wqk
mgOmB3Eadrhgk93knyANdn8OGlEI5xZeB15+VF7CMrhY1AaULyhXWMCVWDjomnxdj3WZmBmJbx4b
wr2hgNZ7fUWx5aaTpzvmNAT7td3MouK7XiS0TROepAwQ0h3g85AfVOEGKBpbkgJxusvkGXKcdd6G
/720s9hrfQbgxjNY9IOtgih2lSZWuMERX2+KXkLvUuDXCLI+cOXBNBnLNupXo2MgugyRCWHEuQPX
sik99pA1xbCtt2XN+eEgCjfvaYtaLyduS6QWqJSiSKUFWSrewukJWKks8erODyvXBn3iapdAgcmR
+N2XWVseodyE6IFSwX1iklqO552lezFAyplLp0BALLjmJ9INq4WEQEGs/HgZgU+u7P2WpdqGMy0Y
cSD/IFa7XVc1D+wXQBd8JiibA5GEA9bcIRQToKVtyz9g0mXv0uKkLr90Qj//Tkv7hoUbAamjEkbQ
n/CRWLplPGHssjsWq5R3LtBrTJ5t6i1Q7iThTjsUbjz+YTW7+VagNxFI7lVT2u7HGDs+rDQL9HAv
mp/mHI3rtQ8VMwWJ9uEoorYy+8huuaQjU8l/qCF2HtMGpdI3KH8zlD4zMW/JJggtHr+4/q6x21Mm
61P+S6d75AQShTS/ctqKTUa60/yZou4srXKBgu2skEpeFUE01cuiTvcCOFHr5CSG9knyxR8BWnu/
a5JO7I32yb/Pia939jepODZFoQoPFXqAr9AP3IbWhiSUkMvlUhu57ukMuJYYw+VEz0KSCHwdFFQm
ZpU2+P4my72wVvsO0WxDNK0fEY64s30o30eFTfA350laOWi8eYrByrB6KfYyZq5zCARbz/uQocQw
XeXkJzSofaKI6rrMlcZpMrAsvgbihRP5O5MhIylagPyGWuXJ3p74jc3cGrNn4jnMYfXXyLskaf3D
G5rsFs1sp41DqBdfollHdF7jIvTPeyjNI+dy9NIRTO0FLUdPV+xmRcPnru2XEKYCJPdRF5/5hpzG
6Y+3bTdx/y62gq+Uiov//mGQhUdvV/wzc4XLA+q6IK/WPGLY/+FYEAt99g/itp4OC4JqCXiiouF/
slv5xrsbgYiFzY6zjLcPg4nbx2g4/dQxOnyDUOM8DVc3MaAheYWwrFK3hW213aZlVsEUWxOE74Qy
kTAo98hJXjmiqcwJ4KYRYgKrqHn+fjRhLKUif0mlBv16Rg+6riJBRI/uJWizeMvyX2fMBz1lNQpJ
9W1yx5Ra5pRAQEnM9mrhoj78CP4ixqb/shb3RkgoDKm9J7ekdesGZloQgKlEM/ybnttABFDLLcPm
geqPw8NStHwTRZex/kHB0eb8o6wFxkaFlh2V8Xkbf81kwrXi9AHFuYbORrAb1j1onJ3uFgkE0MN5
Q+S3ZzvxIlcByKOOLjSjH2kW04qM6buLWrHtF7OaPBEuCvNmjYyJl4QtSpAcwFtacuutfLgDlngg
u/bPVE02VNsBsG0ccwjcmtKFK0HfH4GKib/fqrOd4Xv/Sh2QYqfazOKKKmdeThqa8HFztOJyig8v
DhmjbiSCNZsL6R9EMp/ceQSLcy7N1lXR13dPwDGDuexoaKPSjLy+eOUeQOEPPd7qxw4m6s8O9/x+
dI70oiky1AR3rKuMljr7yGVuG2HHCO61T4MXPDkl3BimJO+TXiFI5ti5jOowGp7sN2w78UI08MRN
WCnwg0rWIyAPFKcuM7TogtcTfJQhibAnJU5QXeJeaMIGdzAvKPXJQ7NmoTICwT9JPyHPGe0klzD1
G/jnECEoVUTTDmtvCqwIf7Q+vfGxqn295HTh0DCkMqEo+YyfuewOfvJRLZNG9gBvxv2mloXgNdy2
ewLr3cY3yyYU8fjlCLWWKdDMaBGv5tbTu5688p8NuoD97nnMLfJ04TTLswBfBZHVoO/Gq9MPd9b4
2rH8MM30f4WVcH3376K4/fuTSmSuu+vpcrQdVYNd4sNE+g2nY9W9oVDbMYLHMuik2IrLPqNLez1y
zcbXvcHv8bUbLkcmmw14Ks650ak0t3+KrRr4/ElinU+ixL1N8lz3dLPhMnKT5glwrunoT9G/riji
yXpxoVqxWs0owLC0Yiz27lU4vgY6Ev60EN+JU+G7YIsUDjuLnHCUwqOvcHYON6y4+IHQHl/v0eZK
NH4OgzpqJ9O+TDfN2Tt9muOGgUkYyEy9Ua18oPf3VaIqNTn0UEnPs/e4ysnnLtQy3lWN3XPVmDlP
VGTykSyaYxTQ11thq2JAWNcN0exIk6WuHzQLLKmnvWezb4rajVucyIlhMjvKN/WDniDHa65duuk7
3sBYlEgYJUtO8M4Zh1izqyXK6mWz34j3nZUahUTzoayuagkGY6N6xHAM2GsbMWLjAVNTksJZGaLP
uwn91hqSrRVu+uQgGN2YVhFYOFfm25cjQa+nD5vPPeO1Fe6C8JipwsKLgaWSWqY/sODeVrOTTUBq
NTSFryOrmv3zPuQ8yelhXQmP+LfJsHJ1M34JayuQGOBcqOf7yBihsF86iz9PFI43hi1ZezFcZJR3
hZCxz68R0QzRBTyf1shGyYjfxhoyHvrOKctS7lGfENC1fFf897+gvt/ssPyL2prw/tXHT1abwkMQ
Ldz04CWnWSQsOCchSamwmQHuaB5V5nMqdx9oaso0+a3wtNFWP2d1RF+CqF87ImErRkDErSFsiuiO
U2uYfcT2b87+CQ3xBlScQjeNzFl4OpDbEnDIrvXaAjulivQWpD5Vt0RNH/rUXW2EFX4bXlTUXD2e
PXD4MZeIl8i1KdgoF1vZcjyviJmKTvPZejStNYG+5rB3iJOkptugxPsLfzvTTa/gmmW3DIMxrGgY
y/Po3WToqjzfCRkIWpc5O45w5smoT/grG2sTpdQ45lb7TNv6/G7G6sWi7qwRYxYUtEDRnHslDVr/
/fj75BulIEyJcOl6Xo0G/8974jDHWmHCB6qBCViFDM0kzarTawu0YXqxYLcVGT9GLm6eanmKgmgJ
ShIoVn5VXaH+IUJusu2DAaAau39hsrfhsV/04QyC6WuRPBnKUofD4zmeBC/qRDIfmBXLeujCHBDX
m4dyBK5A3OEcdxGTauikpaCS/Vr+/4a2lmxSFVtiQKmjvPkK8fMNiny4oxBBgENaBhRbZcw/VWgA
Y36P5tPMa2FJLHMesEjEIQyg/2P3E+61dgnf371PY+TMvw1+LgG0cFkElL2C8//c/lYgWP3zrDzD
JXm+M61OBLsM41GTbTkDOvk+VdTFQ7y37F+8zkjpaeYQJi6DeY/1LFvJXJBfx/Oy3qvrJXDFrBEe
D3z4GNl3HYfZRZp1vNkdsT2/KxcSCRYywIBAwOtrScQNyDbsqXKWq+32W8M/JoKD2hiZHambvNcM
ijXnIj29z1z6WG9NA030yPMyj6Xu2xaWDptkWES602ivPNUfx+tPJKJEhvET1BAJxG7nfhoiO3NF
BP7MFglM7FpJxEkZgiJTVU+fSlxLIcYToadUmiLw+P5Jz3I9geZ6Fjryc2/AYYnwcrQKPMxSv0uL
ktT2uqhetL7Mn2SIiEs2WTIczXwmEBtI/QxGzlxh7TmoLqCFZ/+y1187w+uHza5V1tj3sFR01srQ
w3l0cHf6dK5BheHN6lbX/Q1/rmRBUduztADVy4KRVDLGhqHTYwxNL63tlgtdIwZCwZmDo2ZRj9Rv
7kWFIaE8lFSecIWjMLGDk1H0F5mFz7gOdyP8V2xneK0j5SJUfw8Gn/++q6k8tMUhPYeLGZCL3x5M
CRMI5Knyb/AcB64J3OdjFM+bOVbOJa9WoqOyWzsAA33gZvgoer/K6FhxX6eVuNNiQUCRpTUArf9u
Jv6L0wFalVT8OL9cCNqkM2iyHGrJV+KRl3S9BNfIKkcZgVrnvUFoBRC+cqvEJe010S0Su8eRRgkc
6K76ZUqVJKtEV1EapeMPv4hBClLiVprDXtk5CvjQURyl2zEpa7PGhqMAZNwblIX+nSSSfzst7oR3
1Q6gxGIjuJESazXDP+Wr9W9uo0BY2GqLH5n2K+w5ZmRzN0njm1OVMfuvC+r228Xhl2FFiimwawUa
O1AWdlOucrpVS7B2TO9+wiZev2CeyatECEKH+M6oMGn6asOE/LOsvHTVdya1XtJu2jhunJ0QYiEP
MYmb6Ma3SZlIJFaUBE4SKObSnu00Zxrg5SOCxjHKf1os3rBdAhAs0jtyslN9gezkTZcUIMzE5hFF
gc7LWu8wzrFnY/BwHdTY6/q65BbntOhEax/z59cBR3xcfGvrb0vgEHR5udAT+YgmdhJDlWqORnZ6
v6G6DGfSlyw3YlocpCAvw23pv8M4ZEFlk9yMm37xg3s4UGVrs45hDC8HdTHcZoyxEKx3XwxbAP29
XLrUlpbKuJhuWVlEaP9FiODk5C34AZwfCL4EhKwu5iHDR+el8BZycg51nEg18JVp9fELqWxdeG4x
aNR/o6vnFRgrKQJvW6QG76O24nJBOoipFvrvbbDO/vS/YrGYmY8kMDLoZ0A7XPtVW7nqKRgrooM1
iFwZY1q+FXUwnKdQ36bkxt7z3RrWkxiyfCmCZlj2U2Z4AZ8KXJcUpxw2ZWFN37PDmRP9y/4LBksT
WHa4GGcZw30oG3MCnab8MIxk0VCEAAgRuqtLrtTySTbcRcYBVxSkbmp8vKI4Z7pgitk6+h9JQjxD
SnvutNyZG3GB/6fWduIkuMrWJRHAOb/pp9b95eAIt1jxR3dl682TZ9Q/+MK7m+sw3vQMxwl1fFlN
n8C97EfwZe9AIdSctzL6U1TAbHMXf83/YXihA1MdlMwpz41bWmc2Hahjm1AAbgZYQHYtzIPUZm2I
SI1AxTnwbOY2lxt3eVpH1UVq/CoJdfddtfc7kW3Y1/IYiuK40LmedA4pxsCrTwiNnPqiM9bnTBa+
Hupvt/pqucfJnf0hw0N2Z7wsuVzJY5j0
`protect end_protected
