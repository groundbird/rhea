`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XgIyvdpLvOY3eDF7hR+cj6GG+K2D61nzQWIexteu04e4WqfcO3Uih74KKdALdW0jeCkHR7KfELlU
0uVsvf6nKA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dw4ChLNnQrku7JRvOl40SK2bfzvHDwuqOdM1otoWchbEHA8eCV8ssbK+lt3fWgOqG8SAX74xsuCX
gN9/o1fEd+pklZgbM0tkH7BdxLILtHOxvD9ZtqfG6/xLioNXpALo9eDc4fbVqhiy4nr1uJ0bdHHJ
xeMYzUR6HGY6fLMqbOE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RnETH9tFxraSSlCGGWscyaQU5Tlwq6f//X6FTPGM/d/aKNZThtLhoxoPU/WSfP0Aj5PcmDBVRT6r
cT3xUiQdOvRCjbwm8iu+TH+ZQ/KHkG+/7G7sHZCBsAROgU+b1CqLUj2S3bHBaeqpvXeIH9bfM968
eiGT6xhV2/yei63C7vUzem0KnEAkUpUR8S3dUV/J8vGUVeg0UQXXGyLdUFYtyBn1IM9krt/Wu69V
qGQLNwHH+bVk03ypse3WFHXXfjfIH3rdE5gPJaMcC36r3orsoaWfm9wuDu4hfiMqWAlAxQsPTBxq
Z9eATg8ws91oCFr5Anye/2rY2szhakdOxPMktQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qHUjpMpagkQwbqjk97T172TtOeWCNbNN5mfCu3nXOS5tfPDQW7sJyOBCHhwHpnitlt3IQ7z53/zx
Z+Qctc0gKb11gqbjrQYHgE14JIMh5NhBD3A3efEXTBrswl7Ar/v0dLaTh68nXBFojTz7NcUwQuJ2
lCbQj/nFdHBj1ttiHDw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mU8/+nzM4Ajd+TaX3YdtjKCWp3nLePYGFeE5nFNUxQvWqEWMiYbz+VaA+H2SSlTBoBkpiMp0Yu0k
6xiC2O3EYoTE64hRaGgLjuoOX4Wq98Py79QQQiLvCR6h8Eutl2hk/0vqxY+SQDJdoZPmv6C4eN6z
MD9rGIHiomWXY5L3dwVcSjFR13yD9yNBdHRkVJBs5BvJQrq1HEfsHiATwSFLtUdYrkQ2mgeMsE3B
CsP+S+qhEAbKz5gzsF7x7TshtIoUXgkQmbiq23KKQNneu1r/rqZec1e+SQqWCICVPcTi/zE+7eQT
6aAqt9kMrQZNxiSsBlxInTprlAvqCAgsp1MyQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8016)
`protect data_block
D9XTQQnu2hK4FxtP0K/v6QeWw2iCc+YXiuorkd2OgExUobUQNpnmNZHfvwzF23ij1a7TqzLX6whk
ps0G2defhQKznJS91rd+zCab0KmBITeolWumMMNXGJJFoKxi9zfGWsgrNyxBbgDUdpR8sG1jdWe7
ly/LtWRxDWetmC0RO5qaH62jlf3sQ3GmlcLboFY3AOvBc+0/vxR6AOHYHO5KHjTjjnd9Gmu6iX2c
3E4dOwa0AJBnBNFZKvzqcaQ2oqTYqm/xssCPL6qVGn0oX+d2ovRLe9Qo2AV20FruojKkGYkBFAuy
KDaZZjEAKMASrj5NoF4BfM0O4Adb3eLPc/hP8ZdxH1yNNal6LuJRIJoseEsMl7eXfW4kP31jrXWJ
RsDEYnMvUHEF3BPaeX6/HL7tQ+XpgH/pTVLya361xCQNP25xTE+5iQA9O1Jym36xb7+nqG22vqTd
ZpTrjy6dyfr7TO1M1UamQ3e78b26WXAZFHkcqoqfc0Bm5Gu6Hvs/ZG6W9uPiPdIarZE3O/oVI9Ox
RgjTET5e5wNkWKoAQbDdCOifc7bWzJVCgUfex28NAUpg+Fy8HWQJTKJvwc6RvoovIHXopwSOTpR3
WnINsyMItgx7Bcor7Sv96QE4RaJYUPsB7XwxNaGNMy3zyKM+dK/ufmSFW+G4jfxM7uaDwi3xVpC1
mvnm9un4C34CY47JHZbI45XbTJBP/a7Ykx6htH6yJgqnHqK4n36SGFR41E+vDIceZFq5gTWZXSbU
CHg8ENbvg65S7V3QaQBgHg7gN3kD83ng9VRQgUSlf6PCWck+PpbuZE9peQ6mYCEalFq0qod9H7GK
tFBiYFqVCQCxYXqTiS5nIMKOkhojixY8A0Nb9Xj38dBXftLSsFGxrN21ZeFPWD4nPM5mIv2UInEO
7K2ekXHL21/jSLSHMC/h4suRVnmMrfgBFOx9leWZKmIn/35Ut/L2VTflJFuCDzpIvjqIlDbKXO2z
XNR58Y0sms8M96wd846rdwwOYHZz2/nMRzrgWPFG8hy5Ki63vFmGpPnNK/B7yaBAY/Eiqd1SmO3/
gEuIuEMImdRgi5Vh5EV+xPcPKaDVyMp2SiBEyF9GUkJcVBh7SYJZjmCVX9vnNOMz2rKUtkjahcvr
4NImYdl1kynaGPFgKhLyCVQ/dt7ZtB0CQI+bC+qmhYkiggzWDTVkCk/Et6cGuVx6XHKtC6YXeMUR
AQg0k/i5Vw+bfRNKfPrj/jCKfIE1brns/nVPxIN5R5oMwV0nx+YeiQxdGuJcnlEatfEHJfHgXprK
pstoMmzTZqBX8w2jNDRjUC95uUZ56lJiNE9HbfyYhJ3iuJyTHb0TvrzGefyCcIs3nWEz+RzWMYph
bdTNigHOj0oa2f27Gix26GpjU1E8VhcPgYlkDsYDsw7/vOfbc9BY3FlrsRI/V1ukern2kNTP5zfL
tZaAmrwz4HxRB8vxYDbvaaJM4cgyI1RFdbf1tC58YhJR1NlqXmhR0rxBA6bxsTrJuLKaRXgARZ2C
5+AN5XxS9DMf42FjmuUD4sZNG6REjMZMBewd+a89aMZRcaK1IeTxKbZZ4jS7fW42b/UN6MsAl2MW
sedxHQMlGjVQpe8YLaOz/GcbUfjikRGj0+3TC0E/W+mQCbk4wyZQXTyw0pPWlPbkuY09Hr2NDbhO
oxupIT0zIAolrtYx+AN6lUAqVX+rG/QukS5tZ88F9aAoEjDAhAnXmtw/pHf6Vh7i27B9UkQRnOQL
8ZugCQ2nv0RxBiYvELd5Ih18NpzBEGyMXh19vLFLb4ma6jR/YOu6FPRI+xHnjVftNye2H86WGAPA
qW2PDspwfniaAOzPY15cihft5rFNbW8x+aVaMEFj0PG3qcimOxMz8n1GRekojB+KAk/Gzlbe6ky7
nGqD7V9Ma4PQ8qt7pBHuDF/Ukt/zQivo9uHtpbMBkHf81pYg5i6ZJiLuxfCNw/YvtlA03VgwPrFc
n4fKdA+6MDqoA9GIjR1Dpm7GDpg2it2L3JAF70QrqeVLZCbDXriGChhQAw5WtKwn7/ALuf6YD0v7
+JatZB0TsPD+TQBsbf0HvCNz0qRnI3hwd2hK8PGg4auIJWkkN0aEM+oUNg2g9LQLxTEkpnm1k5j5
oURU3xSX4egiWhLDs28E6vpicxBRYtxH7o2Te4ZczfbQOyiiDhxrq7zXkB5Si7T6uGSzi2CkDd/1
SO7D/vXR8Sa6jnSzgFTF/XEyI/nTsBaLy7AGs1KUgDTSmcZiMuX3lsstimbZUD/tKAH1QeiU5mp/
jySO72Q3PQJ4NqZHX+yspBMeYWnPUSEwkAL6Wg1zE+SqFPMxefqgOEoIO+KonmAF2j897kcpqhnT
y+PjAbDEJg9AX0ejMGG27xAgdbe9sJH7y2pyqzD/uVvZds/5fcjyf0UUxy2RS9G3jqS0VNnzy+Lv
WpC9ZTeyyIEok/eT4/uHnYxOMMEilPV9SMHOqxRyMlu94b4yeiLNcXuIFeBC5UOftawP7QWYuCgA
hBHoKg2YcN60wS2b+Prbmn4sapUdYquX1SthxToUkRUWAZ/QE6czE1U1Aor5AKyiSsxlZjMj+sQG
Gek4IapeMrRuavNjmL7vvk9ZpOa6RHkix2vUF2f/nMcGXZSdejr34Uozh3iQe7EW9nWIDmwguZw0
TYClhSSSFtEVtHfrU4xWQyGdfuo2s6ePBrHtZdXiOZA4MYBkcxo/eaxzVVO4Xm+UXEFUBXi8rxJl
/bCkQlAU3mNBsJqUNF5wryAl38xME0P795aX1pwLFx7y7vKJsZSpjJ+e+qw6IyiLbv9atL+kE8bC
GJov17nLCJveRGDSRRljVnZ/PXbhedwDSULXqLEefUqncB0Cet29kjstrDBDpSSGjYj2mIwMy1tf
kTkhjWf2XGjtPJ0VEarlNzhMwhNFaBhMZ/rc1Uo2rXXq3MBLZtqsM8Z9OtjWKgEXLuUI+Eg+5lPe
BxQSYsdv2lHLwF9w7mHTleHUyM+hiZUtnkSgKhhfsoSMfDlc3RiU+YwchSO4s6kwScuWfWBxlqaT
zz8BD6cNvyiUB5lpC6rZ9bp8A5Vlasnbxe+m2DN2xhERw5bQg4sgKas0RtzwbEFrG0MvDxXxgme7
iUF+ZSFaJeoCD325OLiEG6pFFWSM1XnzMcf4hc1mPC4WRlrmQYmTT0rFRW94+Ah/tIUgGtbBj8hh
GOzy4N22NLJyucJ6g9ho0yJ6B4b8qI6AGHGGtK4gV0CtTFnbKeTj+GQDgK75gFXDuvOaG1oVhYo6
lqbQazStUHlHzOuEdcjF3Z+0W4UVfVnepoujn0+QSvkJR/ulSpuGrF0CC+nTrEdhHkLzdU2IZnWg
R928IJplulAc/6HXOirjI/ZmF/6uWxTZC3jVs9esgmiNbBj+memE84r9h7/xTwJ2hmq3AM7L5V09
S8ZJsZl7nyqBe8AwiNGR7wL+p4ktoTkjkha6JPBNVjS97WTDJ29FxuV4wW9ds/WOBD86rE7sm/jp
vn9EEEDfpa+UWUguKmDjss3DAAuac5v+dq96CQVrYWL300RzYOn0UtZpUSC64KMQK0yzq5RGiSOB
1au1mh0vCwC7+G9l5e3qtcdUXSGpLot5odvkI3hGVnD0H1ZOaRCLgMPNRr1VVal2wcCLsFfC7iW8
JvEESkqB41I16/5qml8MDPG0P40iUK9ElFGbQEDpJjzIcxZ+EeqZB9aZI6/oF/lqyUsNVBtKZ3QR
kUsSXvY0Fuvv5nRZP5Sq4a0Qfm2eRGjnxZD/IpUJMM6vQBDKQhuLwg2PQWM6s9xWUWaXgnOFucpO
U0rNZFclFN2M94sleSb0iKP53NJsGrAQS2zeNI3L1o86BbaK+WM5J+s139Pb5yGfLYeWhCgW2lRo
a4/AbFGAZrry4kZflZHlPb9xUE/gLz90VzWRvJa1dGT7WDj9wOF12LBfUOI1un2d/SoRU6Ps60f/
6/4PLQ2No0/8vUf7zGQnc6roEnRa0Rx3IvkLPdzEbgQEMGPNSB6IkoMh4RU7G+SlZ2zjTpRaLtxy
JztJ5Mw4HZK2b+cIsOTbAWRzZOfgzO+ExyY7eSfjLk2QpEwRXV102xRQCW3R+CTbrE82entGrPnC
mTy0F/S8kH2YeGZefLXUAvRFVaIZpTlulUsdMtPc3q1JZcBBlGYiZPR2/fKtElur8FsV0+DM/jRm
hdzjsgLEHkVmp8s0+w/tfljYXH1iPk88yPmDsiTf8kTxvDPGliEQ+ho8YjJwPCbDv8KfoL5FSytj
fQwS+/pJ/nPgVvrW5HVsWDtzjlALiDekRpJ1BVadmlAoHI88fObXJY3YlARzddMnkXCYrTadmj+e
rXfdcY2iMRd6nOxyLBkpbxLPb1qjEqpkkeMk4Ua/uGm1i/gPVojaP/LkDa76cZnYS/U5j0KG2dL6
bq1ZrHT5jJvOcGHHatXMJu2PPDASYxmPf3IUV7eXXK9YssolrkIhO4M17Cv3ZIIem5c3uDhaXxSU
29NeriokM1HTHtziviUEShXjpP/0rr+jHxsvegRp/hdXEiHpHbT5GVp1g+rk6MjzzbKuDBm6T5Oa
2DxrDcg6Z0TTMoT7AU5hiay7DKuQIOCSyxjTjDIOOUS7ZFTqDIkhgEWA1dektigImLq5Ffa0fY28
PIZhca+Ya3AtGRc5HG4SgP46NhS4+PRiUT9S2IiVy8lS19gRtHWAYl+FAU2k3wG3bXKzYDRn5RvP
akLnjzf6TF0FZ+caksp2QJJ9KrdFWzc7z7CZfEkyfBQHWCM2JpJnkvmDsTjvqCqjhRNhSoLo3xS5
pmwspT/RiY357eQcsjGhP9kTdOSrfhum7aDtdsXpWlzn96pZmSyAgEn/6BJFa5j8KfEcA1a/iq/+
kg1f0t1v96Y8jGUywaaToC6NjyAsjnJF/HQjOmJrFCgTZs/BKFsrya4XU/t1JqxDUj+CehaROIRz
Dgqvg2Yhvn/L8ZfYfgTo8K/0xctzdsxpDMLuxIZWvpJyqo65HiTR8Uub1LTY+2HP9iDWUL+42lPn
HZm94lP4r7QMMTU9vHUerA43h1YwlfL6ZPAtJWcV96idGlrUEDbwzuBztUf6rGbFr/syvyMReuc6
uMEehITL0lCCUID6Dp5CHQd8XqPc4FOOqRCek8b1EwSTHpq1F4/A3bnNJjRiQ2Vf89xlMBtmFBEe
DtcziupDUXFEH2adFdFpazyvRc9f9sHbilHr11ZtvUiyX/fFOB1vuk+zNTUTv7WNFcVxsxZgedC1
mr4AyPgE8f8JdLGf8eFMh/uRR+Cc7hnPuZQyJv9/njHPcPHpUHVOpCnd1+erZT9OfKPp1lBn+kvg
wMxOQOWofdP/dJELps+uMBreyq4IJpuF1i1/hRJVIITAgwn7Dl5HsVKpZ+iKtdv9MJqNRf0WNeHD
k5+ewhaNAm2KmOnTdCL/tjqlS41WTz+mTJ6l+PrMbCqjqfP7Rlqd6HxS6y26zNmqy2hlUelvK0Iq
Ll4BaxgapuKVaFoDzVFo0Jx01it6DivynJ1mUsr/4SM3RRSeq2qyFYKMYA+7yzsLDpXA+Suy/MsY
XnfD/YPFRytnM/AyBDYmqGvuKQ+4aBPVzQWLPxLgzl7rYT6R4Ed8kDiHHtgdt+OqClwJn8O4zbla
+KfFY+sg9gTyaT7MYTKFzv3dYodohgIcFW0LxM0GjOTg2LotJu8rRuYQuy9jvofL44BU4qkIS7iA
H1Xru3GcjEZVolacjLKhMhshLe9c5g6W+3ZQLhEBR7YfKK7ljLyUsSabjzNuXNLPT2MpuKHjer0P
eJdGutFRTly7tzWGykamQq05KSXefcyr6Afr3yOnXo6Nx6GDIArMtQywsenwhB6+QyvC7waePA6l
H4uMLzO1JMWL61sgudgC0vjAtb9q0d1OV3pB4YgVMlPTLkDNbOIbyw/DgI6U03vY68Esk8Dhm5XH
GmyBPdRrvfr2UEv5W8AedMl95Md85L6nUjv44kNNvVh4jaMb062yIAt2MebcTseJyN3/k8ay1Ynh
ZqMAFM31L43bY4i3sYxvRSOkpv41UgBWzQpccb/dOsNksjefTSGdjBrk5pF13g9ZqaEE+k3OXe2T
XwaFH7ugDvz7wZLC5AaVn0NM2l6RUtIo5ISO0OEXt7Tke0H8ZlG06PYyhHcsABTMx7DMfAG824ka
vTsqx3nw6RSXWzTUGozwI6Gz5EtwywMa2Hikf4LFQM6BHH3wsCfOSbOAz9eAfCe6ViIZCQmOPxcF
hEalC41V9FtcoGj9gv1WS5T49hEjWQCf393r/6BMgAjegY6SKOtBusm/DH0wr+frNVD7sl7ITPHy
fyKl6Y83oAYJiSFvjaTcK4KEPQuiv1gFgtGyhlcFQKXaJ3F/2BJvEBn36+lkPea4gLSfCn5XLrIS
IxVsG6u6d3MbkMLTOWTF8svpOh7Kn8oxPP/r3w3L1r1hbcWweKt86gNJCJok5JZxwgFieFO20EWO
c93kXNPH/YMXgHaW9Fyaq3uMPbaSXm2zex4/dgq/PWUW4krcndVM3X+ELjI6M2ryiN2ot3G8jqVF
DoinnR1K0g7amEUnUv2BgqP/THidgO45NyB6qMp9V+DLYQyJ20rRBEDprErB80zaJxzXLUAVGvU1
3US+M6feeiJ549P5Uyw9xIqVFNFb8z7PBwuf8rK7eg/l9zFEX7XymiZvAKABHO+9oFNroZuNnedO
nbpSk9sEzEIimRzCjdWva/n9m0c24swPPUxtTkS6TOfBywDGehlNUBgDvmOX9ztL+vQL1fYlBfAN
j94BRquoUWe4uXeZ5ZE5B0RosMwJmceI3YjHfsflHzHiu5xzs8OYCr5RHcEgPs85krsI2szFhGMS
h4rVsrTRLmzQHEo7mdtWGpbF4iCba4If6GUIgTG+GalyxzbR5lJEp2Hy42C0oJ8/drSV+BehXBby
WSMUNrYEcdUc6u0JtuzZzsIwshhTJyEEd/GMkXfXJprKCqKWQPeVfat+mFamCZcvD02l1SWoGSWv
LvlRNqzNI19vn4yd618EgtGQnKV6yY8mi+1A2Sl4Ms48mFnZP9u/U/pGu01y/izqB9IFaZ6y4Zcm
rAD9PzpubG/w0P/3U+uK6cPquTVT7oDS9YjF1vcG47+L1Ignw5a9LX+bAbcG0OVo1fXFLI3McU2N
/h1mA2tYaE3nDgxvoefBFxWDLCUhCcuHx5EhswbMnC9ZN1n5/xnjUtre941oamNd++LSG+i7NY6d
MuNL0Co11IU34AjiGBH/kWMK5gqi2YYfPYUTQ1k9/oHR9G4eDMFNJTV43ePQsNCi2IjEn6mEGzfg
WdCoxsW0BwdDV5WG4r0OTB1t6uvX5eeiuPHQHHFCax3v/T37Te6t9JzoINBBHc5ldpWrcaXZiS0a
M4t/Poe2eD8erlpA6xJcUuFWOIk1QXiWTNUFEewOiJz8bzKRZ9j+VXJRb1FNLsL2H3Xa4E3FWk7a
/xyAyqPdPakjZyq4Il7+YPF74+TvwAGDIcGp7c1ungV/dlzTxtqqyF4Fbcd2AwQyhJQO+b0jZTt9
EJFqKReEbPJbWNytZnWzdKMjkhEaMudtrMYuk4dBSbvbRdj/8MNG/1F7GhOlFg6ySP5YoCeXcwPi
r21YphHA1UfMgYnbUE7ydZe/oKp9sTIoHgchAcKC6EsuWkLQ6bwLLJHbNzkQCLg6ugjV1zQDH8Ux
RtWvBOXhCUigRid97O5ntlHlzmVGLgUDXWuQZvRHpIGHNbB2BlE/HBdqYj8Z6sVAXKcnC4IgUkza
G7Hdtue3NwW7AsltJSlk+CgVi4IVASgZsaHY50gqsfGwxIqKJSXzhj9NlA5XQJIOQOLVISWZ/ZB9
gDudM/p+Z3oghNcYX1tnll4ABc2PweFv2wldPJzhMFF1ARozMRqVryd4XZUguEaFP/jQzj4CAOab
IN925KHAKbAkHcbfamjXknsKtdm5eZ0j1emMh90CJNG0MzN78mEZImbFsOpQAhTqG7j37Z7xklDR
rSQYvPEH1h/StIi8DB5E/earcoShz7xu7PTzx03IvSmEncg4RdZDlUyI4XcwSV7hgAVk0+gKWIgz
eVqZuNFyGqPXWne0xTxsz1+9pXmhmBkk/T4hevb7gu4KGFJOiUSEkEbLH1VZUP18y75hm3tBEgdt
GxcnHN8vtJOSHOCyVxdAwuJt0Ry83hAuw8SLSN1waaBY2tlsVqZlkevzSb4d1MePyXXxRqsOWs0G
IDmT/9uEPmunfqY1b9CjsLrV9iYvLZBjyj3aL5HSxIshvZahfSTdouTaaWyk+06VkxYDhGQ9YUUP
yeP4FcKPE0IMgqlH1nbgnDI6aQUjM8IyEGmD0ms7OmAZWv86DQNryRCEfrb8X07d2d7Cnb8ucsqc
x1zxEFVSgvVXAFSPG9que245lHz/NeN5mjiM73JZHBibO7z3Pn3wpy6goj0c1GOVhzsgksXt6U+A
tGgRDwhQQGGOIHUAjRz1jNmgCX24wVH103okCs/EiJXzu6N6QW/36DoZ9yRIUs/ilBbEZwbvLibQ
MQ494zQZ+5KSLYxhsd8E1VsSEGdB+g0asoWSVRlEFwcO1zu6vhP2LWToNaVUeg08ZQUt5JGhu13H
96+n2IQ2FkafmxEJmdw58KX75/sOM9wgJ6l89fqV6vyEngjb6s81AHU//zoTo8D9pobxj71g2U1S
zZ+yz9fUhyR3ngk5LdWlGgVTFoNYeGRHAKOIcahhp2R/Sl4kOzsM9ne48GNtw6RlU5DDdq94El7p
UuIR4c76vqtWQYlQHfZ/uZxd7hrR71/1WkebjKnlk/+ZF8tlV2BajgDt5xxfy4asFMGocNSTan9U
xBsR8WxnUgUH3PQEWGZXsIGpF89MB/4AWS7VC8c8iFoSDkO6xmd3nmfuY+CkkyAs72m7G82Alxqd
EUaTQYDzF5ABfMpWzojCuu3QZ14Jn8odmHcTTXir0ZcaZJBpCkhS2ZflZim++rhYTIo7gr30LSZP
y0zwUwwfGd/81XNALp4M9OXANcJ9QMnGHJQ0Oka2R5EzMedR7QtI33ibrStGCXTHbapCQiu2Yvpg
MTcqV9mslmhrObSJxJ1IFlUcOcOeMqWC+omnfARZHCEhy4CP26JGBzyd13p9GywlzcfdJNgVymuP
svhilUPPtPUSAADGBUoxAV+8kk45EqP1sHRf/x70UIhFvNh+jeA6bpQZT4zQk7Vv1ox0DGGkCeHJ
wzJHsSSXq7s+n+6zWDW28iMfpIfXa/wzP4qjBVNXaaEkB8JbbOBzhiZlNezOi3RmzaPpqbZyH6q5
1K5ISxqtLHtP1K58OjSREEjQZeV4swXgI7EtRrBYyDzbBjq9iaC90ger9rOjsDT6Iz6ZMFlQe8YX
CCPyB5mP3SKo8utMv6jBcQyukhUzxKRYAetVqXCF+PVyTqLEwwMEnh80aNLwWAkpshNTYINAMwRA
LL9TQE7n6TJGpE8XZ/aUTu1CvvvHV74etp+zWCXWF0f2ynZFYzpdaCrlkxaU8W6yXOXgiAiKQqs4
xXxtyNiDvcUt9VIN4F8Qk/1OgLma9MofGs4GEroHGFDOjeUnnsiEDNthFVNtDZdM705xkZqTA+vi
bysO2sVaV0nT0Poq1wCKilwYCevEC6VLJJwB75MCwI66IvAlpmfrF52FQC4UFNyW8/Fzkqnxvkva
/HB4R7Wb/TfQLOMnQPZQQqJAkheICZmqNDX+k87kFHK1W0/6ZgKiWTAj5KyJKA16uHFjOM62nWSQ
8xK1YSuBEk9UlRd6u2TYLvVgHmtWVaD/R38XVva/BmMX4D261hLgY6N85LYExiySUCQBeysVrcDn
I61kC0irCLf1sFjU1TfiMm6rqUiyX2IXtcbMwvdrPjfgQ+C5QSfGq6eLg8dvJbOyQRTxI7+I6tbt
IelyuuSGBZp5ELU0uYRAojakXsa7pc3mJir/eiA7S2Om+lzW2D9nBTx22duj5aN0r8NFAMXY8oTq
J1aj6HYJ/SaRzDuGfm0CNMHNvC7zMnNrLSBxg667k5uESmYqDI9wAyUhxXD2oebr2MW2s1g2Fb2k
ZdKhin3nYE0ilratwDRc4z1YCv/wWFr9fGQfeMF+6t/fyFC6PTOaxRDnwLJHjDlz5ofFlrkxSPKq
cQGscRq8YFRz8rYUGx4JUPV7nRjVWK2GCfUYvie5zg0Pv/3LCSe/5S1zpoolI7i/ZRD2vfqY4Dat
1F9CH5aaEQ9jQI/cvD6TzfgQpdwSHgjt+bvURwidCldN5Sy8dGeV7eSEUqyfYN2OZ+JQEpaPcBxy
3WNDTvKKVcl5Z9OpjZ+kL9n14r4pUiKs4eTatLoVhhuzlNTP2EZg4u+KoEi7haF0+dIFqIk7M6TO
bPPzBUADyktzMyk3bBenkD/Oj40KP9+WXAoityzpAhB/xFQ7ArbZo+jKniNxtI2aGXLo6aVNj7eY
8D+Rnu4azVQKBr0Heurv2hhfEOMSOJBN3iLQjJjJvbgyXWjOZNsFzSLduFfWrQ51d95soBeMVsqk
bnSAwdPa8BBsEjDL7/Qtv7bj3WrefTNQ6o4167Qpu291In+BGaomT/A+c/IeHezeRa29EspRiES8
Mf48rYe5khKOx76cT/BFu5AtpCHrUoXw8FiCpYGSkmq0zEywlpH4ofxw/oKILbesstAvXVpcZXYM
o4s7VUaWpkl2wqTHQUTlc7mfJ2cQK8BepHgFogBTG2rko1sT
`protect end_protected
