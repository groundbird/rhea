`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GVR3tpUqP1D9tNDew5iD61F86qRypPsSkj5QVYxZA/F1uzAofhHK1aXv0F6vKNSsS6JPghF88I1H
rM1nqgXQww==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mmm1Pq3qArHf/jIhaCq6mqdek4tqRoxjIXwmX/UwoGHa0kgpqw9xmrl1KZCzzLLJydmwjSDgTFlV
mr589U9bh+EmmLK9uqWO/NVl3pja8a8GEocGg4gm+VJMOskyZ2EnWaHVrG6IUp/EQzrlM0FDQbu2
EZq/a05s7D8woIGR3HM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jD5U6zH8NXmm+3dRqg3oV5ujJMbmxbS2TpKG8Z4Pqp2UnDZ4+V2I5JI2pz9X36W3TI7rI/jZSsDT
V6eAewp+Z9ggYdBGMLrp3vS/4hY+An/aTBrZAX2bt7Q1iDIR5cbNaqzn+NSKYGRjzzx3uFlpdRkM
FCqyqM5RKYzUJqsR05Nz23j1McD02w71bAqQID33x+z4NzPlz0PG0w7hQcxGYUEPw1ZuIxAXQchm
FimO7dOAtsKoY7WmmGlZAEtta2h1IvtCdqnm2oq/gVSOjgPF4FwJuRwD9/Z3EUHnOqresSk18k8q
nO3FuUThLWCb1Yrbc/+nCHDlDDi0s6eYVQ37/w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Wi6cKNdp3k34AFvSYKkcflCpfKrpDHlpa74x8+mfVoq1S1+O3D+wL3HL156n26x56Wc3MmsQ1WoT
M3+k5XRVb51ydqZ6LUEySwxE7y/dTTYuYkUm0qgS6T+e36P1LQId/LYZhr+aA13PyJNWFlWqxNY8
U0To7NHmCqx/UDwcrcg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aPYILVcRPSju9bzFnAdELiQgmB1nypc6O+VPeNMM/iWt4nceR+1cl1DvGV2rukOC7tegbT4g9NRa
+jXFqyE+jdj0NLejps13j1RpuR78w5WER8LhNHlZChP9bYZeraPUfLuQp6nfQ1iAuB1ChKCW5YKL
yROQmn/uQMh+Uwdvz8uO9gSj2M8xjNpkkkYqGDISnej7Jtnty4fm7zZ82E088kee2doQc9W4DvEj
8T9IbPQLyAQULvB3cIZHVBhxH4WJaoVzfo+3Gj6qlpNR6uL9HFIk9VYCKJhL53buJ2rLPiweOPgm
Wf4akPPkSo5tphBvbcKEDKNOLxq8HrfHpcY7WQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16896)
`protect data_block
X40EzPOy0DTCJSMgwe8juSduEmfWyoL+OapjVJ1dpSXxV/l4VNM5DA+hUGhJ4wY+yfBs2pT/sP+v
CWeiAuXrxhVujA8XAVn9fMn+ocOqWhhuWq0jwVOvO/bGVvsnb70+bw20tDZf7kxWQsgcE7sk0dyN
yfQf22ZjRqgNvZVJQcj6XG5KRyrfzDef0WwKlldIkqW1S9qkKCGC3T9En4V7WoIL80JRc08wkzJn
+hT1lycYuCPsMdWZ8Sjgjvy9TwwWENaltAVvI9HKxTDEW/+Y0pz1qUNMimTBpsXW23Tei82KFGdw
kGtjUX+RRTuSRaULlR3lkUprp4NNSxcEbrIfWcHfCDOKtjrf2N5uCBV6x4HMp2fHaTiyjs+ylOUn
LKoV0MMHtN+tVMAqMXpBx3Vnl/C6izuwGibpnLTcdYjKgb05CVEA/RlnijRruN/WDczxe/ObUMCE
d1J+NJf4vqYHwiciAfKzGDB9MkKWLUWTW4Nh3IfiOx8V+AGNXxWIBbFBrV9Q08y+LKBvEvOYXuUc
my43TnmskrMpmEVKTgLFiUZEcmuOeYjFvjLH1GHQTRoCKt3OiqdUSrwkiL34YiJVcY5jrXa87o1F
1ZQ4VneCtGkyaKtBgEfMb+rDjtY84fV+kqRYvtPWSCGlMVgAXDILwvpg/aZv6sGO48OmLBYwFPyu
DErhg5dRnU+0NeC5FOCLwspQXxPGd/ianHF1mOY/ZUBMrVZZbodozqXdiVRHfzqz5yzwkp3WLtSr
0/UYSFQRnEzLnO0jq0qnCN3Sn15a37mfSStT6Gz/n3Ja1u4Ejxv606nWTTbGy9dE4HpDSgDvqTdy
1La/Ts30EZfH4Ptdguligvcg8uMibI5A6XAciGMKlGYT7ayouUsxmW+vwYs53Fqb3HG7DH83Gl+x
L5DH3sHaXnuBVXkJ6BpTGxiY/uX9J1uq8eoC2lj6Qb6Mfw4AHudSsOmU04Gn+gvNBpwI+WmBS7JG
Su/z5lJgJ2bcDPH9d5YX0M3VdlSTMufCnsbs1rNwIE/mBUm+F6l3/eN0vlJIlFn9V5rVUyAUKGXJ
YXwnboLkscACfvS31xmY5qGb3V68xwc1o+JxwqCeYuKXTEOqk2neZbloxEwTg3J6UDFdCKP2cc0q
kYa4RXNW75Pj2ob/o+JaN+crJ+jpq9ob0jqfAEmR5PFUoafySsohh3KjEsVnJqqI/moVV4k0sVau
RQWC9GJNziDKSVT/yK/AO8GVQVtkqw3phqE5QbBM8bx653v8K3WvmgUGtnTF0VrCU4vTFnXrGHqK
meGJ2FhSWAhnR0kjCQaGAvAZKxd/ODO9WBIjrj+odYkLXslSdGec31L+pFdESxU5hR2VEySSmiGN
XVq09e+30lLnT7cmrd7bspQUCdhrHHcMMZ8pPdsyF29kbYcCmoJgiu/03fcmiIsOG4ip0tL3SbpY
5jktZdwx0I0FQNI5N0ZAYe4boo5eNgoA4BrgYbIi/gviX7Pni30dLGITrmm4sOkZ6GXIgQAsam6X
yZcHfLWx/7/fMGYo3HAEf1xkY7vGVhh1cQKdofMqz7Lui0On/se0WN/tGmzftjk533C/SJTiCd0m
hmkgCAJ6OUgaKRL5mrxSpsk4AJzNWhXnThffIAbpG9bnxLMs3Af8tkN4Sfl7yhFyWFIeX2jdwvnC
0rOIMiMKvfwOcGdiuuYeCm37GxcYYUC5DCjIHMo6vZdwQNTepn5EvnMkcd3oUZGnOpVtXmEF6fsp
Gfu5MGxlzzVb3qH1MDuL0pQe4BR+UvTjRcsUVsT/b2T/Nm8NrhQkmYON1OBY9hVA64McIqwTGiha
gRwMJEPDU/9B5aqoOJ8SnzeGYNliI7GitHkB1/0qruuFRcBda2F86mpyAxl7/YyNgmh9QibR/NUp
Z40MBmtgt1xCwIXvQH0xksAM1xzz1HNcGQyzbZrJaInMoLIgWPg4oExOrS/t7xKpc0qO5mpBH936
q6KmB0iEgQXJTj3st4Yf69Bt8GgZusBxI5yMZD/RrzbroZncfuSFhsBVR2NmFFDg+MSOVQ3O9R4q
8Dz3cavNrpAKlyCzV8hXRhvdtQIG0Vs3dUVsHJTWSuHrWN5ttDDtlILx0V8AaosftDR/yiCCmNKD
BaUGpqm9E+T6QnDX+zBTYiEoKEz6ucBpfEyEj2PjFfuh3ZTl6jr6EEcXRKytVPqMojVIhHIkh23b
JGlWDlZ3cEQK/uh0qDorKqWuUjZfCi8uBu3urMgaDdnrxdXYgmN3rCXm+sJqPOU7o40tr0FzY6Az
AI5G2G0qAq+QVYvXAUAhBdo6KHMRxY4tiQg+3W/w6mFo3t1+alLGDB/bobUp/IShEtQJe6asoBx+
w/4q+tB09V7kI5o09csIsG5ToonxtD3RISjQSj3eCzjGKn1SFIOaeMEAxQnMYvFM0Ar8+qMeMvdB
tax+wzmI1+NXcctgk320J1cka1xVE9uRDGHOwkCm4dBMJHQhpgnuhphGhQGDbrUmZqwNezLOkCVQ
WM1MnjFW7kFrQhO3xGeOtAZy3H2A4NBHjej84LOYwHXG/eV0NVYI3oCsOCVCzUBv0171fR4CgACn
9qQYGP+P2EZ/CYibtFm4m3w+a08fugen/oBtnABZmUH36Jp8Q4EiiXqGO7+YPkCWKiFPXQ7OstFq
AAjNtjeTHxiqgEbDHBEHldLH+e7Bv+ylIS/BBKPf0jZuwV5cNhFcg6190nRHWVxS3jM91zJi5ILp
i8tE5ue1QcEoS4+LNC0Z16BejoVlWTYiX72+qGXRiM9VKkHKMzrZnAzqsNQ8htM0xrHdNE98EOw4
O2dbCXok7pAyzaw0qjcSOUaQopObOh4/ShwyfDg/S0MS+c+5JhTIrntX07gv1yODi4VsAdlpS6ys
NID2MHh76hJ3Zj8FpPaQefnmoXuGZ53LRMnix2xXndwsPTINbpo2ZkFRLil8NY6+lSNOUn+o6kXG
RLG24VoE066aDs6HlcsI8liDyHeuOlXoobqwXOCv31XRZPrr0fQBHALpq5yKyoAAJcDyW9YgolxF
E9ePyDx5OrAAutOHL+cSoKS6HS7m41elfjSyVmZH/LlM9CDUGhdl8DwXIRq1UM9Hp4uiJYFlDINb
zT3lCzfuiuobq9PiSNF6p7j/Y08MCQpWZkIrp3hwhjVKV/KhVNZhWM1PxYA4sSpg1N3smlTAytpp
+zNUWzWIkChl0N4W5xwP1JSw8gOoxGiEGRsbco9OTPzg+79gd+bWusYKyhydhkq3jpgZkBQbXCCH
ggPSkuViP9YvAn7DzsNqSWeW39K2FuBq/IVy2Fw4AB/ldW4fBlWrCa1eORTeWBlNqpTq9WXGrMUS
WDXnWL/Ii93xrL6XYD5AzKZx/c81bQaLjyfPOv9SKMigyMycuOstw1z6FXv9Qj3nA8ZwsW89iyDp
B7y633frheS1PJD4mNKK3DfI8O5KCx7UnJeUZOOvTtPgc335EgnWmx8Enh7lAbDqYebQU5BJojpt
0WH7mDEL1rmLXFjGF3LDb2mHfyO7RhLhfvuNYWcD35G6Bii+TLSwxoCpBIG1qGTc77fDqjQSJKy2
K8GW+qu5ddNMNSco79ElBoWiDrKwywUqxJRIATpI4U393IwVEuJ0rZMdp7PvanCEJkQQkFxITaHL
gqmiroFkaNpRoJ1J1xsN5yVSzTNGpPi7Hq1VMlPJVkLmRJm8SLLm2m/mz3N2zT8Dgs/iYTaYYnnM
GxHMki8miWVFsdxDdPshltf+4jG1D4cR9S2Ve9BcDUtHZs+ZAddEanWDP1guosW8hjrQSAtT2FK/
WR4x7YQpHAhtzJPS135WLIGrA5lpalaqhf/qBW4HPvv6vRkVubZfzoAzLKOziR+8VOWuJlC/ruQw
o78/MZXBFKxjeQ/kkb5XBE9hGMckW6vuL6jAhCoPDr6UfnjLDOKIp1I4xsbnO2F8aNsBsiX9e4GD
X+cUMx2NadUf8cRHS2i1fu9E3RWhdOVJIZT+OsC0J2U/vuAlJnfAdqJftsWPA31yq+BPytJHaeH4
ymXG4kCbzp8eOWIJXN2lMkrNxuCbK+9PDaJd8RRKBoa6ALtbTGT/ZgLSy7EGxXUFz7Te9c/Pd2Ct
NRcstAzEPIKmOfQsQIuAbhbLFvbIGeyFgx7tu/hfKfHQE0YLW1jm5XFHRXT7akEbgKtorGPXmDbQ
2wGviCHnkEzDtdrfq0Tf0gVe0U6EGnQQGtFnDwgUJr179iQIfbbt5c7a/e4QGD/Iszh1oDzhud9n
acOCXlapUcS/kPVEnksOA0k6Rw9xC6LiAgr3s1gYvJ4fDd519itk8sXiZQuwj/pd84syuMiuJFNJ
fV3qEWWGo5YDi1u6u4rgri5IWuWwtNf06CpFCMOU4YZFfv6zpajHClHz/H64qanzkbeovfZYZqiV
IUW1apSpU7v9fPLStojj3qOJTHKeHW85oCemL1A7kUPCTc59RFevW52mCQnebfjI42y0y9p3yo4j
hxq0LroANwYoyl1TZRMsEMIHJMsPLKCVxSeljnXpsosQLQDIZJ5i4Hni9s7dUkFACQJTnilM1hVG
fBvATRApBrNKWkqP9QXZ6Q1UxqEUVtfXTQ9nqSCztrzGMVoqx1UD8Eg4tN7Bw2IJjSmjOXmJQQDi
sX3xkXP0SH0iaatGk+9jiRvK8B0BQ4doWl5uQKnmLzX2cu416RynQZfTXG7m09FMj/eKXv1IjHxr
oISIZI5IFIgHlfieXOufCkUGFheqGMji8QIGVV3B8XSGJpWLSBxASEhviLKYdLC86E9onXRZMh9X
yj19rXK0yyE11InnglSCzBW+LFo0pXfaX2imUlp4+MLV4FhALsmC31i9A7E9CawY3L4R5+X4a9+u
gBLSMdXpUJSOvXbXKUAgFNiXzQrrpAByKFMLVUk8LRlEAqwfc/tnHTcWjtxtFvW4xCPRIspyJqGC
EtHjde8AyW/UWEX/8quMx5vcDbXdiroKHx2vE1gWGngf6TD0aqfADX+1bjv1OrJhjuzu/QccFf9I
ZZcBh3K4fr2K7PLQ7MTGz/uFGdulbJtMy12ARRhi1iXbV2MFg/OK9+i/LH/aQYqOkDMPV+dOU4Cw
vuPtjChl83W2kUVHI23mVlKLGKpGW8p/XI7slU/Zme6fpdbd/euYUy6W7LLz1F5lNwR72DemI+7C
ce1AJIlcICanNVnnwS+acQVsItS0jpNPa0dv+i5kpzsoMNV1M7EEorpSOAz4FDtRNyAE5flWqKmp
mdMQZt1tC770zZhkB5zY/uGv1iCH7aGMaenulWT14mYw4fqtkLJRSEiQXiXPJ7VHpUCOBlHv7g2v
nPKMzgQiybxWBTKmMNB/BvaUDN399GXQjGXhJvkamEi5Gr+Ic77bxH3A9bKiwch8NP8g9nJJ2KOZ
6mzPwGEWxO2U+WT5XUdwhmHyNuLaW9upbsa+uxgjyWXQJ4tIX2CUuC5og9g0q3QMc/89WPGLAZwn
Zc8lMRdc9oDzI53elWHgFkNtpvhB4bVygi6mhzLilpqUL9WKp9JUEDuu6abBUx4ELtAPw9XmTjeO
tdOPaQ9K47T54NxVeIn3Ijmceto3xJOSBeKz7tYp6Oo6QF/3lC54metmlv+7T0JuWIdjsEoWNs3z
8hQBaav6X4iGJY9tlXLk8+DrJmnZOoMMFgRtKPzesH/cOyDKSFaqA7MNICN83lnh2DEhzq/YvDbm
gb9d069TfZj0INLkgEk9F3VN1NmN5zFqzu5zZRn8povmIz89EwlLOJGLnEU9qTrvYZZ9a67wL5g6
mnlvOFDSnh3Qg3OjxwhdrvYMM7aHMmxWxY96tgKfEHt+wmV/gHvucYS7Y+lnmmvV3N+pI2POKs6v
nTkkOAfbTX0GYNDgL3ZG2+8qvnxW3i6lx3uzOlwAnRCiPZQlSp6qvbvBwlqDvduMKGF8kQpKKFl/
NTF8UqMXkkDzjFzXPIukJIVg+sBUVOUVJxCB0LeO58CRAbyh8KJ10kHKzCuYGKwD1kMQg/iFCZup
sGRg8vpLNnXVoTJ29Vp2rET+C99/EwZHYkf6TADAPOESv5t4U8dKWp3QHe8WI63/eVE2yBuMseSU
43rq2B2ow00Fgysv0Yugi4poNEgp5uwVKbJYK5lGv8oUA4PNMxlXky5lxeULO9Ge1vDtE3w3a+72
SPMWX8/5K2FreY2V3TOx4IZTcY9nSzJd9y09Rkh24iJjnrZ8wniAyzdkLcXHNMiE7bs3HITPhjI6
JcEpJZ6fzLm2iI4d6CY2dA0KLXgVsVGOQxQkiEnYAzFXyfy6es7rmD8GvIJlHZ6iUWylzKMl8OAT
HjIIlBmKgm/OjmB49JOnF/bi2p208zBnn+S7/d/M6Z081GdcyI++DH2/CBm+0/NLwQdEup+HPaMp
QZSJyaAYNx3T1GiMY8EJhQ1kpaIgIGP4sUXnggX7lZId/ovgfKaVMVJYQ2askuL5njXSse7DqdxI
d3QAB4KSHItbIYTv+y7YnAhEckZqXPkMm1PJ2lH66AY+Uij8QTpFcCIXnP8kp5RfuuneS1lqwGv4
Qkqv8+nddZg8DowTQwPx9czXq/mJVpvXYRkrIkmBXtY3qwfn2snnGemooUU0xxOjeWL87+KVpCjI
+eOwa+5NZOIBZ/UN018VHMkJNEBuFQ2OfLrXlJDRsXb0rNqYHeDrVpJX4X6VaDHV0Qxi7d6qI43m
I0jwnjAlP7Mobne5h26qZphrNOQ3dVywncJGxiMosqwzg4H3cjmeI9oC6XGeJjDk5Ka+xi/J8foY
fKCp3BCF1dBWcgQs9SRr2jrWD7i++jpHGDKPyZxEFn7yWe8GCVo3/2j6TkO94vJgaDO/h+yPPu0i
Tg9VI1h9k+o0DPqucI8jCNPrpSAks2IwTQRUvmCikxEa3tuSbdT0GV2BtwBGIHNiUs6jrYxnEqdr
mwp4VlCjqCqea/LDPK/3nb2mjIDG3EQWoCpwET9JADTeluLnhmvlFjZBRNjS5nzjZQd6uK/lLtTf
/PacZSlohcJCM7OBgaemVg6Q48ZmRwxery+eUNJkh6alqpvY630MEZPjwfwgEbbwWz/KMx4hMNWI
Cs/LCXaSmZnolkhEHp4S2LVpYPT0sra2GDQRXfWFo9AZOHlrUTGKve+loLHoD6vEPQktD/ZbcvEE
30zlhRkc7twI5R2pkfxSmJTKttAo2eL7QYYjYmoGFfF47tLyMadL/t5MBJ8gqWQoVyovZBBAEAZz
bQugAdo+3QigpDA1mSE/h4T6YzVSq94hhH7XDKzqWDU2Nm1CPaeZunYnsR5GalxxarbCDLqtL4eB
wcWS7bS06j0i7IUcBylM6a+MaPA8xtxJHxlbVgLzQJGcFkqbW/ximKm00TWNDsBAcd2UrQNR4v24
xC5Lhk11gdOFvvnIcOU7C798YIptTOIVcOVY7kczDABgs5PYfwHPsg0I3p4vM/u7FaCWYJ163n40
wlFl4kOzesNjYg3P9G6YLqVRk/pfrdg69yk7kyv3Kk1Q/kyTkz8rd2FvLWO8/tIxNBJYq8zHe3VP
vQl2sEeSrZiblsSJBgk1kSqO36ajiSKrSDe4TDbLeP4MLATamOdEIu4UZUlznvuyOELS2KXMYB0u
uFLv5jXpLSEA5jDscUuN6DJQRqg+AghvBs8qLgO6Sqbftmkh3Z3KHbC5kNKR1y5wIJ/XYxivNYG0
6pYtMhkB6Eswh7oFEjEd9j0gU3kE5wNoEnEcASs6aC/6iMR2eXKAjTaVokzSiZFUBypRD4sw+O4P
OeUpqLZaHjjwDqKO2RUb5LBe3i04dZ3YH+0wJrGpKLG8PaKwfQ2CioQUQEDuvxgPpZfAYTag/3WD
dQKK8gkHL0MqeIu10MOyHUb87OI9u8/FgbscaOCaoIuSGmKjlBKQGaq1/ZxNDe31m429C4eZuhre
A/BVE8ITGvfnUa9FsA5IDidmbxmdYTDZb1MUZUoO/74AXUhvhY4LEvbydylzH/WNFIVhQoGZ1ICn
kuHSX06CW0foeJxsoXka8/vJAcqxqZuaB+CUuVwa/iz5Vit8o2kgRv3OP7rT4ewLKfE1dFe3xlAN
/ZKqmS+ZS36sCWW9U+PyV/xDfaylnRIqPYC0w1ipMfMOoMaHlYjzDRYwL+gYY531tt2oHye/DqxY
RRkp2ta9N9T5OeU9u99FyUhB12OvlLajcAqvp1+Btx0KWNONc+bZpMX9colWLyupCBsa4+x+F3ig
bPrEMFX++R2izaiPrQhJ47KI6imJ5UPEv9bpUWfPzpzc+VGsNtakX7imY6YBUfobaaJEvrmn3Pba
/gcoAyT3ZMVNAVM6A9ySar1Wl1H5Vt9hc7AIgnO7TrOX9EWzrOyZilcQ+QeXQsv2dGg3AbuREEBd
48lVLA85pClZqccSv77MUGYmtN3LSQ8cHdVEg2RKhFM8TF3Anblzy/0PAOB4nIhiliYfWji0p9Go
e5Mp1kmZZlq6g6Cc0fa+u7fh7r1OOt/cuf2aAEGmucrXz+sm5Dc292XPzFEasZ38xt5FSa3J3FJU
T4e17kbdE91LGGgkUUMdUnHsWUcu41CuXFV3ZsVWKWDXsaTswUgrQK7lLST9MM45G1MUC6OTrv7J
Bc4bD/s+2fpjQdlzFek7M4OySaZGDmiej4IRQzS41tl73B2ifdgUTE+KdmprmhXDlSees/5JN0DI
tb4+lVgRX2RFxtU8Y4UU4GLSS1X/CBcY+jolRpz22yAzJCFcakEpruyFwU+DpquhQi/p6DIc9xOp
TKfYDaG15BWE6w0H05OlbhwQ+Su1SB7iEA/6IFdcMGqh8Vwm5xt1zjZptmzaY0rz0dAlbGeV/OGP
0TmxT0EYl/bkRWBarsNCtw859fHp85dEIVU0ecl/YR10w87g+IgEJZJSTK24BPj5Mtx4QPpsodVd
jXepUYsn9cUoXOeteu4SoUhIxd9k52OpgjZESOiJNCI1ArMjAGS8uOoVlYDO6SxVrif48fdEHDBS
5XmUWYDVpPsYFP0HuPcc7OjBdVvaa1H30A+3ZNiWHeiEjUhioN3V/VdecPNjG8s34SWsC16QTiot
HfZAHqZHlPcYc1szWZAPRjuN1QxbYxWLnuwqdFc+ieJ1IYG5uRMmSzTeYq+XmQiVPI0Pjjp+QqwU
W5k/C/zE+7dLQvGp/QIDbaHP3Jhit3fmEI64XTpqLnaaKtNncGWFAoUXQO9ZmU30VZfo5zTCTO/C
BkegLBBpAvPRDgn+k7pWQx1EfLn/zvZLsf/oF3yFz3MZVNWOdipxy9oJiD9QcCel+Oo6RObVYOEy
iqUTx6qkb8spg+n/WWS4CodQAYk+kArZ+6cRL0ybe44h7yibnuB104xIQG+OlmF6N1lJLK9dDiGx
Ge2PBG7LEzeJpYlXXqOxEWHbXfuSrXzI1nveHZvEyHXLJNR4ZkuSykycpHOK4SBWxEsIpIna+PN5
vWvlTgQgM5mPsabYIRREvhZsszJYW7jQFxJJs0QgfYqnUsvdKpz1bPWhcNTGAq4SDbd+kwix1bcQ
bHqTE2Xl6Z6uL+DFR46IOFUQCE1fjXOl3dGLMRzuhdpdN3cgkdeh+7PFvAXXRWKxl3rzumShjy3F
BzClFRdQgw1bVydFssnThQSWNvfA51JviAr6G2VAbpUwDtaw2uUuiaQVuUnDYYQlhWFx4EwCxcK7
PlSrbmhm53G+bn+mX8p0eDyt8ngpe0a/egfoLJJzpoKXHulEWM0UwZWdG0akc8Chm0SMN7RCNgBU
ch/7c6thcIBprIWQXeR/k+RC/nzOh/KA4Ud1SBI4l6SAGz/GQ6gIRWlaIMK6L44Og678au/Fmz17
aGrfH20pYbSNBk8JAbX4DPv6b/MQUDZcAr6McJkFjo2985OUGX8HbyVA2Z8CuMtGiTgBKgOlj65b
+v6V6sK5+LvfTbzNXLIOmVZlvJXIQHMUxVNWNsP6qVEggVmWWmXmqfI+c2Y3rahCG8VZ0P4Qro3k
rVHxzPjRHBefI7AJSRcfKFvmCLLT38yr2VBvySbzXewrHOlKMnf2xoU8aTRVi6EGTxxqOkqtKOHy
2PZEVGGWD6CnQ4n1204RB8EeO+DjmC/QDPZjT5pb6SykJO7xPtvaOfS4fykkEOjDTdDphdD+kS7V
8kpGp2/97L74L9lvTFAGcYFCNWlgrzT9VNo5fyXSakCous3Pgl0zP0ccgnJ22zOyXBENDNUONnlI
C9HipOfjUx9j6JfMCEHGXHaBxfD+V9awNj4nI6Aymi3sWT4zRHCGwtljTtEswU9ZNYYgfExRhShR
I0Hvs+xzM5TyxaOplaK45sOgvpxLuKS44xDhIOGl6Nzq03XYrCfoOi0EJAVqvyRBNLyxwKcJlRE5
2Nzxaef8pbpiwnG4WAJES/M818WD+s9m1K18t0KSvGg2+kRCQZ5rfUqtIwlHkLFqu3gFozRUTHQj
JmYudEqoKg21LECqD+X3Y4F0DBwaTqZTLvpmj9Bj+m3lf0VMrX1baLdc5XkCHVfTlc+OzoQFueEi
HR/FcnRh6+mPq99sZDE8KH/unAqahJDudRjPs/bJcPfwABOpOR6n+qAmlsv5xJ0q1gu+DMNAQI8K
bxdHyMFljTUpntU2nN/Vz2khVBUPZvEWbiysihLHKdUXq6kRViaBqSUPWvawRFS58B8NBOBWh5El
mEXoMktquOdevZ7kgpxRLTalmLbP74HMFKnBnQ5m9oI/OfrA7v+lqEHyVVzJw/PCkd+j1IbVTY3T
GExT7FIcHgNgodcnAfF3X+gw4aFd6+r7i7LQeaggnhtQzrFyDZ+xrfJ4hHnBAxwfuZWSRB+jDtfK
kOmWQzuP+3oa598uVpdzhPdSweMqHAEm3L2KfOMBqSWSEpTpGfDGbMzJ0QKINMu5bw5iGc4iwfvP
AmCVHQhB3fKTNiCCMA4O6tPFBq8t9dQMPdpb18UC1mnQ7k7tLpNuf+6FaTBqRSvFaAHPild+SWKd
mqZficgJiTOt4EoEgQ4+8NmNuaEnHaa3L1AUEwXz8xAok/xx5OwBTjcAEAxS4RTVJbfJFDl1O/Cl
ncbYX5fOqX8dFmbgMLIzBJyYRBwmpx/hpneXifQ/vEYpsLPspN+hGczqq71QsMR8nOf5KmaZfmZa
Ddm47chZuuQmy3F/68QtPuJjDrXuwKrkoua0OG+RSN+Jovz2Mjf20+dd+KK4vEg5lkG3Oege4Rr5
k9q0ZEcNhHpe4TFfN60YSCc9xFOddVh78CEsctJM2sL1M7YVU5zop7/1WhVEt2jWJMZV7iHPX3AH
QMBSftvO+Ul3pds9ar4CcEcFNNwbklmV2XtCvXHG9Mp5tqV6kyvg96Z2JSSYu1qDTtRxwWzc1Tx/
8JxH6+sqKsP3UnCUEe+mxNldEoaIJaUlGYcd1CwQXuZcS7mY7oAQYWWh/f4lAW0JIzzA4gJ/M1zE
tlVXI0Jyg6ftdvz3G4FWSDsAPImfsSkTqTg6vrjp4n8Wz0LqAG4tidkmWF3sHBqqgOt5k9S++mCi
zZ6lxjXeem0z4xQK0sYiAGDUByAkO84hkI8g9LA/WcrUNGXDzAtTs211BHWMEvW7SoPhB51hDVYo
Tajm5dUypjenXEI8W92v5g51DQQWfaHLqpDD6xH4pE3uLZFp75tkOt49i7vLa7X1YKeqD/rlHUwl
75n+QYZBLZkFpaUR6Ex+mZcyt7OMiOSNISWEsRKJ3bLIA/My3yHtDoBxV4E3QlFIUEZbR/zvnozM
AJovV+gDJdXHKg48xS/kOpIov6Ub3QndiBrrh5XWx9Y0maNmqm1TjE4KwWQSC16xgdTeGjgpqsfC
pslx/WPiFRhdTYSqY+SGFVT1vDMweg3wLw1vJ6KxIlnNvuZf67uQnC3Ps5kxKz+ThktmkUR2oRfI
Vc+oHCq8cBeXeGiW26diBrgZb9qA/xVRtuAOGz3xizD61Rd4VXs85pfrkwna1nDgNMfx7e+VqxqF
HGncyNI1ZPJ55J9O+QJxpomH3PcNV4FpToLBZ7WlfA8pKi5TMCzjbzjvqoXwJuAJIIaIrjMfFlRs
O0SgJTjMzks6tGrlLXXC7RXcNbVagKQAYVGelBnCxhU4hrq0mdMmMS0Bedh9Dxk1WR4ND/lgjf2P
KHwSSccZCY6KWmIYxLtG+E20jAfopYGo55+E77fj+yD9G49yf2tiOqp1QaRIpIXUpw5zuhIzYSTp
ShRCQKqOjFDHvwSwpzzvgLgJgZUrgVdHulpqe5HpZsxNQmhKnL4+DrstbEZS+c3eFW6FZRgo/t8e
RXIB/zFYxKVoUGLvDJAfOs1DJ7nlhk6Sei5tQZ6sgWFFqXRicppMIAso/1zrz6wWGeJ99dkyetCl
7FdEtuoXgm91B8Tbule2q1R5TaEAMsl9ZVP/ILGmLQayY0FWj+A//ryHWo7HMvqsxMfr5PzxmA9g
55mTodW9c9sy+2RI2AufPLDdzw/mgE2NTexKMoU2sCxODKmH8n7koQFO6cJxY8c/T0cQiv8gpqzi
Uwpqxluw8vT+j8cHG++6xD1LnAJ/8s6hI/xOvfOHO+1B57u5mNzqfug2eSo1mzK0PZBLfnBubRRz
/uq1DTzbJn0EA9WynL4TyK9eilZcIoZSrBYhXuo4uVJen6HC0vYAZ6Ue4KZYMolZ4U2tTgwpVrIx
atfgKjFSZtxZwgheiPOpURpkzi5GMm+57ElnLFo+nOPOrlFTCxTT7HaUNzut6aiJWpuJp1qsds/4
k3UUgQfTIVulkiJ9K5CyeDsf/iK/lVRoarQXBzEelXQG/RZd+VYB3LZMhTskwrxVkN5dpfAIcgyy
BHtph0FVzEFtxzy7vVxgoOVn8q3q4n14mBGLFE1MK5/OrXMRYEmAfnFvjHiZm0yT0x/VAzuKLFwR
3U4sKmaLI2s5wdmIxPKfAOh8QJixzofpJbag1MwjVq0QQwbr3I+Zo/YoMc5SVAgcOfM6z3CLEq4j
YPP8aOFdYGdrR0z+3nBIBXi6mn/6o12oR35F/A3nqirtR6GJVeTW93QvDWxpo3B7P+SkOXsbJPci
PZrOyMVpWVl8uEGJpEzh1K5XYqLWd0me3OHySHD8aGAecyq98Z4GTkUcqRSYOuaeygR5D1CFBElV
FW1uWVsknwzSGmU1gMEOoLqK5VYkN5cOmHwZlHJzyluCgGxT8BSRJ0KjcN+e0qerfZmF0SDGXLAz
6xcR+QXANbYc6C72fMG6keqdQY2HYsP/1Dy8+kPymmWiDQgr2241Wo4oVSS2jC5vS2i3VqoYlzxU
o/QO0IHQFbUtvAf2dtDL4c+4xRPMIn4twzQe4VC3B+hiftuV29tBUb6jkq3nY0EPzN08jKGSwY7B
lQEM/jVRGJIBCPXzAhZpFRUKB/S2IuWKFbdnL+/q0mO+/qdOy2HQTc3ITx67ix6c31MLf2kfPAaZ
rh/xGJ0+piR9ptGnLDT5NzugPC0CV0INt4RhdlrkPeUzdRQT0BN3C+DSr0+y94MJqA57iPOrvcis
gX8DnqRWAEyQO+LzRRAcJv/L99jHxbzV5ZTWhwuniDeL9xWr128gEFGzPHMAYVhwc0JoOvjhL23H
3XcMrCiY2YKlwRQxax9sh6oXQTZgb/S0zK3g2W6jiSk33ofi6+uSJouMS1DgOM0R0y3zOL82IBpR
vvA+Q3TbV5gp0MeJzUj8u4zKQ4Y+UrhhFTxOSDPfBwbYdYtzQEOjkeePMROgiwttP9J5la5C3fks
/EBLFjtETvwgMIeom68tf/hn8D6TKAGXXEZt7lr69k//E5izqSpl0fyEnFEP1KrV0OISaa1V+YqO
Y3Fl2s4DVKfppDWOgvZMCjxskAv8i+Rw00Ud9v8AtMihn1jgXxrWhYiQWe662WKy8tn5a6cQCXL/
7QsE5HTy14l7+NrESbFHhb/jicd1uIT5GHElA4JmANYwbQVfTkOEW2Wf1PNY+pg7Y1DEZ73//TIK
9W3HLllFLkoAgQHRBghVN2gEucOn+by4PJsdnfhb6K8teUqsEsMhmKzoWVwR1OZffs7ofhnySDBx
0YnXHHn+4oCYN896+d9Nf+aGrGREwPhwwLksQybDHHtyEhjncoGBxb5r+P5fKm9a1AjjqaWrMGXD
33bPcsWqMKJ0q6JfY/t3wUZmw7IqW1V8LaL7z9oFUXyKed7kh1k515UZDQUhd526JeYTvuICju0X
zsSLYRV4+J1hRmcQF76QJ2i7/XD7h6j0iYGbc0RiyIbN6D6AHWj8dh8TXPa1wkiKLjnu+78L0Vle
C/oMiuvYeblOaX19uVU1ztv+5PoFg2LDKFlpWVcMuiitPYySpTUOItZYi5qMu/n10mwA3Kb7F9ft
vqBOrWS9O8FyUOXe9I3ZknQxr2isvFp9wRpMPwF4DD7TmbJi05MyjBnArBsz7apWKTT3LRkfJCP7
Sg97MnN3yjOQiLC8wbiM4yvtKSwug+rupTtKjCWETx+ZF8oC+s8Q5vuZ+YqFg3tK4XHET/k+WO7j
nG95/sp6lF9ULBFtZigLe1NKwkJbP9HAO5HuEeD+VqQ60a82H1p0L+xpBV2YwSPlyT8+4JYixMtW
CQSGY+I5GotO1jDJpnZNYsgOt/fwKWUAWLRbC1TTvyBc7QNWkufEevbfQtOC03yB8QZsoiMWCAz5
9v3usviLea0WTg+huxGwoMD8NbXgm/g6C/lgV1ji+8+euyHaBjbcY/3V0x91EU+KVV8MiAaR1mHj
8ypcZZLU4DEo0aFR5ASCi10MiU8D5jz09fbCfqwhaMJ7g4XFm77FsgYw5fX5p4aZG5cHQT/eFY4B
dRWptrKJ7zBLXVztrA6tzbu+cjPlc/DX3owjFmA7306h1PS4zuVCrLhdr9oJYaQsfvHtGEAq5w4y
a4mt+svrxDRsUjjw7qHd0a/11ktcZCg4AVW2uqWqFP0Zl1Hj8MJqQrfZPMOm/iuNUpAUp5H+nvAG
rr5Qmfhvpr6nq+QG0tHvvNjJUN3/cP0uthVjKXtflokcIECFPtwNAdNpbCJWZwV1qEw4NZzmcNKR
PHlQF/Zzws/m6KhYrif4hNw1fPw1v0lQu82CqpAagW2dL9Xd1B33XBQZhb7qah+Yx+Q7KomRzRFT
MekvNBEgBbI0U6uZgG18ZWniXFAz1i6XwVBN7gIfSboDj4Q4dcWfqskpMDUQsIlPL6whhEZKIsbC
bfNzS9ucduz+lh18G1RPsyoshFG/isrNQ1Wgn7LjlEFhnnMMqA22TxIPAsg1QAnpBbpCFwDTPc2M
1uuNAddMJgzOUj6YsoxnvixlB1apNkGxG0/N/75M503hcLFvUyk5FvbsdnBTPicUhVrmxTbjCjSs
hZUKmwrIweOGNYVOAZxkeGWBeGMWLH9msJ3at2O8Yt2f8G4Sw5Rrij90Mk8eB9CoMOqQz8WyNuzk
+OELSpwoiRM3ChGBn5CKWT1+W43AyfbmAUeeig1aCB/s5bYkQBPO1SLl50iAbu7yVisSoKqduiYf
uW8zrYhzik/UhtQ4Mq0ajGlqPR7iNBEQpa2++netB9F9w6Ok1fheZ9BXndl0jFCAKbqI0PFvNZC8
u9GAAgYPDB8pWjUvhGvT3VpwuuQY1JsSlz61LY+o8r/h4FR0uXlFeVxIIFj8WMuG7tkofdH44J0D
XQG4AGTs3T8qWZ0DE9RoACLNYJSKg4wgGpbYQszl8JEYIfJSzGqjfHR1VENoAxaNxttb15W8zV5C
n2WR+Nea0m4pllR6Ck2VLStdRW9CqWEalQcZhQpj5YIc8VUTOEj2YNDtvUBY/l+EuovfaPcjp7Vv
NOnzhTr6V3VfcN7OTvdvxzZQLDo3f8CbBTvUCvGkh6dkCD/+kWqBcvi6keZK2UeoExfi+I/daDyf
wGMyYPNFwJT8krMbmG/rqdC1qciZTl6QIcS5GgkXrCDs3NeTu6NwiL3Bvrfr6zr7CLOD+hB/LNiX
MWKwBKCTvk453vdb0uQj2ucpVwUGTKUCLcuqD86qME84XbexMwMJ9aQ9/Ob75oxBtaSQvpeMtKBJ
LrOOI/D6B0RZfHHcmlu1wg/xnErWvLszZKFU00mO1y/9FNwspADIswU/DR6FSozDxX/uZK7aPLx7
lEQh/+NOpILWwIPlLNIokIBBmhLioujVAKSpj3XwsE6r56ebuNn+tkx8acxxX7dSmu/nJTK3ojYs
Iuw6c5f9tk167EdR/QNoZBog+UZNDNPwAkR9fcA2327OeGgSSXrSqc2/6J2kn4uBLDTTle+yvjjy
lPbelRyuK8rglH0aqe1dmtxavnyD+GRfgViPUn4GUEy05AUyugiHUU462eTeTCMCPEL0unGsHcOe
HQS4Q7+DqnzuPE9x1gaoRicuGGlhAyRvTdEN7+JsFQwB6gVwicYmnloIvLG6v7YJ7whQY3NpQPE6
4za5EHxvBjTBfqSnD+h5Cbt+2MhUmjnLjIr9aCef43MOpFQqy92vnnYKHlQtiCgdlznXdLkCeCrX
VD1JKpUVkcsvWxa8CC5Gw5D8pS+E7Er8x/qgoRSKv3O1t0xXooYB5yG8JBT0Dg848jXDEs8rSDRp
E0CMl90yj2rSPfzzwo2Vrp1caJcm9SXa2eJDPRjxZEGIhi5vivX2uZLlkLbhK5XtEc0anluAUna1
VYxMfPV61YwtxfwhQ8q4q6ByF0Fj+GSTxAHlf+K5JDX16kMJ3pq6OkQ7Re7fO6rBx1me7VqBwydC
qibqw+Iu8Sq8K4ZecnVANxGlqYsUZ1W43i4uiNNVTIQR78WOsN25XnjDD/QXQuhchBP5dWCxo/w6
LKicilShB1v0l5QJKCLpu8K+VMPbQnSjYjX03O/ratMNX+LSQXuYbNoGmQjC/ZOmZnlwgE4J/gSR
ay1NPC3AWfYGpNJv0J+YliMhFnRarkbX2NEUlmKXLoZzt6Dr77ZooetLVca5k3pByz3I5ZpLh8as
2pCkIi4SJTzOHvxkFXntK8jHEB1AgZ0/MNx0vxI4gE8pcMWQ96iv4zMSoCsuT2HiUDe6gVlnz2hM
cbSS12+PlOxXQlqyrZ5VjvVAXLIVWrx1Upco38Q96/vl403ZoAsDNzlAQKrALnb5DIcpJ9XIiJAT
T+6mSI8tnoG8oRQGzfvugSypywIfVui7KBL3l+1D+LHATmZHloDh8JHXvhrG11N1eNkXS3AvTQlM
OTqgdXJoKXf9Y7u7gMoY8Aty+CM2WZEqMvt/UakVarA8Sd7xVPzEj80TFq2q3yTmH1iwK3wA92+m
UfEU0WwXN6k+wHx0QV9m+vrE6zgNcr1aTgDh1Stab+5uwMa28WWJ6rOt4zcDMVyhNxpcnKmqXxox
KKoU5jQjpK1SskbhFBloZITOOhLazlmCMiowDtJEspIMcGYvKRxDHRqOwkFT+jdttLPnF9cZU6H8
1cryL9mULPz7tnEGwhx1YqUrFnXrpmISwSadI9nb7xpbvV/bvdxB3kbn79ww6T3nFepp+5kBoRZ8
eYI3WkiGQxR2wwDwGpcllEv9/tl8msvJa8mRC7pqhxFKO8p4jG+venIz5+g/sWaGJVp3EaLUDUuU
U1b8WPMfL25JtHH1u3NeXqQMPBbIZSW+uM943cIlrHsbVZtpPZeaCGF9THx5pGC3PxBRV6a/C9ea
moNmiaIEGNkh5avm5suhdsW0o3kZ6BWLdnBszvBv1jOHmWcdS85de21tfsGFk5Y31mTBfmuUnY3W
dZOQ7mNG2ghsKHrHdxFttRFrJ7YVp8uur3I+uj+RKOP9LH03q5+ISphazWJ0Mp45zXC+/COTlY53
eiC4A9MpF1ZiTdPGNyWAHaoDHhyi6M2vvmxGmUijmWMlj+zgVn1SWVClr4uBABji0KKMAIK5WLN6
y4cQ59ewIPZvH/twRmLS5oWCHOcrphT0nTL6bKo0Hu2tOytRjTNgJAvuGcxqHnNaDPeB9KLMXO6Q
/xOjt/kaNWmzZlvu03RpbvZQDC+8FslDV9v2gpifhmGcEm1pMHHPtaOwMoaknJQk1j53b95YLP9N
AdS1zNYO9xhP+PutjpI88HW6ktmgd1htoYyfSfFgtD8d3TfUelALHpSTpqrusRp9vTRr7zrPVGjj
xC7P8J+XWyS7GQtPDX71eL3x4RvItcZtV6POoJi3/L7y5H2Zaw3m6BjsrUwEEFh/YRAqzqnsqd7s
6jMb6KW0+A8GH9yPuC7C9CEboPEzx++J09oIuMtcU6EWZ3+rRum15NH1rbVwz9o3/eKS52wO6TP3
Bws8b8naF1Ah9jSnsMv3AhoGnQwwWkGrwcr+OHD8Bi2rtzI4Y2x+DTIiGpXiz2RpulaKdPBWHyk/
sTvphou9qsmeyDS6cUaJEGcRdq7dVgSay7sC7XPinLLsEJMPhaRYAXj3hVUM3pq+8LzEgrFfutwP
9QytJElAIay4asXWm+f0FWs8GpFVTo+jsfOwOunhSw2TqVjppMOjCUbObXh9CuwL05rKf2Ul6Zz8
MLuQ4xi/79KXOEgM1DVKQtnL7VRAz7AL9vP5ViOH7eAqNGeg4gyDRTPFV7dwVvmjUJzCURpoivqR
R4t90oLTcPMC7t5UKv3FGnzzM7bMvYRSSnQ6Pi1oo4e6O/CDXNOEWeuE2yhAdCQDRXH757kZ72OC
rh0RAiRLrLpGLlbc0qlZ6b7bFBjP61MWQKLsQ0nODpXRBU+/jf2UgAA2QyJXNmaAEVSHrOJgUB4T
iE3vkT/h0bmcxD7ZWg3vqADXK+xqe2EZsT2YY155PgPQBWlx3gf72lFbxNdF1PqYv9e24f4rHyFs
IF4LZu4XIg1H82kA6L2wy2yJXaQ8KBBdPiMKTpuLxZMo/WQV5tRFRUgz4M0C0ZMPBZQWOgMp3S4A
tc9cp8/Rikse4XqZ01HzI/ZYs9MAqgEpFd5wENjufiziiMGrXPot7iqQaRAQinB+ZdB3jIyJmRp5
ghDkv9HlUHhLM+i/pSxpQQK2DfaFahllfx5CXWM0EDnDiX10dDIfsHCCkCKI550LdhehbOb0i7Oz
I9KBa4w63TlsXO8cTpLptMW3tmufKz4iWU6MkAzpJ4HoD28WvkWH5gE00pmnjFGa6XQSucGDGAdU
P+zkejw9d7JArNqXkMNajwviXcfVq2xRSUfFhElxfwJPrdSBes9w+4O+0pd5/okwuFenT7rpk3p7
Gz1ikCjeHbd/YqdMPCE2IvtqEzXIfmWuq3GAxuBN4k4cF3iXOPe/N2m2XQyF+VQsivDq4YRZisPK
3rDOzQDeIplooIp5PGIjWbwSeVgEv5KoNyMJLtIh/yqUfyRUJhnijY1crEM0lmXd9QBRliu9s5Ik
BvAx9N59qPuAbAx7I2iDI0WAWTtbuV2T46B5oeNFQIFVKhw4WzQFJBbzuJOsLc2vgs3LfMumzqZY
axp0g2mAljLhXMepUu72ObrjHU1VzZxoUgoMwyjQOXRADj566dlkYOmVuYk1Q6iQ6lndCqRiLgQv
xg40RclXfNUt40wdJopolV1Sc8DDgEfgyFb88wX85OMWM0miZF9FDtfwpC1ecrWytD1LYShC12bW
hPPJZuZZ4TcQIu7EEql+tvHJiDqdb7qJus490qkIgWNbgvTJH446ts1FHUo3gZyCL69Jlm3jJuJF
tsq4tyrQk3pgv3Tgv2lreZ228k+rz/w1cPksG4VSKI0sSiXDjaAkkBZnMNkx7G9zjP2Eu+q1qxy+
S6uPgqIOvK9M5WoQBFT0uptBPM8V0FsZgDSTdusBQjDmHBP8R5Qtf0/CzUBa4RyZ5G4nn9BUTIZe
ckL/Ng4aeyzIBlhaCNPf9UjfBS9VPimpsixPVCuZCWXL1o2JMHZZOQh9ajkNS5LUe3ZmhL7TaADx
riwuZlPFhCodKWxB0UsOEFlQQp5eagZhhCWoweYWu5O8OSkyF5bnvaC04vUrwuYjhOSs5OF9v70a
jbr46YhHU6wXL+s1ENCR/yggz/EN1G8q6KzmGtDoOosToahSSP1bTQzNzHPn2itXrSW3L4r8d/Un
KZ6ZfeI/k1NKYEgmpe7b+q7PJqFykJzohWgwwLKXt0apzPsv36azbm3e0BpbG63vl6VPHtq5FZg7
VLQK0ajIi4SNx/PlcZUyiBR2mGd3JYhB7RrzsX8kcl3p/Qk5MxqDxYiLuNigY48PPiA1F6N/I7Py
RBivj63a4wHGWid1npjjBdrjLlng3L07oUCvBSOcNjxNScjHoXVexx4MvBr4ZNJPVSVcjfpTHmGi
c62IW4Cu3zlNQUjrL+AtF4afzSGKfU5JpNTldfs6JR8Ns/WNny1KElpuZaRfmsonjtAKfb3zUBBH
brnjvuhHS+W8FJKflrEmWz26K5erIduC/fCsz2ZP7Fz/sCXHSZEvXiW1ACqsES+oVTRAo5lLMJti
XDGl/PjW4RLpTGNymvswaBx5CoB3mmTh6SV20jqbKyugbYIixAbwyFT4DGOyboDuGGHJKtt8dpSq
2Z2uIOkxVKZ6/PHjTuKufKD+3TdDXoIESETuhZqVNPnS/Uzu6D84pg5PWb9Dmizi1eDzwuMnvYYo
gBPGDBkTNMkeM/bKZx7bJOy17OLb1oywkQFL7uE2ktYqlSImCDoEOzVA1vESh88WiwL4aC3LX29l
m20mfAZGnkhG0ZzXwccZvWOK/votowuQ060Hd7J5/7vzvb2On8tWX1YlFufiWTfl8EByV2LJ74qP
vAj4RMeTNzDUykyH3K7U+0jFncygZBkSqaoutdFEC/0f37GD6lCm9ZR6nyaxwRqBeo0K/TYI4X3n
v2uruJ7bCPYpQSqehPyUvLUA13VvWe1P9UmvaidvPRrhPQrtk2aLshzjYIq0zjfZ5bt+5TY77T0M
KYwHtx2oopUJs48U2Fip2uJiAKkAkAMwKWbgI4Z7pGwt73jsBswMzr72KjVw/z/931u3bU9XZ13c
sQL0KNZdwVdgCPm4EcLYr5idL17U5Z3ebIsxG3mbmuHLW0lTKqd6+VcDNYZXD0W+s1vJYjCNHNEp
G+htWevDslf7vgq2QappqxyAn4/xz+AOXuBUgIIOGYAsiupC7z8iBGjK3cFvif9wcW+OAbUXliQq
s1eeQ1DG/z5/J/ENGgl0KyA55xJxd66Ku0qM3dvszoUYfwzxAYj5VItnZazQwzcKQBUIg64RXqXk
mCiEE0b1E99/0azqIJjN7llkzvIBC8VuXvW8ffbsSbwTsFcUrKSKsgaOqaLG77/XZV4vnVEHwXZh
0rOCeXd/GKWCF4nxsFtVw0l4E1xeZ803bNjUn/Zxocb1lJHVGDdl/qQ5tG5/+3vjUN5qHi+8YgGb
+cR6Da3pbLgBxrqsyugdDI0Fu6eKasubR9DbRVGhfINoGMXbKORzBY7JsUvwXdfekkWMUhifBF+4
JlXHhH+g07g93Xd2NnDGujM/j/2+4bbSKOQ7JW92CmkdTA3H5LS4gMPyx/X/fJVHR6G397CSj3U9
H68s79xQQNav9qK2ewQ3eU/m1RNGqtA8vvOLYNoxrYGHmoggElROJES+wzO9oU/nMVSRh2X1/hRM
sVQEf/bneb+fd8wlYp/vIrfeCRMO2xISnqPX8Tm/67TkqSrrM9WPa5j9PjQmTsQaSw5bvGLeTohO
49B0f3B7i9ZUcKZzDW+XYplZVBUlTOvTcNF3diLgm8f7Ij/THYM1fAI0T8ft0uV2UgB5ZxvQCTKN
U7wCVFJSJNWeImA9wrAOAlJLzo//VZns736mQNBtL2aFUVfT2cp+cMecpkz9w3MHjcuA8jSfxu4P
eq1tkwRqE57bYVxV7jDaeu83qGogk5NbpW9oqoAy1YSxd764lfTTdxGlbMkPuw/Q/aZeat2bGQSg
72IDn+LFnYqIqGOfnIgWO8+fFREWi/PASylr29oQ9J4pyBq4vH8OLoCXo+ifckgQ+4/RN6yWek1p
aW6IkOHc+JXnL1U4PVXeXqbyTgzkMtGObyC+ixiYGjI5k80166esR3khK3vK5d2nQKvYnh9A22Kl
EsPaXSnWceUw02Ttu22lOs/Mj7EfxHwPo0+gBeq4qI2ccqejyjRwl/8ydJQp/Rx6oTFOGkh+4wjB
ZG8IWGNhXrxmysY5p/YRwGK6mZ3xfS2FvBTCpIza1Vp9j2UApN8zlBnptgSvqYlIx64DURWrKGZv
zcKyED2wJwKlet1dHYslf9zZbUZ+53Z2NXvGtixB3DbXpU5lPJuEqNaGJ7IVQELgH1gdoN/v3Ou3
dHl9eMYvFI0Aa3tnz//KbagQEx/AfRc1H2lE/JbFmVIJjz34lWbV5pdqrLsfuOB/n1Ynk5dCyZhB
LN1iWdk8lZm+0Y9wqSNieHhQA4YTEXTDCbGU6RcRNOarvAXQxCuHrM+3FoluuyehSGU8jbIbQvJn
3xsKZkhmJGRUMyFMjDyYdfaTocmVvXaUXc4AH+vqPmvIGm6Mv4jbI49px+cNjM+e8Y5JgtF9LoXn
kXp7cpWW7kHxddjV4uS0kSL22rwQUsGiAnje51Qjn3UHItjxVoGmS4tIh2iRXbwgEGclnv4s2yPD
f65TFs+Vzk+rQ3bxf8UZKRPwI1wnjHEgvPot9VAvc9NrODOTOaTWh98b1Yzkwxi9Qqu1VkZi5rWX
T7h5jvbmEFsPwNtHqQKMrC8J65lbB/eA
`protect end_protected
