`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MTntf+vvcMesKQulwF0lhiRFzw34adq8ah/7Ft76irnExKwN/kZtzX4nCBJ29BwcW9Wh7FyMy583
sNrDyyAXTQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ew5KhFqUWG78eZajA0cvxYl/Iwb3lXL13yq+2PwXOHpUT0LYU9w8GxGqTgtfpxjUbnoucVy1Nk18
SPYHAevsdLmFmdGi0jl/6eOnogqOJQxpJO1W3ug2wZtGMzM1Ei2YPmsDbCARZZOJ4HbxVarTjQsE
9A9Hy+jdJWm5MwbcUGs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PS7o63c+KoLrCE56V3ZnZnaoPB91TrEUFmCPE+x2IBrY4yqY5FbnkGlHm8m4vmviwtG9YOunwN6W
moW/iozSLjJqC/VsOnE4371qhPRfkhjDlU2tRww2WY/6nrJr5mEKAgbl1D2P9bEAoCB5QhL9gEIg
6inRqoWZRkMboQcmP1nPSnWj7sPBRtYUcoVSSxVVkWDElqz/VfJCK2+a47wZUqaQZBCmIjL+BmBk
f8BpAMlaCZ3OgekPMtvcWRiZawKhjjBdwLVBpB08XIeTqQ+alruVjNz+JOzW1HhN+8c9zom05NJQ
orAo03nNo3bRmuQN2PU/WPyeid/ZwO7e5mhx0A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u7E/rN5D1GFcBL/ioIqi6P5knAa8cU27XVaS/U8f0yBAQOFrlClmKYa+DncXAPJZnuvc4Gq9jBXT
Idr7CFNZ/e9vg4dv0aO6Y0zTgadQ8HUSsArdwK8MY04f7fy2SfseT8+XNHkW1kSGDZwSIzjYCjwR
xXo9jwaL0JsGmTtvtV8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
reo9LJmL7wj64QcopiSHUPgM4uNggSRLpwwvzVReIsBoJCYNr/NlfaqxUvis4tP+KhPC1QRdkrwj
r15y2slQ2ZO369PuT6+90SpEPdkxgzHOZwaazp27c6QMo5k7sJQccQdcVvZpUdBGySRU/p11eZzC
olCLUtUYbJWprdBPk8uSDowOZpdZe+qeA/SgoNOe4N1jwhPtz2HqWpCQIsNSDzcZlF73I/XklOwN
gBCF+gkGr0FLJLfquE85yVHRAGMjN40WmmSVOZyoVvs4+zUTBYCpXTlyTWk+NpPyxi5RvSfGVdrm
pnVyd7wVcixjZbX0mEnhvWxG8/2r81YBTv0b+w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33952)
`protect data_block
Sgf1Cw/cqLagInEQdE1It2yD6NHg+sjJnEtQ2aG7lwpbTt2vr7zsSjbB0+lcokHGcFxbJl7DGpCa
deyl2jZ7vm6WMw+YVrGw/jfCl9PRxZ8m0A0mFQpqCq0PtqB04MlP1/ZMlUYSyEPRCpqY6kmPFLXF
/px1BAAhcNVnvTXf9j262M7LLFhuH8kXhcwdQ51+xK9dlVybSSjSGLTmNQttev6hE/Fx3KMfWAWw
65qS+QbGbrixcl5TwyzMKo32LN/f/f+eMolN0CrB9u3xss/Gb+7d81rIYX2BgB5/h2HNsD4C0Uav
8YswfvqEBWenyx6ePQTvdCEbDbdOM17LhtpP+IZIhuIUpIADFiBI93HGHmMP5qjCTPc7pWRI8bjk
hPsO3K9m7F4XK311BSzsx4V5IyjpaTo69oJP2GPbm0nXPPB62UvamKo9qMFVAWYZyIKu++kilz5b
E6Vm1rteypTSOeIzcyo98jrkpuxFXQs/EE+Q1WxAjVH9qoXZ+RePcdji/rlz832zPlZbmReqD4zY
gVMPQWh9PPPL8/rVrnZncrMHLg2s/S1f15saodDXTEfwC6Vrn42CLwmbR5gK6hsJJZ1mAlR7JEz2
7EFTjCBOsig5HKKMjqYSCaCpF5FCwzttKBqvXC0lbgrOv7jz0V6CmMjK/k8SSLWdsoVjcXf5d9rn
IzHVtz/L0Uymd3t6zckFuXLRqJFw2pX8TQkcLbkMC28KYWckjfrVOLnJOMQFmM59vyHgd0xlfa5B
ubyhMdrxJQwvvLeAipEkkHEMAsBelD9PEPjH5ZsDI4UZhXWcYpg85nDeXU+nfHhxszVCjOzvBLz1
f4xyIGds6oaHglC43Gx0CcAtwUB7ilU1ZcMxiRtjGVforInMLWgr1WZqBZgJChtjQbiDD7mvQriy
lyiklq1Wf/hMknT5bymdDvL6/1jeO/Vl5i/j/SlTT9mZAwxS6BDXQ1Yb/yL76oFavFWP5Lrils/g
0Ypm/Yq1EM67tEvVIe3iCQGSAoS+IDiB+VP31dI0F6ZXYO51yqeknpU0i2551bJnUNMpU/A/80dm
RHI0Sh7s6JqiP+P+rJMmDO2O4z2pjPb3bdVbOkTbClDccBCHxp9/NdFtetaWs93d0XRUSmR+w6OG
4ox9H8INNcB0VyA8TQ94locDjO3Xw9YqvBAVr9hEvi6c1MFwiYEYR5XJ4Oxy5izSNTbZHf1KWUGN
zcfUwTim6/R/68MUl5A1nTTbtO+j2/fyldpbaVHOSGCGtXSnRy/73UFL1fNzcJGOqifAiXp8HS/g
p3hwCiYv15pnx2P+tJ1FTblS86HXf3JCNkjCOEp+jh5BJjj8OtR8sgf8G3rW3/yLb9z+niaIVPrv
RtBN9sQz0oexCLQalZMBk0UwVi7yl6xgjEaMy+SwMHp8+Oa43nH1z7xSjZhE3Yt5GUzKP0dTQ638
yKr+redF6fjIAWPeERr948LyBI0Rbt2qU9CWcDLW2JxODsa0ONIIg6cDDoxeug5kalQZnKsf7iPU
zQuiCvVJs3HZzAmMU/d2CN4fVr4tea9lIDgaq12puNYOzwPjNIjOygi8aybnahgVR7ZLGukDW5pS
OBGIPhN2Ef0IV442Yg7FJIlk0wvySdYHKdCS3ItpH+KJqrbdc9U3q73a0zfUskMF2mWBlw2j27le
RYzSa/KNDqcKlUMZV0aSzrQ9MULlECnno108FUQk0J6SDgtDf1fPE0XfJdHARopJTvcsFg1Ya0cK
JSIpq+8tgsoiiPi6zot6+nl7Ayge/4ehf1P73jyL3k4zVlWUJo7hgJBwV99VHUTcwd3XGqOY9gzW
NIQJAuQWaKVPXhS3fshEIOD8dgZzNShLCqkbwS5EKLq0gUZf4/h1k99b7yVTd4LMtKqJXgi72ihB
5SjFVlaFD+KjFBGv9mkzKBeh7VA/tjV+080gkqBKPML8qt7PZFoI1hYjGpHb2oabHKnkuYDDMGWM
lDnonz9rETEDyCAfrYxRdb7RShH3AjlI4mfoeGQX4mSb4md0GcoNlhCUKlVh+VJlNXohA1NmRzbe
3sBbKgsud51JzbfFidWp8oj1UKbi5JzkfMPUjBqXx4QL6V2P0yXDad9ko8xYafZCaVxqBsEsyJe9
L+As1LmLfVeeaO4THzZvvsAjxfYuHJW4Ztp4OI3h//vI8FcoHsyZ2WOHmcuiB73GwEHfkG63RkAe
xAmgNd5RbNaH6GWllHzS+SGurYTiqrY2BNfV3THwRz8s45RKR1SUtVjUkYtrsr5VdCooXo4V2Spj
Z6+jYnaVrBgq/A08Tj0L/d/fq41ASFUWyEeqG0lmC6c12HYsQFms6e5iQjUED/gseezhBSghccZo
D1FJA1cDaL+/1c5IytXThy9EkD2bpxmPIt2ldGdYlMtPpkFgjDCrr9yHTBkcd6w569WvxQmBHAnm
CH6gQf047DOos/EvxqP5PVWnbfO9mG+K36EkCQmzKSi+77PNrKrcxNf0bsZypdyLckftWTHhZ812
AU7/1zVRDlKUH6Ejw837g1MMLVm7977UpU5WHJ8702+MqGsxV9Uw+Y/fysYM9x7MpdzcW/GdTv8Y
M2Lve5B8Qlub+IQXs+26VCqZ0vKqQoc5rD0zKNIkPIh4CpZI+IHBtalJLgD4LRHyXZ7egssffPS7
NVU61CjP8D7NoRUnoql1+bPAw6R9G/IMaLtLos5yPyaF1PGMG1vZ2cezdUsKJcj+QQIQK7PC24T8
sEKJxJWqHx1aqllr9Lad6HPfiyrdZfQCfmWKhUGBE+k4u7fbQ5E9j/jIkmb8ghrSiBegIpXQs9Tn
KB9iRvFicM1MrbBHq9vIY987QZj0AU/lCq7kwMn/X52m2xPQs+aZyByyCbaGhW9ou/+OUlR/Gb2S
55PgPi0+YKDSm/0swXK3l2i/8lGad5Ddl+WySX6Ua/FTd1omlH3SCw/St7Cc0DCq2ti1K9sXfRqx
3vLT8tfDM4szN27FhDxUKfxBKvTczTjQADOAUAQtZ6iKWePxjll0LT9DUtD5jiHR5x14QDoYqye/
dwEBqyPCsH87ZYcG9j/MOL44s6lGGrNMnMOQSFmuunMiGgdDnMhPhAa5E7krISSPnfO28axnhGYH
VqfH7FHB1NOg9cj/ZzHHn79ykdzj/8SWBI+7qHMwbrnzWnbiCitwBB8r/jAum0BaHev7LDjOkznG
6E5jQ50XzTh95u+y3JSV5gaJa6gTnuxew705MaIoQXSKpLNSQbIgXOswvVqHSq0oaPCihjA+XbKn
OeIn0YZ2ulVRQdj3FkLklVA1BSCXXvNO1rHC7temGO7+TEEBTRraSp1a5+B3dRvgG+5jA013Tbzi
89mRMpThIzmpo30eRVNtZnGWX1vj6J6QRmE4ATEGYC3/F6erHVR8zNQA9NeKK8NDh4dcfrJW4+gW
8ZwVmw2p64N6Lol4WJLQK3BB+6YEaMqKGrdkr89kVWmrkfE7ihNHwOl78vsVcFYLiB43KShmqx3S
vC/vR/AiLI6PaV4kAafCrBtJytzI5uMA3EPJyvQvjQga/05Q8O3C/TVqa5/rOQm/0b2N+8Om2Sm6
aA7vFuOsLmxxdXndwNXAmFX4b5rIsCNQRGI5gF8vQHEvqVcyTyBsgMydDnPTA7Eg8BeAV2vEhMEG
ceTNUh+dA9vSyzPbtAgVwaPoGdpIASV8RZKIdWEHzt9OOv5avzYcLvuELExphhF35rMHULdbFiX8
uNhT/PK0ZpJTbFiMJNrM1UMi1CEYeHRfC2tmvKP9cV1Q8TF9znxuy0D2SWwoEXkXsdsavMZM2ril
uwnkUv2YkGtc1YE7sVcN+zxSVQcgJaxkEuOXsRTi2P9glVIYly5Zst9E23+zQ96t4gB6/yAdkBWE
ATehTEC2gaavHYheb1OLFGJqlUBgmLBpjY82tFWgV9UcceWI6Ry29FTVOgSc/Y2UiuJmj4+zzlXZ
sIesH/xVtQaqsAnUDO0SDfw8traAOTTKXJ4zjR6NtY7NxaWpNTAZ/vBXgHxYKgnxN0sVBizwZB1H
hOLNDDu8NTzYfii3YFEqAVqTWoLisonCb2U7uO0tN31jwQVHq7VpKk3gilF7CaJrwu51zedGI3hx
5g3mCpcnwQndRS2d4ZzWiHRpzfgNOICNfCy4a+HynM3ODdxI3+UYtt2nOq376OT6SGKgbduD7PuD
eOZYJTYnv9hZVESB8f0ikWXfDC2rv39BwM+++upYMos4W4n5zefAN9boatUx3IYhYYp/cXupGHrx
WXwbPfZ3UeFNMf7qtEt5Cw/AcEzwa4tP+oyciQQS7RB9SL7NM4n2S2ILROvcCJ3Y6iWbiDiH1W+Z
kCl2j4V1kOf2I/QyUMqwPkSQek7y7HcTIW7XLLkvIxR30orh3Fn1T+/gGhAXxstrqLa9GLJKy5rI
4aarULMny08Yi3MFa+cgpJs18YCUxHqwEq+pIdk+tqXfGOJxa0ecde8gcwPFS7wnUJFD9CMJoLoB
yad8wDUtQ5aqQmkVEU3mcqEAoIx8Z/QaQGNEMclbdgFydHAJJlqSa5D+++Pi+OBqOlyt8pn58Fkv
83khVp6FjNozFrzOPJ53J0CW1s8vhOPqf379cpYWhIeBJtKvhZ/ElO2RfTH1NiDL3X9ClQvZLdRW
jbdea/CafkSumF7VT4uc9hwpcXX/0lJiF0m3uZmtd4B3vEqjeyWe4mcL8uf+TNUvQ9tcYBvdOqr0
409bSpb9gwodTN3me0d1UTQMi9zp1RC3HluHbpbSIrmyLso54XEIEOcZvgTW2D3Ojl/hymmay3Qp
1GrmO4Vv6CYe1wS14YV++zOGK2XRi2ulYNWgKWLs8c8M8T1mRe6S7EzpoXpbWJjLOI45Apx74uXp
hI2pP1wDKvOs+TJJmorXSvDlODLQf33alAYVEjyAlPSoYb6VuG1LeuzF2oMLh0HcVvb5Pi8+pO6X
GJwoVKyFV15fSmb5gpFIRhV6RCh5ZZhI1hAlTBaK7os+eykzZWrIV2L8HcXGLn32C+XjFZ06wElO
ooklvKGVj+4wxvYv8GKq1Yqc4g+lbuRfFZrCFNCmuwaQcvsiVIZaG02ATZ6M8YKNer4h63IGDIyI
SwAkg5T2z5TkDWioYw4OanCeA8Mz5W6xorK27rpH/9daABzt86J2Ce8vQJ0f+2Ndzbfo4yLQEqwj
uYg88ErkoHAN/YGa5LC4TlAdgIHDJ11FAKJRDquJQkmhW8iHh+h7qSGOJ20P2M5hwCIGDY11A/Z5
ew8G88Kr3sSGNEVi1jQAEhW3oKGFbcpVJXrlKWo4hNoUcTnyWQNkzRLFn94jhlxe1S++OW4Qk9D1
vuu995lTgIbjUxo1Dyu6tMP9GqCgbnPiqob5Zs0Rsze5ZHvgwwHVn4/GKWrGWbjU3f3VzFX2MVYz
eQNHXPi6BhQrrm9zzHOAbV9fnQfIG/9tG0XyJD3Snc/NnFAhWRsr280YX5pZ+hywoCnYYEBi5fFF
8i4XhItJ06wzYqujhzgaAhTyop/MlE+OwUmBCToaPP53LxeVpjWgkY13cnouQ/zEnSf1EJimefFr
YXSvl8hKhri7g3xJkzu4bHmEESzrRCi+DEKPMdB23Zn7wuhqY7Zb4eUvCduG8R4vlBryy8z38V0j
IJ3F7fHCutqtealONniH2uJjA75fT834BU1bPmXyilmroLcs6qjQ1Beg/OW573uVzdVgPByrOmlb
+pu1pcfwRFCwFg728snHg9hf4z6e1WyrbkMWu0rYlwYvI83YVm1i50aFJjfQyUHkzDEp69Ildsk3
K5uH8shVC8/BZ+VT6I8jNvO9Bj99nr80RzxYbPHn6D1AFYm4ghQCCaMR8rDd7nlVSDEMuk0Bm4WW
7rmNnjzpLsboFXx3+EwPFa7PKS1RQfWJh/XUYqwSNwN+Uxy4RvWpFs6Q7kvKRTJK900pjdA4PkJM
3SUR4f+CZDb/Jhgkr1+dk0rBEmBaupW6XMw/DnsfTs82cpzxNXtQsHbnTKK0fGrCiiMFPlTG0SD9
FbZ4zp1AEy1TvoZ9sQYbW2JqbimlDv/26h7dJnEv4DWCSVRwoX4Gg7774/lS3nD5SOPiwS0mDnsA
+3DyyvFtSeNHTLePfhrNCdmFl7bCpun/iOI0YDdrfCfvHxn9FQPBdyJU+npDqURzJGfePWWexZTm
jgd59wFhQacb3C6BYQJ8KZJdccysH65VORSvk+QAY67A4max+LShITxWPRvdwn9mFW1Mt21f95aJ
xO/I3tdIowyME3MqKg2UqZbGIgO5+jPc7HL1Q7spcTivN456wKIdCcg233OySjb7dlAuiLU2Hdpw
9XDwAkyRSNKdzFZ2qn/EK9dluZbxBnPl/pBOpf9RN4unUxv7uDMybUciL/lNtSqPqRyimAT23Qam
1DQr0Tlpf9NoT/bsZDnAg6LOhrSeT2YzYXH+dLzI0oNtJCJlprTY4mVoLhLSCLUaxIncMKPO8B7c
+XsuGWPOdpJgu1yG7MF//I5AHpudalmKvyGrs7H2rMU43qWzDc6fBbIHN9NCn3S+bWmXk5L/QW+s
FEmfNLShyurP/ebg1br6VhQG2h8f6vRfqbsC5qYri86eWCkpcLzWuWkOt29mQxckC6RqRQUMNdHe
c8oIgMji3v06yISdDxlY5/ef9/ZzSm242i3+RHYZ6grk+Mqs7VOrXUT+c35QxVq6uWSAEPukr97s
RwEYKcNdClAakBfHxncptZALVSHsx775I7nyo2OjsnWSubTSM3FU+5Ay6wPE4I7dYUTtS6p0tPLd
aIIErEBeoVGTaMRcNio64lL23ktatm4oA2Y9CkkNWnC+O0lUef0BzqCIdxOQ5h295ldLR0RZSALN
gRfLKp+IxhRU4S81Hu9SuLPOZWnjo3lanATyz4nlrdkFn1IxN56g1G+tlYUinhWababVrO8bo2Qx
SbB6nME8oZIsFp9zTepfwZsIxYTSoudkVGx1u6bAxRdwvsHHRbNCB2jmpFCLAl7toe2enPLISdTs
EOIRZjrNTBvtaRRMVP5I7jMvlW+lqz/xIIsmQ3AJ6qwUJs8nDAhRzX3HJyKy/HBxPI0SuKMBp8GW
zskrPA77Y9Wx5Xw1JyYlb9nBYjU8cIcfuGxa7NHCLGNd13jEhkfai79J967Iv5BgG6Hv45RvB0Dj
ufR58HPBJwCoTkQCzpFLt1q/nG9uJ5qnmugMt6ymTCri7+KuItyZa/CGEu97BDtjHz0SZkpkRZGL
8Mfwv1OeXippv2yCSTr65vHOC+6uJ8Hq4BvA9ZwJ0CYN+3mdhS8Dm8t+Yc75QYUVmpp17AH4o58k
9paDPbv2Xj+dK0puZJkCa7T4TmUP21Pn97ttkPODzHpe4Hz/n96lo7PNP/2EFNR8ZoEZzFPEOofP
L6FSjwl9X6FmxKmLmG6ZU0fvU+XMxgjeUPuIfg+B1a7551x7x2SOyYvS2sTLP24P+cax4GW+BZTL
NQtfQGTI+fD5q1pwnQH4INc2Cfhw1PMTJLnJ+WaGWcr5+kENxU89dcpdWdUT7mREMUWXrJjIn6i8
CryRD8N34IQrRgJmKkHexI5KMNhuaUDYgekS2mcF3v5wC2/1zMTyfSRqEDgUEOhwMQKVOTY4oST0
6mVabNqiySzcfidgpDTJS2DTLh3O8bf4yq+Ey/XW+88OVl/18u+mloRROlVUCbAyQ4jBCx9Hi2+R
AGVYbuDfW933agk7MqKw/ZV9Q35xqd8gtp8BSD/hDClIsdDk1u0GF9ar7xjVrTBY8YwxcxqsqNSP
21VrhjH8jgQj+ASYVvjLm7zTWnT90maOSHd3oqhEnyJcv3GQKbVdaLiw2guITjtHbcQqACYNZZyE
B03+g7YF3PIhHJyt3jaOKKzg1FqVmIfD3bkH4eo+rlQCy3xIDSSnvbDguNADzXQ134T03z2GHnjx
BPxgX0HALZjPy7VmY4uLvPQ8uP3O0FC6nf3qCkcB7JlQricGkldVPhPrH+U/tEsqE5PYujSKofpf
u9hZmFetk3WiNclLbioqpXKG9qVhvMC4qJSI/D1zmYO5OEq8FU143SMlQvbaOSU62PUwt1Xd3eT6
FlddZLukjNTgcuWQHc14InviC5ZXO+NaK7KOBFxLYBa373//C+c8mtBhscB/fEHNKW/0IOCcLW1n
Mw8zLioRsxYMRaYcq72wIydIYFtV0PyFZlbDl+PaeKEVw0iEUPQFUc8Zj9X9Nzm2GgqJX5BLllv7
pzSAnjh2dA0liAFZ9K6s9H1uH/y3jh9FU4fyuFhLkGumvjZrskfCqup1bvrvGUEkMNi/v/uIFvPs
Q2ENLZud0YCggSOLyFU41tFUIweau8oSZofYJFE7SKl8E8ZlAWIC0EZU4pGqDO1+hGSsW7QrxQml
hPistLUYXYbLIce/Czo8W3Q5X3P7J4ncZApPTO2n6DZJC2tlQSvsEQB4rhd7oUH9/c+XEbmSyoqS
EWKp0ipi+DvnRVR7ESFC8rHczdP6gQKXiNxgLYclSv8AV0ENGhMV9vMAWX5iYJuS7wrMt1AE3o5B
2IVMBDJx+5wYVoLM1AmNj99YBwA2ZNx1pwjgopDRdfCgGIt63Q7t4P6j/mM9wwCnGq8weQPGwIZR
ij9i3l9jRT5DD4nDd6QWJAyFwYId0WJv0Z3KmwuV+uAyslL5NsvmmlTP12tA+kFbWcS0yd+G1K3v
xVbjtQ7XAUYOdg+qER+/yxuvksTnsFyrCXaeyFkuaNEpEhEdi8qUMkDuM/eQ7FW+JbNJYCeLBlj+
4T3Xz+N+I7/PSVynB56u8s7/5/ch1x9vXjhkEd7nFBGff2uBfmZjQf0Zp6qAdFLJ3pfXHWR+HQqP
9CzyDkN/madU1XhFFKIQhRLFKNI3IMz1j4gQGgWTErU0rQD4yet1nB3cU+73j+cSOlGVEnQFL/nn
Jli/DS9jA2ZhhNEXZ2XJjIf+J4xeJIYWNOpf3WAKwy4A7rXDsicfKXad9tp2zhdf+lmot0tlq1SF
Jc4o9areulafOBmuJt1LcVLVuj6JPBsIlscxq71CaiT0PprENr6XNulLNcmND9LqDBQmDkOjpq82
kG5TIUpmdO2kFP/+EE4o79qCVSa3hSuSBzEO4+eHkGRugAcS0Ptz6pcncRfupjqkJ2yeqdIP1/Vj
AwS6Vkn3ctbsJzK0j9iz2caEKn7vQXIIHu4pcojG6fvplskQ03oJMMMffihk1Uwe10FWGfaAzhFk
0Vm7NsXVBxG7rvXFm3XuIoU2D/cNeug/FxzxUNjwpkLJ3UNA/14qDokDHkShoDm1E97QgN8Kh+Mn
t8NEPNRIM2TBih+oNPfUChfvz6DSKtrOhYyAzJjE8yyVD+kwexvucCCI4ueoQ5LerG7VWT67WblK
EDI1qhTS3pKZbEZhK+36Ti/P/5AIMSXovKWngYvZXmVchUUvX7/QVkzJjImUZYn6TdKkHHyMGYNe
LOnitJ5WUIDzyLvsqe4Wojlve/IqGjivuHewOBopgTmid/kZdRM6xqHc+UpCkBwYNJscXA2wCY8f
XXbga+dDM/hsu/vNCl3+XoYMX+BPlO97omWdRFngWlk6p0Lv7CcVyKuchl69vR4d3Y/ztwTVJxSJ
vRfMnnzPXyrRtw8Tq1Abw4EuR4TFgmwsfkeKogoWAipYiTqP9c436vjH1dJU8uS5ilPQeAbg1We8
boTAL+PW7ils32iE35ymEjePOFMdG4MgmUB+Gg2zMLbNYSEakwbHjAiJ7vn+ZRKdfjl6O39jBE3q
AzAx03c1XKQJaLY531vnvETOMvsC3avPmO6BTHs7m0OewUcxAlRw2XlLL9cYbZhsLINFgyY06FTt
Ro3KR6c6Yy0RVU93Rq1UzirbgPi6vVa95iDtpx2yJ5cSB/B6NqnSXOp6Db6YbUlvgkmm/lFFjfgH
wDQfCwExKUE4M1MnU8UnZvYe31d3HjNy2nOSG43P0ZdxroWlrtqkwah5wJ5JBff9BxzpVfIwNFJB
j9p3gPAcXk4AEj/CqhC4z9ABfjjlqUKbRpNBOPUP4NPDd9q1qAwnJ7v0MLpVbTP/aUyYPcuImavf
vqAuMcL3ZGb8lHWg+D20x6xcUnpHI6s3usH2AD0chmzHlC33irbZoZbfJBQ8nxk7gpCAEikJijS8
feitRs2CNV9WHnxjLY+PHd2dut/5ToRGqSh9ZsN/WLTX5j/kKyjynlMC6IT57/VvPIQnvEy9mmtI
+obiHiJRmVH3mGFIixxJ/9Y8YgrSAygqfyta2xXl3uvWX2bewAhqT8DNAjG6+8GWWKyUlT/Ic0Ep
p4EUBpydeSAWOVBBSL99rmGunwnHhS1vVrhkjroO9Q/i/NMYgM0rJ8G1n/yoqKT5psMaOEvW1l4x
3i6GM5DDzT9IjUntGLVQmDdwWcAFi11uuJ8GFONmY/V5gcYu/xsy+0fx6pN5oxhL2+nYr5CrV2HJ
zqb8fQk1r32Icg04i853tOeZCjjLblppX03pRfy8kXzOKMIitz5t6GgaieNX+qwjHFTCsFhoohMX
BsjHCalLAAZtFVOfwSI7wpkQAUbtlktLEAOl5QJmatL0VUtxPcrZYJfbpLpaNl2GObAgcsYMvO6/
iwrEC+3/HGZoWFb94aFicG1X1K16odtwjRJxdB4Kz/sh81VqWZMZrP9s62EvTWUDE0ggkm+YYBJQ
2Haclfv3N8sYwVeRvVhK1ksUAnkP0a7zfiIwncj4LVXQzzfKp9DOIX4qEbGkXfL5M+x73hlwJDrk
ZqBC197czbFaw3xrBsn7QI6ydmaFeHWidqHLUgBn98lN2Bojmv4SIGKuM/L8avzBEGEeRB7QbokS
WeJ7UhyI2+w09UtFqz8tXChQubUZH5evr0R3D4Q7ZtwnhF0OLcVJTnSNDOqkCynMGJsO1INS1HBW
MOMTXRaJCafKpxRHFJUwAld/LbdbVDa/ynG4b512y/yvVz5bQtQqhkD3fuRDP/1+s+bmXmRA5l9F
7+qVUN7I6MKNNnBDFb42TOuliTAx2D+BH+O10/7txcOzrOcdKeZRZd7rpu24x24MbPnd5o/zt3gO
Ijxncr9o5tQ+xGFscICnskryoGC8nNN/Bfl1UtO/0YprZIeqgJr1sZPxD1bVCjX5LQlhK+hqXOhH
34ABJXGAYr3gt3puWAAQKik9ZrNzgEohNSoFgBTmDp8PVRXJyTLszzruWiFSRz460pc6jgJj7JIr
Efud+MS6otSFbDu4ujfgAHIwM0bgM679XBrBgzzuzeQPvJtVLh/ES7tebqIkWrIDobg1LBXFn13n
BdhdJkgx8+jfgjiBfvahaUp+BMxKLXGvf4sq1gHg6oDt/XGsVeAdQcH/7hHOHWM1JbrOpyOKzQEW
7g1+kJSrcOK86juzPCQ2jNzZkql1s3I1MZtJCFsLWYyDlTJ2JFxRGnFjVgN+VbxoXfoFfxtJgs2I
5VdpEn4TdwjrPOXE5z8y6eASFzWCM0V0X548rCGWh23lUT/mva8GA50xuNrTmvXrixWmB5gMy2lN
+1dNsbdtKBcPmgLPmmWZ9VM6l2uhe9z/pUt5KMdoiy8pr0MMQnZtpO5EIxdH3U9ZFywrNfgaKDVM
Sa85uSf05UakytCUkXCh9y8txej5up25pguvJ+qgNyus11vZxHbMcf1UG3b8SOb91eA0mCc0Dmsm
1oftJhuDOp9Xrd0+QK/JHO70lDvGln6La7Y+iYEGQe6JA6p9+0RuLR5NirmpIpoMHs3G2F4Dtpjb
M8wJr7lbPt4KL2K5Xq+2uxkFYygzOof9nbxbIAzUnFKdIQrnglDDDyP736Ee484Ah9GuSDNSuVg8
SV2XF4Kg8fgKw4Qbww97iLcjMeLjIgT2yGWbeLLS+mCvm7dKKiahIDwiNaU4ffXo/xspiysasbJA
d56a6Rx7qJEAMPt0EXUuFt2a+Hkj7vLrvPx8QHhiNNWchT1Ljk2jneVQaPDyknyjtztOwaRF8xU9
argCJ7pSjKkWpYwhRD7JasfOGdM255owE12Z/W7WomeK0O3A5UAf7CdVdnGVuqvopCMT9vaWm93U
jmMcIH7Jd7rl0yolAXTaLL1lhfrgcyYnquf2NuPAeRBCWfAaCQptx+WNthwrwGn4/vlnbKrsLBHi
6QMwzFF54SsQGLvN0HDB/pOWV8fL5Vg4rqAwMRQgQXISHEvdSFBjd36KadiGbhYHREczX2UbU/zi
NftachUr+IqoQ50z7xznW9ThlfRWcbQYW+XKI2hiSrBJuHNpXRdJ03FdhdSVVsEhHTMXANbiv5W9
cSFAecvtxooIGs1QWf3rPlSjTt0ao/JXAQ2c3UY5WUCGxvWEq1ZUk61KtE6iS0W4yxguc2FioLAM
uh5Awy3jnimlwK+R7oeO/9+4p/wcLa/Ni7VC7R8aN0Hx2fOlWhmpton8EtjTMVH2l07wREHqSAlp
rIw0fiAtAHrXpulj+OCoOxT1NyXUa5WzPoUKJRO6LKXZ/6S6I0LT2JAMOmUeF4LQ+lZ5NDJ/W8mE
LzGR1EdrikS4hclydxrtUv/ajHn48qT1OIt0T0PUJKwyQdlUDnRMwEuxqN3CPw1L7e/riX9j8+LF
jcbbbL4DHcfnjt+2BWNckguQzYmUJfsU6Wb2dS7ox9JA+ENPpjTlPaYpI2934cCFlj0c9rDR69r/
/cfea3zMTLYkNH52k71UCa2LpJ3IL8uT1ffqPCJgeRtLP+0UayTrSHBCJT+IZlZ7d5r//395ZZiG
UawTIEgnGYt/OqNvZUPh2RFOeKXx4AtEObJLToyBSyXT2Qmsa1atRIzXbU0BAyXsqmpXHmATKTDL
8aJQKw3c2lBSHb2qakScnDNBRLL2JSAhhxpDMke7khG/EMicSwjDIi/yw08sO0khOrvx+DJjxcmO
9PZRmyyxAcuBvy/GjRCkoPovMYWZf+V32eXutvb6Gdjf3VVRrhD7/vZmxZDTFZamyKIG602vk2/W
RehWFG61FO6v5q/u+y7RTL7cHTHIwpm9GW0xxxlq65n0RuiWH7ddzrEErLJzUWScUn8oLhvKAwpU
ptFLmLJCuyPM4p1+sDiBlyOZYNANGQF4dRQSubvQbphNL7xrmHSOJ/ZMwAiHNkj//JmtG/Q7OUo4
NbRQCE0FU0+Q0P90DxMo+HTSxdbP7muQjXFZoXj7Iz7bD0eoS5M4Dppg4jh55RO1QVl6XEpBvrc3
jcotSkJl9GNZtSJHy2KxUPGIKfkk+8DkonzYNuMxMKNM5+fO2WMhEL4emwfJSf7WRWivpmH772L+
zA3n+n1bmdXqhRaUGjm+k8M+LBVp4qKIf0PuzBzzUZkAEc1Jkn68ZDEGFrGUp3FgcUpPq85aiHDM
43PEv67+aQAtTRKu93eA3gIYoK7zUiH4uzlBQvajImpMCRoHQ9M7QAK82VDh3X1x87x/WCJOr7Hy
M9Snp5Z4xA9Mkcbh2pKbhD4RKwil269aBmdn0UuLkNYwLN6Nw5ZYUHQNORqHbaR5LXYYs5/e0Om2
cZwinCxM3jhZpetMyZnde94jB1iU6U/ttQVbt2rzmoAfAPlbypkyZxxzQY3+42+L65E7T2hb7Dzt
tFj769/336BzkfWbvbz7Mb3Rzi/tCY7zp+bcxjxi/AQf9r0ym7EdwbLJ/vzz+MrD0hZjxsrG0L4V
Rd0zEzlI+GpzdttP5KoenkxWfwi85Rp0FKg3gzoIczgSOIzVGDalFbR45ulPyTF9sKSzeiN4sEK5
WB1X/tNO9hcw3TmYw1im/d/9MzpbOJctqmaO1684Ncv0JA9HUWVWYbTakW7SxvSeEC1o2ZaYeedH
tfzbiGfJVbmi7nLwlyAoxDCn8nBb/KydcoStTuYGk3q/X2bwBDqLAUPVAWO8PAj+dkskCkv34PhN
duKlDlNFbi3EFXWj08Qm/6AcRg53y43XpYcVa6ktAhCKqyk4fzeQnLnjQlNxP0IdRq+bCkAlfXm7
EdtvVSQIPuhiL1yple6yNAd8IYW5VxAtVskAGZgv+YDFtloGnUKfp705UxQ84ogf252XCt0r16VL
+15ndinRU7kBWLXSujVGsPv6ZDmwDwbjoiGHzj5nZEEq3Ez3ji6A7db1bsToVoyPr+B/VzaAqGKc
9QlFu9Ndhz/wsSE0ImXPk7j5Iee80JdGJk4kdd6TOpeX/q6Nsv6fKJpcno8kI7+mWAN/haOGydkq
aP3fxRREmzyhgUJ06v86crNIy+gMnxL1ukJigIVbAvriB8Hp6dK45QUfC1p4kCNfeFPwZyGo/F7T
a64ZTHGcn86oz7ZhC/C84R/YrazBo6bAvjOnQeN8LCf6G4qTwGt2yrd8qISmR/OQ9f0Ro1orJoKw
IqRuQyAgYeXT/ZBm2DI7GmfJ9Q0wVWzJ0XZLXjboZph9x2TQRzh18EY7oqD33o9PczZbK55pn4iY
7wRTCm9/QX1PeV1znEJIru2BCb2fkTm5GT4H3hYpEIj5Q6XMb7DvB3QuuchOj/+SvHDAgQihFMRd
/P9mf1wUuL3qgDzv6NY5nexMPjTCHCovwrrvhK+L34Qf9hvu64urIrE04hVe4q/nWdMgsywlujcg
kcez2z4CI+n8cVq7b8mgOxC1eGH4I1EnGDVg3fe8VjNSiZp/6JYko/tfrR3c/ZZOtnvvty1Ua8Gx
NuA2Vgkc93BSSJ9O5ryAldYmABEaO+w56Y+I+4/PzLkeWnJJkRmgIF0MuobAJ+RP6HevTarlTHPh
noiurt2RF+SePKQgRmYXFOyJ5Ci2m2TQ0EfyN1aD2gHJEKAef/M/Ow4kyrSmn3va/RES6+Cdq+Pc
OJJtpgM7f41nuuCtiVp8HmzN9hVpaUGDKDH90LneEx9jU5COJff/m933IOmbSkC9MgH9erSSX6Pn
N0DYXO0gGX/Xe0ganMpPbdDYsc4O/2yBHvmVlxd9j8gnYkLGMk6iuXNf/2Kehqgt3n5SPAJ/7X08
o9evcRSV7tdnxyZZ6+SsVEnTFby+5DJCwSpJenP7UrLiKQPC0bB6x/ElBp9Wf8EVzmXxO+XDKSYf
oRdE/jvke46kPN8MAjRpR+y7A98KyLzipkc/AeaeqxV+x2sM6xKJUB6yc2dpR3KW9Z+NfTtqRAfk
Wz7XcLNsjF1U5jW9bn6ZuWE8uyQMrfdLh6bBX2ojEF7FSHNaYw3gyKdLdDI00snp7w+pNmP23XaF
lwHvzNGLOrU2SNXaxFqC37E2/PcqIfVWBlY+War127lt2y1Okm260WpYBgl999PRzqHWMtXqkZsI
DRFRkukQVFGkRxMA9N00Qx52HtOxxcUfn2HU1477edRKCp3imc8NGE+V8/TZZRN6CRtOy2QZQlda
LA6ATI/yd+gNuGfNBuNFcmdAqkPOvzFlUUJpmFPlXqYD+ZFD5eof6mWmD3B98VHMrnu/MtwXU0MP
LemD+JNbEcGmrhtgsJrz5/19SL4Tm+Eca6e8xDTCCePmrscjc+sskVwrXHjZlQzJgKuE1P2UfEyE
L7UoiKzQgrfxmq9YyEOHUXZ5QicYpA1mj/L/4P76T3JzlqWRQSC2jILuQT8cK8h0L38z4RaL/mXM
MTRFXEMeBQECV4Tuickj5SMs+rKHR9K3JhGtEekDk3FPXlz2FLiYQ941WE5CYqj/Eb59zJmWResi
GHZG+ZWIroLwRwq9ds2/YqB32p8a9IXKawOnc8iJA8hkfubYYqHSxwLhaXhxx/AameoptxKS2zZz
L7DJo7961qkv5BuGU0LMQGD1f+PZCFiqFS7jelk9iY2IRMX5A9b14Ure5DGszlR3stUeKWxuLkiX
2Z6eFKfUPy/uiQKaZUs7TaW7wBMvLpXPmapldpTC0uT13zp8DA4oaUrLAFZvE8wRf5VIJnvLVvId
/5XfRCl+nmfr5BngvCIAPyH9LTm3rznmLpiXRQb4dOlB6LJrkVuuUhp2TbR1a3dEcK5zcOExXVUn
swx2ZRNfi4tK9BaqvjZGx5mXM97N1iVh8qA3RjeG3/KS8e6kbxEsP8ijqHD3TRnWTVwGADTU6+go
B501vcP7BlxuZhiZl80ocNwt6vENBZcLtcM+UA95Xy1Uli8LE6HemMDeUSjyYCM8ixT7w2JZAeqp
qlx7YvXaiMYA2pYejU4v2iHWhWuh9uECa+hqT4CoMKIkjynTddVTSB6kBe6uJi4jj77vBlN4ai2b
hKcouj+u15+zOg37Zf1646vwVybRGDA0jraSDN5lVHeINU96zklCHXigJ3mAhE+gjHbpGgzwGo5O
KXDPyE8km8fu1+2KBYa/9ysigq8rmLdF7mF1nU1/dm9t3buS5IYwqIuHmCuBw35v5KltqjOq5AtA
iLw4VW2ww0RJWBK9IJ8L8+CxHS/UeLZL/sqIyt27G90+WOkFDarA9Z22TZDINfYn2owtwR8kqPJZ
Edg5Gn10P8OuNwoYHwgSMBhsNlF7dvyfCtPYDK/YFt7y2HnlPGPUDBSAf5jRjBr6zfo2pBSPFScR
O2NLUCpaODGJiaFnVOf2bBXbDenjSA0Se4ym+mNlpdRCJ50VR+zMnmvykvMGLJToIj7jVGc6Z9xx
NyfhFWd/EmpcfsCY/2zUmdQbNafT9jUJnBqhwcWvZC+0tZbptniJ4AviIWk2MK1Pd7KZDL1AaIHX
6Wr1Wxqf7RD9xyUBI9VF10FklhJsNA24gM/ORWB1rOxTEaRTvkjFlH14W0KL1mdCyN3he4L2BSqj
TAU1WIhfu0UKe61ULp94FWLw/IcyWEib6P5YtYKTA/qL8vb9e/Lwd+fvZ5lhfToePRPGnRIczulE
txbnUgxT1/hx7M3k4vcIPMNPC5+Z+6qGdC4zsv4dxZ0TKOOjdLLIv5ecviCzDJXFNzZ1qBb6wWY1
PPURL0O9SJH35TGJSm3LBjWHTCvDVUZLa0MfR0aLpoPZF+1/n+xvzP42363z1iFMbOfRp1JN/TpX
ZyB603I4APR6Ia4aGocs6nDphj1p3GepYTSLn07uykSwB9uImPiMtAVeCyxFeBgndU6UkjOnlUBJ
s4Ztqne74qtSBDdwiPzDIKgFO/44szyO1KeDlnaSrCIjgk73PBz/Zt8T+l9S2gyr6u/WMoYqP1jS
qJYZLItquDuA4Fr40Yn7yA2zgef2Gf1MihxRXuR0DWx1mc/X/GpQeS/ODNqVE0BtTevTLDtTT9Yl
nCHOP7zyge4CC2pKC1w5XE6vQZR8VQO1pdL5T1tWhwJb4iserejJ+8OsLrIEAee9DtVQiX6ECMNC
FbpvuqNUD28PzAUEcoiIZhEuxsPC1NuHv14l58YlURpsGSnXWvqPrjUHzaqyHWB8Zvgh/oVdNXLT
OfBDiUIUups88ujumNXU60AFwEK0CNhjeiNQV1FNUdGIsPjJyfHmOctosAobgqX24Q97Up4X76Y6
xBXqJ6A01BZkYUr9JB1XMc65QTqBgHxJL+zQ7gKyGi1MsgZhoEafzx/B+uvOUlGoYouCI7KWQ6DR
Yt8JIKgIsuX4Jt4fgx3ps/Q+JNPRGZjvuYFUJ0hxnj65h1m9MaYr2ROj4HNvksVUMTh+0xViAlTC
Mfppv0ee52lNZead8frDKiYQeDXtDzvc/hKQED3veB14QoAq4s/8RVwhRE2ptI+MKaVdNAXxu7JP
+ygw9mrQ4Cw/nvAV0a4YCpcGQhv3ZzvweztU2nwfNj0Pe3p1lNRQEoLgH4wMr0MWSLiPeqvlLzLf
wCfl+MYKCWSvafvY2EPi33DtRTB+v8TLnK/HWpAKmGC/XR/EUzaTSIKegYxNt+bAfoW/LPF7g7Mc
G7zJWULv5ZepHxkCvAOPpMzrSgRhHs2FjxXg0hmFFwW3/lAm2zKDPigCblSOJle1DBmeFgzHmUbQ
IOE+2lFrsELL70CY6QwP5g0+oPmLmG4I1MFqhAHsqV3R3wZe4q/t/vb8u5uatqG+s3NTbzeeNq/Z
W8b1IWrnlDvpf3SMGUhhO9DVWnGshCwqgvMOUEUKPND7pJw87EqAHStXxZUYtgoKBw1ZxKDA6vwE
zLr8CpBb2vIED3U/sfgl6MgbS3auGhKVh9EDOG8W+bhi/ek/Hi7dtcMABKLhGu3MxPPNWZ2cFqYs
VbE+kqF4+7G32jn8EoewwEI7RGyBfjFCAYExKmFfY6LJUj+2OnLgxItIFtFgq/yVLFMtxzSAmJKq
H+C0cCWaeUZsGtHQvbXpop9Jh3g5uRDvImSwmKMV/7d/KlfKN4ZpYbklj9s4Xw08uUiAxMdFKoT8
QRwDKMhyvBUm9Z+rPXyHPfmAE5E8KBwdT1GHqdB/uRFYefYDTZJJGDiA4iw7pK4k+OFnulxoJ4D2
HdmTT6UQsusoxVdiuNUdsn0h/+Zq6H60sy5gK9AiAEsunlxIIfOrTtcZxrShBE6vjXUlkO2PS7kF
7hkv2yDhe0rMjM563WE3ToPPCC1N+CHW5CVNlPnirfcvhw9rFs944xsIs5hGZLMxPT61FXxpbIC1
fB0nUUrh7hkm+QNGrlxell0UkENiAdYkOs/HVMZOqIPeb28B3IfvqD6D2keIKECXaaunUFyeTxuA
B3wpZdFYG+Wk7CJWjEyT6Ua/RIY5mfdputeQwpz8X1mctlv0I3G8ZZl0bf4Qs+Ug53NHkBi8vcuO
GKoCyeaEXJC06LBoONLcLy67RCJMAgCAIOcvVJrR0TvCZFXtTvMh9r9obLHVkDQ7YGtUixGUlkvs
o+PZt04mpL6OatIPjRDQ2iqxHfJDsIPtjbWQm/shXIcRBO/fDc0IiPQjV/hhSkPHTKpP/cfzv0IJ
EO9kwQ5NZdVhcCZHJsLfP5BFeiPH2xtaFCdVMzcNlrAtuF8nyWd/zo85aDh2LJD6R8tDbn4moHzJ
fZAtfI438JDEr8Mfb5vtWtrzchdyB0fN/bs192A1PzWA4c7HMVpxbeVq1QZLz3xM0rCfNbNBh/Pm
3+QbRWVkwpCJ6OeTzP/KuTKhhQa7QQw+Byt6q58ahbFqsD8OURF8A7O1tWHV8h1Kh0hiODmgUhXi
GWNwwmZoQCTU/Aqka0GtzLannP/3A2s72flNB/EGg6OGHv1QqnpIIrIj4FIAeO1q/XkR8PwqJij0
2RPn5cegIeKT5nRGgW16362p1kvjkAEfd9FPPuCjq6OoshcfvscijVKEjeAE9Z8NCuAucUGq6zZs
5wf8q5PaFsjf4lho1DyZjHHtYXyLV3b1khdPa95BVU64qaA9cSau7vHF9RItiA4b9N1hNjRhOqPS
jj/29xp0d7Kwftl+7nuj2hEtt5yn9SGs3XizS/RuIir4rkw/K+hbMTDeK3djntwcSl6OZNsq839+
+m2OKhqgvMPb+xyGgDH7bve2Wads0sERp3ZaMP2LtDwJ0dclmU5pABYScw+sbM9J6UbzYaSsOPxI
ww8TRZcc+XGV4T9B27iY/iEcnRmcjjMeSUaPzto9R+tzI1bELsxsCDbXMxlXY1Uc25UYR1lkcf9K
Gdv3eOqSi0BuX9k+kwxz3tBAthwwYk6fmjyXMy6JbfoI41+gC4cdx6iWtvariKKHP2LdlpyRGdc5
FzmjJ5jsJt7dzWCIIvhJeckNknmAWm48+BrYiCQVy7zjkjo1IiXWYcKccqKDACrr3E/gyjXZyLEL
hFeELnSyyHw0ZyJULWz8ePqzROzggYOTjaLcZAjQfIluifNwrAFFX/DF6RiIz4BFB70DKP2+UKAV
nIxV2YA01an1eDVxILMEk2dSC9M2WkNXXvvEyZO2zMIprnY8++nGekhym3FHzTpFdrK2QFXZ876F
SpefxgGmbXYR4XyzNSeqadBMaejx3KHx+VvN6eZPjHDK8yENjei/elI1tnigfN73+eQXn38Y8MlT
t4ENC0anXLmWJFt5v4NOnj4zaMLzcogLw014VZXoiqsm8xraMrMD2ztZWtGb2USqj1EKkSOhB6f1
3wPNuSBg6Okixg5/8nEPgVIZevmHYm8x4xuTyUocsk6Be+1lKMStL6XM1XFw9bRxlqE6r47Ecp+f
ekeOH7bQ2EmdzJ1HEXLcOu/LqejvHqqb3xzhrNM8S3DhWBpyFEJGrjHAIC38GlwzvMohmmfFgqcb
y2/2cFJTJ6n1vtkX0fvLQpcpXO5KH8Qrz+Xpty4lyA0OJev06SlCFdgq5m5+KGAxIa6I18fIOWtf
1bUXIyjmPX0kAeRtDIGevkniAIva0oxc27Sa5fFrM9J1uOhOf+EAiajqH1+jsOkwHHp5rEWkAtqm
f5hhWTwxt2q+nze67nycmoseWawBAjOXpGsHteEIpzW5Y5pspMA+48SLLrLyC0MVy1gF6zgDZhEd
v7aC95ksO7K18j+xMEmGDlcSjTBUe9nHGUGmaXAlq6i83ZPmvsIEO0Z2pdfdryqn4/7CjwImDskE
j/TZMP7/PbF9JJKcaYBhGbxy9Gtc3lq7RpESR1yciOmeGt9c29ITNjmy/Y+BRkd115YTBjJMRXkb
1E++1l1Y/pVG1BkW0KxFE+bpZWw2wwQ1Zap1xVE3fW5FyJxd+0vCnEW56+wvoYs0NXXBR7XMtdgO
UzpAswvyPSSg1J5kmV/jJ7KF8k9H93tEXMFD5QFrmxwL0g+lP7y/4x6YRdIqjRcE46UiQG9Ilqf/
uIhP9MtffWm1wROyQzB9ET6KXSfkD1/3J5KbVvybqoeiEfeY3vTj8CNOYIpdnGuu8HlrR9erc6n7
XrdnZu7QairFHl0p/ip4Fp7Tk8986lpHxtzJfCr0V8qDaXENwK4GLg6qfmRBr0TOBeID8Qd12P5q
2mYMxaAMIiCdMCwezDlXz3ZhT4vZ/w480Nb+odrsfyLLA4Lup258RXCLOykwM1xmuoqf4DEOhxBQ
2G5EH61R7B0zDD8E4nVd4ISH3FA9C5GZaZ4w7cq06KFhIuOnyt8iMbzGBuZD/dF4gJVqIoZCWFT9
celEgyEwafsy40Z5gksu16Ld2xRhimSV5M+HhZ8hGZGBNXszZilKoIau6ERGWr316pw3JZDJUwMm
BBQOrxa4pJMzicC6mXrdImdXayUIkQQQ5EgmYBPq02VFGx8lEBlL4aqL3d12R5q6YT9V9Zw+JdNs
xqUfDSvZRyOsIYbAvICXfEyz3zuwHmRy4Y+ZdBfusSnA124BHsVhmmkhGwFVHmjGsGXUHEVM1Xda
QFshnl5ZGTn5aDwQlfNWppqQVDnFBqWQx6AzPzITE/s6vlUyZTF2/a2rMzYpGksJLPpEsjSuh7/P
RoZEncsB/cXEKuAVKbb3tETrEUi2SS+FEh3ww2wLYXpQi1b3PhSWJ9jGI3fQEni4s0a+I2MMSLb6
Grb+ZJZn6zdpe3syO/5tIVLvPvYAXdt54v+WMUe3DsjDNoyotlfZpnoUQqlEGKKBrzB7c3SUyc21
0yhHLyR1P6BYMYn8WcOMCVnhABwDzB+9Uu4TfXQV/H1LIB68SDBjjH2UY5WO5H45BE2xkuwb85Bs
s/boyjcg74wnt5aUatFOH9D3BYrw9ygIpt6l1oZunz5VwnOmLnnmGKGsZEYOAk+CCAxGWGxj0bb/
H103vdQD8PuN+k9nyvp7pUdeutbdOi5FRfAyjX9q+8QNfSNt6iStZnz63Saj1pRT+GUyjKIleIpb
Fd36QOijSl7B8Hg8uuQ6N+/MflFWbXDYyONDILb+qPQLZV5oY/MzAqKLgwrAKyLL2wKD1MMrM2Xh
Yjuhkb4VWzvo/533roL3pVf9WcU4YNd++F3TjyU00bZN723pbFjQsJBQF0zYyIv37iGXhs+QU5x6
Pnh/kfr7VCeeoFJ242I73qJ+TZD6fc90DmnumwsWkSidUOEZKl4E9HU9D1joRafGmKn1n6QXwv/h
YLXCMU/PS+QJ2sqilT1aMckwe/iw+1xYrDixo2CF6HlcZsE51lq522J7+UpQ/9+aCUwXbWVywEKB
Y/tGO0+uXKJOvA9eddzhEtwh8glPzLAZGDmdlhE6R2KJLkZdJSf/hxEZ3+v4FChneJzioXr2WFbj
/ZoY4Qvxzo9R8SqGUzB+tBDAklqfBB+Y73nba4xMIIYFygW5UBkGH/l2V0DVCQAm26VbWlJyeWtW
1vRCZFYNmyW3rDHg5BAZOdToiTweP8DS8k6qTiq5JP3sqK2P5ZEd/B8mep3Xsys/FBcOKHaYpc7d
0QKYRW7hvenVVCNbeB6lPZd5MpQqUJ5QFckcx84sbzLDUe5iMzT/ci5rgnzqhZn1xEGxjrnLC4M6
6olqn4H5OAPXpYlc4K6/UMak3FQx7J98ahShQAI4KynAdOb/ZJ6GYUPC2vMKEam8G+JQhTott6zI
fISnA9bzph4f2ckMYO4D3lEbGdyl2ed8hWiW6ig9XO/wcuYyp10Dg+rR5FeOS1G1PV7uasCgUSe+
Txxx47dVh1EfKA3LUeAB510Npay9r9sH9GSWaS9FtURfZSFrbX2I+pz4Glwvfl8dB/f+mO0bZVx4
L8+vf5EPUI3Wl7FwMZahVqr+4AiV1WMlTe1c3Nb6ij76oRqi+bm37flMw5OubcyMDtfNmLwh/LtY
ozvP5v9ItqsWtiLSuI58j+f/oclOMGz++7TUHH4GR/SHLkQQooHucgZkoovW3w/K2RZTqBH5aYLc
m0GJEAWof3AyoWGzx34q6gh/tc+bgkNcvfwAD+sgGKbyokl1jU/w2vp6ixixtqqviifLmw+HbSIz
8au2UrQNsFzk7GVT2NZ4WgwjUoZDsv0D1jnucPLtFmcHlOWQbzBwlBHO5LXcB0yFmTRFL5BVyOXi
GjaVcoA1x9tpR8k0buhFtK8XxAc9dgrSTqsn0ubEVvWwsC8kzQ8gjBOVk++pbGGl38ASI9M0Zd2S
4PiaZhixfC+yqJ/JuL78HZgJIi1sDjGmbHcrYyg8CbKK684w2PGLxktdF/S0aeoWagKMwIHyOzIp
7Ydaav/mgmo74VMUiEeZF3EeetS0M+7X3cn6A3k6LFZJntw6CJLGPMH2bAB8f2Cz7a7vnw5+sB5T
jkKvXbd5MtSp7gbqhgLn6h/NIhlOQuYWBLMSlM9j+Rj6DeHXKSzL4S6zn7mjr6slF2f9YjOFJLEn
1qUwaUtZrQ9pJ53EMQ2YwpG8/XN9B6QSL/CdaB388PT7e8Sc2HJV7mql4H2+Fi3awL45EQj4WRrD
FQ+Y3q0enknmg/7P8y49mQLjSA5T10eTlMMhmtDhxb9NPhcZ/GT4j38CHQLf0yuu6kcJxHio+ecD
6ojCDSwsrXfQPsy+647vZwL8NsQZ5tzsMwcy3LwpOc+9btTnfNbg1lhxybj/PE2wqJCGphGuLnSP
c/kd8U880p4XL2zS3HIbZ32L9huvax9yyMCtfNeRrRTTw2qMBlcIBoW1tO2XFA8CVwoL6cB6H++W
NcdIMAA2TMpmB4SJtDFYPWEFQKCbCgaqI8Iyw4c4NZwQ5sJdIvBvPfRWtYszAqIaWP0O6/2sHkxr
VUp1s17rgaRS8rPt6tWzDbmd0pmLpg8npfKoiJdCk24bup71ZBV8kMUmMtj1zvcesPqgUhAttpae
5Hd27EXT/dd5AHyLzLZWxzslN4HfdOD0xN3rSnJBmpj2ZNgbBA3smBu7om/6EL6w1UfeS1DxbZr0
huBoK397H2Rl9x8hWhASnKK6nvbc3zvxndlPqw1DFQ4VDfC1uBYlEJ3XaHatxQP2IKvGMyZJq+1V
nfg5zD2DLvUCphkSVAtxxZkth4jRhaccU4Haah7MeHKA5MiBSWXg3pcftsUP7bin8Tr1drX1jXll
+5p6/g+RsPI1pFsLTKoj4XdsO49Rdjtg0EoZxSWYwNNh6xcaJ+cV0KsbN3LRgwcCtUb+NUxoOuu0
55rMlctKBKn9ueyJuNCbnECiEJC49ntFTq0rEzJnh7jtf5pHmho8YVaTZUv4axI03t3CDLjziRZI
PBWEZD6plDVOWS/wLq+Vlq2qnmvvd6ZljSPDTRHj7pa35BtE+YNdt7powS+emsu9qCZzD83orZ5S
iSZsBvyNpW+TL8EW9hNrSDeb99tiKBs3KZOoy4K1u5YhPrjfsOQDLuTuUrdF0YsFoUc2/NbRK8/G
4Uv7cOuuiTlphE6GEyW6tcrDkQ6kqekvESoqYeFnlPfAuy/7ou4w6XF7fsimLiECGVQV+ECRzNzG
9QMZVvxVc7Y/5SeA02tx3EkwwixFcWWdaXTrOc3wFH3IuQZBq8+NbhmDsuw2pgE+2mCXGl1iz/yQ
ZJht6kEo+qSH3KF8Mhn5Kq/W5aEIswqtF/MXIGN5qhgEsRk3U2JzZLtWemwtdRg2T65k7+3J/5B3
NyDPLlSt+ZTgOBZ5niZoanS9YT/gqODqS9tKpXQCqPYcEURsdQ7IOTEsYI16Kh35wxIZZ5bUINSW
EjzzYzRtDsBLCtrRanoin+9weGenZ1h5jJcxfms8uh8FrESoYqd5kVM8QKXfLaqBqvZ/4aSRLDks
L8LbUCZu5VRs7HRRgM4bHSvTwxXYf0QL3Rn+YeLQ2mwuKxL9acj9LTYMZCc92gmw5tzkDb9l1MuS
fGaXaBJ2M7Etux5AapNHY266+ozvIgumohxfcvTNdRTTPEkv60uqVyeuzmZ0jRXic4UkbxcSW+xx
tvRAicab6qennQoNogrfT1be+mWwrAMUE3I7q/uixf+vK+aCNGKcoxzlyBLFAW8gVMQ0FvgB+H4C
0fumOPo3Ix5PcpIdCRk2mcPgro4txJBBHi1NREQOnG1ejBJph0aGqFfy3OgTmbEhWrjujCL7VeJl
Hk6qKTDYYV5t7ivLqhtkfGumLFgVH4o7JtCdsCMKD/jeV2BlOtGvg2PHcGrC+iLo+T33I07K+a30
sPC6pHuf9jgTOtwqhNcIEL7Z9FYN0hejmFXuXtNSYGL/bC4+Wt0J1cNefwStL5pVc41xjifNSe5e
3Kc7nVANk1qUVimCgLLzXYnsqCnNyZK0qSVN4fAzYEW5YNOaSaJYcEDbH8p7ATYE1wQeiniK9ITT
UMSM4pwKlSoPGXZ3csZnQEIP/uOE7IyS9+dbYFD+G+zIxLqqbaDULCQBOXwy0L7haBW3wZGDaa44
ekpBMw58mTvYJnXqt+I9rj9IhNFEnpp1Yxiyw/UtPtSj0xOYJwmRhZRnAmudS+YQgOIWpTxboj6f
bgnejRylMMpUV4gwUgHLjKJ1j5ZckhJqLHIM3j6ehZwfisATDhFzNGnplzuZFpMvt4CTmt0l6QWe
sJwa5dVDqR0TELGl6yApUZ4SR+yuDLmj+eFtwkIGEMLzaIDqHs2DSAD06bQVfsUUge52uA4aJiJt
Vz8F6EpT0Xf0c8hym+EJ7GH/kL4LcCX1hw/l5mFliIAChqEIH5dO1/q6eLbttL6DHO1upkz+6SQ/
77CMm5BF8ydvAoY8n28AkAjA6ZFQXnel7TAOJq7jW6UtrIYzYZDUUuvjXXFYsrlRQjuZ80p3bidL
ZJ2y0gMvgkE5PPtTdMMQB6W3fPXxi05CihlHJWzxmWvmRZHEd8Osjv0pWKGWCDKfWybzfYTYwDQw
GjITZMvH3bKZhdqNcWvpYLTg/NVSYt2mHP2Q1QiBUpjW9P74LG7crg3qkrApX4dfQehIWYKrHE3r
rdOtrz+ICG26BEbWawHadWPY2iwjqU5MGPfewiB9/edQoRwRNPUmjjdjqJAgSrG14sVcLx2UgOHz
3EdMO9ElSXpHfo/HMNyDKvojHPFhOp9ONwpccbXre18ynpocN7maQ0YRRmT4ZQpwKfVdWUtQ51mI
3Doz/LIHgowGoBw4q/m5EE6lm3OBqZ98fGYLgGJ71zwzuU9ke/Z9Jrkih4QE+N3PLi7GKspZjtHG
fNM527GpKIDhx5qoF31R3BTGuCvFqgJq8uXUDHLy4nXVmeVZSD68bkW/W7IsXTEJXN+LQLo/emxv
b3JlfS/XU+nClWzzUcrYRJQPyQ8K2sE9xr+L/K1xa3JCZSKI+hspNMUgIz+VDkSwm4aNFZ9FpezM
8XWjEdZT8ADMqMpImyylepxQPAiSWi7tqdF5cjrgOguLyDph/PXKc8hLz0Ug2xwm4YgBDXMPyJAN
ry/7DdejjEA/ZDmT1Qc/3z9Yi7yy0Embxy9OtSg5CDHcTouD9BhdRtVskqx7A2QEyy6LQjZOhjHf
WLDRFVx2068242mt3O5fBDrwilRZyUmH79F8cCfS4e2FviRxatPYNmHnq8UqRFDFSGjxd32qfV4X
HTnvYMlyS9jSTRURM4mIspOb5iTHZOCxLE55rM8cjHOmBBLfeWzJfQOUeaAh1GTOc1djbkeF2qmt
8uFG/4qWAbjiPMmExSlUOk+E7Caypy0MaMgNAgWs4WDkVxFvA4cor2aX+VTpKRj3qyITjVMnbQ01
GwrUd30dxxKp9s5ZlTHtCp9oXjK74OJ7STc+o6RwEk0S5qt0+d41tKoHYz7gWeUzgYgDQl8cBptG
LgzS2azTyFOp3F4o9rOseQdv4TfDZ8TF7GwQSo8+8hoFWoXzFnjLrwY9HqGTHBOYDUuVkJz+/cPc
RhjRUUZ+6Blo+FwF4G+yQKBrssCqUbnIB5SGgFaTIpQVrmfrPsbm3RL8kXGb/BQGWdAAYZLHLeOs
AStFemfighmPIvmAgAyPWQ1bDL692yuk1zmQHGt37zi80hgcvuATqCyhiSwvzZIPPfAAqykxthrc
ETUfDUby/7Ho4O7hkELWt8CUu9JSswmvbyFMBS9zJhCT3o5SQq/77BLGdVvb36v3EQQ7gAYAELcC
lgjuxx6kcezqkgcK51aWI39BVyxDXsgc7gZ+mixAi2sGt19zyXNi1gcsDDtB0Af2MmSll7PbJdbg
49dJTHkoP7giEi0o48g4zJaUEj+3ePWuoyDLTVtBfSZV1rhtJRkixFUhweCsO3rwbho6L8aKVFiG
8bb2TzA5pQPsNlj7DGMaoRJvvkHVHTYzVNWDHX/NamGOr5kW4jPwXTUh8TtQnU/XxZjP5RIw85yB
5nyBLj9skE4uMEgEwwX6S9zg8AeWrrfNzufGkxpEiNxtfOrypxCv7l8DK9OffOYDD59qHf8sU2u2
obuhj3mdA4N6MfmtEhPufC8EDkE3jAjX3EKixdZ9YduJrNNuH4mQRiCkWB0UzPAoQm55N5kHhoVX
r0QwUaR1z66lOINIz+IAbq4UJWbFroa1LI3Wgyg8kSVL19QYDjKHOZodoaK2sHN6GzNRFqZZ1Y2x
eaAwgsQyntiOVJEoxBWcP/9dNuMU5C7kdYf1IKWvpjSf7C/4fYnLHTazyZbAbwkucIgqKLghPJmB
MdM69TJ9OZKQTqh8nUV7IysA1UBi5RJM7aTj+skL3WScah7SeupJsRxD8kzSp2CwItEN+BJ8LiBU
1BX8N4q5u5kC01catq1CjMY7MpLLeoXX+QciyZXhc7WTXBRwLySu8VPbde/DJ8gMqh//tV/TxkuJ
SHOjr4Jdl+DgCrzjayimmj9PAemXe2vFYwA7BXjO+A+kV2YGvqQd1cSfTM1OV2hL/g0ququ7ms3s
GVsN8jiSys/Yd0VbvkayxduDEgQSrqeylSNLvYskDVMoZUeA/FC3GHAmEkX2F+lIQ/6fjN0T/G0z
aJV2G07knWuPdKo5J22kCpJbVpID49uas2sjjsHu6cygUaN0lYKt1yJGUUO0mZTXZAtSfVWyWII4
sPpqW5nuSQS3GQodEPxCYmtayLVgm9pUrktD509LprtI+GRlZojJEiHcpnkFMHy9kd+cz3P2JUYJ
DUXM87x8r50fU9+oU0oKisptivqH5QiP61GGHBU2M9JDjm0DHtYQS6BlleKktSATNWM+4DoRxm1m
IrbDB/lGSQVPTCZtNAwwRNzScw1SNXa7RhuqWWAMmueJ/auQASNPmp/ZvOYXI4C8royXqS8bwyL+
kwslREPjAmOnKiy7pYrEocBFVqRffCyezBgHZ9eerQc7RpGTzCuP7VonmkR2kXwYZFYvVv2jCmJy
N+L7Sd6FwBor7g608ZUSw+u6Siaxwx0m6wotYccgHCHoBSd4MviKZVKzIGURRttyFtwNqIo9RNkf
IAneEouQgg7z50V3jkBZg9elO6wjZqxkm1jFbWlRVzn3IOHSe0offloQmtdizLURuHeGxEBsPF1N
qou8Y8tb9z6kMARRklU436JjsHTw4IBfKq+ygiOadqPsRrhgf63bN0BLBMoTjC1jOqL37OihlstB
djfok5HrwU7zkGyPBmu/Fnd4n7Hy0MQPhsrqQ9GqbZaCSTRBJXTl8QIB3b/t7OKQ8Zb/DazsaMpA
bUDWh39iz2iKzjVmxtsY1XKy7IER2TCPgQGXn+6U7KFr76F9Xc5Urngr2fnSRMRcD5mOXgg/EwY6
r8j6Qq90kEVoGlzLcwrqc/FiVP/FayhujonRDoDGf4GDsS/0yt1p6dL0nWnxbPOhB7R3WDwOmiEW
bN2Hh2q9af+HFOPNvFEwAG9MGzG0w9JkcjZM9JeASPp0SNoUTmlw8gkpEUOflI2XVBNByHbWoeAc
jARVzzL9K/ZD83EUS68ebZ5wEa0CGrcgCkNfFzyLnWVW6LcmoCTVo9rMh/FUjZIF3gnij4dzR625
py1PT0XfQItW0E+n4szGGCv5ZJIqIrNIAQVbBVXOytqXv+m87K/X2TWx0DcD1jYzXZOUP0GHAoeR
jryL2+4iglh0POhQjC3wMn0nVp3VLN7//IomCGihIGgkWh12dm+N+EtTEry8iLLy8tgsk2MJh+8W
rMy0cfNJWEv+P511+3Moyndh60yJcFNbS43qeFy67OTNOxcRvau/jbrNCk+wC7Xi5W5Q9Jt/yUAX
kkGQohI4Nnt0mE+Hvj/OYxTqRlEmaEbJyCXJpywNWAcUL5WQPRIJpRl3g6CrzWVoHDFkdzReSovz
tvhitvoYN4oCjV4/1GgjhwP0XpVhuSEP2EMJ5vv7cS5/vef4Sj8s8xYu39uDUwJZzpHRlAq40ss3
UfGcUuBa7ERUsUY7GAG3dw75znMfkXA4fmvzJcGO4R1mTudbpwoDKVLUwA0E1flsv3x68WeX0A+k
2Ob5xH1h6B93VdGybZamcS912Nvhatw6hNinWIUEI+/oNEyNFDoxZA/RH9wpGg4kmizQefPjczCO
zny6ZlNM/V9l/zWBStd03cUdTTeTwQkTUJT5JA3UnSaGRYmZWvXeLq2bDXtJ8P6EOfYu3RF811Az
00qEg2wUc3KJnIi1LDv/f09HUCSaAZa2xJnR5KKS58yRPsooYA8ISrDg6CkZwxBN/lu8C7oPMQ5N
Tu2NiHJYlP7hOVnueuGVcYZxJTG2WsruxyLaYPWJVavOxjQJ4GA0ghOBQMZ5fvrRMEz9oetnDz/r
xDVjofa1LDV81LR0pdUa85520ouegeC6kl0fY6Q4kPc2TPLytwdCEOtpUqTCZ5F8Rrp9SP7Q2BnB
E6nwF95nWOcbm1ZO6QJVQDM8+V16YVJ/IA3KaMgCjHpxPy00vPN9cVmA0smS2tVifTcwBsjw496i
DzEBwEI/ATx4r36buC4IVWV94CveOYtayKT+nC0MoylSdNdEsuYLn/hrjCNCkNwoE8VIWMsjci3F
rD8Eai/gPb/1EWyDyp8IVCVzArs3NXlkwYfmcK3LS+auk/Gdz7G1iXyEd5HcE36MWapTGcz1Tf1U
h7b+VdIOqZwWQtgqSbFzMuSIY1lWyj3zDOl5VjsL9DWHRlHZM0viq1KiQhVl+cc+e+h9Z4DqsP6p
ivwkv2HEDpaN5snYZ8+16EYUONh8xsh0IlSS+mbFzAHT6Dn/NqSHDOLZuqqDEpdhDRp44gcGbJCp
LJvDNFqy2PPvP42C5JcewZQ2CNPXQ/cwQVFZAjf/glq3mVikPRO07xaR8ay7pXvvY52IDf2ZwLSu
76ETv9R7hCmpykMdYK8Ktc636/jSpsfitcUNJuLzDQPwCw4nDM9ig83of6440Dr8AC/PV2/1Y8sU
JZqB5FeyNUxRIUgABLQRNQQPetg1ATLj3A2R3q2tQPZpZ/OFt8B7Y7K43OAvI65TxOlt7IPc4kDH
QazYiZHPXQTaP5kyrO2vqlG9S124aen2duwnmuPneVotomcgL56wcbAyS1z89umZvCoTXftHXG87
EReGagSIbDKPeQA5LhiWrlmgjDbn9wVCNcERrHfJd2IY/Llm8giq1qEgU7R964hit6bLC+WhIG+j
axZPSIQkSU2idOACpQ11dUyXDuiYM8SYZ9TvgrvYmla8QunYYxVJunEuin+o6h5hVw1xWTMOokhz
2tiHCWyXh53dmWj1C9N1dk5ViPBwxr5rC6c22vPmaQL+NwugbV60obO71phhJDAnEmMEcE/DYD41
zTbQyXPIy3+WIvpjQ7DAm/SOoKpkzj9DC8CMGAKsAibpk7GqlUdeuAcm9J2X01LJnQjPM1Epid5w
JHHUEe4o4FSPWevC6WCNVVDAedVWC3DNtiy5Ch+4tZpkT3eEVNcV8EBV/h69sjG+im2d5ndONIcj
8VTHF5o1yyybFeMZ8dhkWgNfO8g6otemgsdvdQk8PR89IZYkKHYJ/igB51BnBNY9ngTQYMqoBIEi
8c4hTXHngqQUx/uW8uo4dGcB71b4rYEO8QQpPR4FHEPTi4MJvhvKrzDxqfJv5lzo9k/3YfVU7aUA
H+qMDO75x0JCiS4WI/v1W0etLPrSXbEvan4ppxfhADHzLTO82aRws9e692wlQHCxXMU6S4oYNj+1
7ORyYBtpo2eXgKA6f849TC1tO4+7JfKrRZRXxZMWXTF91vG535dgFChF98gUtlVumQ5tAiUatIjb
WaHCmXDmiFun7VqKZlq6PruAAUlO49qMyM5dXKnhlRyL2LRSvfk9DmblYF2VonrKnAqQ9J2so7CO
ZZcPzdCWJp96hfhkJTpceOSwuFkGAT0Bb10FRf9lo2Zxj12hgoDUwx1aiNu+i/Q1JiZ43GifMVDB
L0mNK0FV9hHpyQ9IrpfEljOwLtKCOKWXtvheixS0hU6FFGWCUxKPoIzM7FrL/6garHwFHuNv9GW5
8NoKN34Mny951M/eD9eNq6bnODWk1bdIbfK9av7fV+q9Oph0O1sTII2VsWSzmiyhr8HGuVKMIedK
kwBMW2iG6EL6WPdoCa9os752TxhCDtbZOGkf2AWGvQFrZgC/toIXwrOi7k8L40yhNOIM74QzaQFl
WcjFblwt1rPRXP9cSGIcSzp500RIOX80X/c+/pu0qFX0ChF2mhMc26cueSSrPcXKtGm9Cp2m0Cn5
RDBjd4LMlRECP8A9ULDiIytrgUp9HrxUbuhYdxxa9MA9UE9CBd9/QUU1AfejD4qQdCWf/lF9Ly9W
RVxjr4OysfH7Rd0SLg10Y98yZKhtUe1/Opugxb/la2SBHWOmXn0JHKImGEep5w5E9y8hlUIrAD5M
9rNlRNZ0IDMkn88f6ql4PgMzWuHRMHTkBiAnjQCYstlePuqsm4UUWc543A4IunQ+XjptXV/EoUgT
6V6CQYYpyfYp6LPhp8RYRIdB666KyrAExRv47cn6zWGp00cEDCGaEf8dJroEJIQhLvTL9bD8R/UP
lg105XXe7iuK6jDq5FPtJ5VUCa0j1b8h7+4lFnWD5m2iD2uP5P8Py9Hp+LxgAo+lxknW8ihXKdrA
a10pwAPxMzPE+NiJiH+EfqunWrfPugzTCvQjXrtgrSL4gftFGKanBuVEdJBt5FZYZ8+Yai3C15Jv
zXb2ezyGK0P/bHwnkvzFYXl5NvYDFupsBJFmlx9vER6dMiIftOxDERGTNh1dbnT0WU5+9hVO7B60
yfCx6qNOb9hsxFPVrrkP2v7bt+STYklvd2Cp5yN9qloJuk3lnEa8nfpb3wpE+f5IvBCqMRSNL8LH
te/89mmINfEJ3eLvv1F2X+IiHokSm6+2ExtW2lx6OqWpRuLDldl/RbQ6Gb8RD0iVJc/Jlr+zSPbJ
uXcpQM4rx3dIXi4YV7Bd65UXJIcqyU3waaVSpokTkNT+ODWUQxkeYsnEh31CJnhEKz6sCQXnU44g
DmsQvuGscurWhoXRHqsTY/RJMIM0IS1O9R+ATSRGEkHhQgrt8iHUM33j8dbijjC3kGUQzRmnGBhm
/vDXuXOEgDKB7sAOf2bGKYw4DDemw3KDyrRxYqiIh3Qf7q5dTwJRcMOZWEwve1x2xm87y7Tx1oCb
GE96fGLptKgqsSFGnaVCuUoO092xMbNzrVuLGViOGesRz9LAute/HD54+595WHb91WE+FzTdwCWD
gjp4jqCzCgqKJi5x4g61QvmWoi/0tz/f3qKBVoiODUJR0am5zjmoAWHGBGpyJH62U9f0FF6q7mT9
R2w990Tjf4YJTw0drSyh2fMTxr/A5Qx4fuIfNr8tt+vPCE5X8BCNAAzGcs9QKfzAj2FXeP1LXiIz
nk/YbUohP9POXzh8eE4AjC09n33hL6XXOsg2+dX/cc+NGmFagIWslly8rWcxanK5gF5Kqd+KM9q4
2uZfQAvvFCxWW+O+bHnA/ctwUEBwCTtVhYTFNN9wA3vLy5QIQmDDQcQ3eqBMZIzE6GJ1k1iANbNV
Xqj72LT2/GpK09W8uj7JhW72IcafVDGFhifmdoeup5rKtUscT33mvqVp9Sb8J2lEDvCDY81kbyFJ
cNqzjL/2yx7XAbCKUL21JsPmrIeoS9kCSyTnYHeew0AFs/I1GpXEaFyCtQqLa31C3BEv1La5rqDD
B1NnbXtATJnRWTHoSASKQYkCE87rEmNRsFXAvkGcg5mDLKp0OxlKBNYVoYBAKPPgmChqO1/mB2fT
3BbOHkVRmaO2Kf/rEjsSLO2feazUXbvrkK/oWHqCF1J0h3LQtnxgx/+q12dxIDSu/viz1Vt4Jmi2
6KzyRqQEbP6loawMMYuUOGFPrwjFlGI89i6exk2/wPetceo2aZa7TbC58Yzdk4QJKrCBYstbdraf
5lEUT/rcxEPEgSvFnP89jFRI2mv+exw/+10JHE5z2hY2zNpf322yJZB6KlbfWArAgSsfDPPDuM28
Kz+z6SjqGXbL+MrWWqDKq64Rn6jRPU9hGvMOlmeHikifZgYdAIr6eaz6ZbMuf/LG5oIZHlBEwIyY
K9VIYq6qnNRdtnt66E1htruiuD+b3stPOhFDixf9MfhwX8VXJdKE9+WvU/PeuDCK4+YkCCYpJJ2W
0YLPK+ZiS8C/V7W77qaFEiNpFOvyYmEy5PummQQtjIw01mjUnocg9m0imZkfIuGTJRMOsoLkk0V2
vUKeIyXjApGLpT+wZp3a5KXXXiZdp9s48AqNSHH5XDWaEsEskqqVXGLKvpZcD1AjQfQ6gNo5NLjm
so/d6aviJsiRBYymg+DX+UouF2B4E7ar3Oc2u4QeuonVGAXatEuHkpdPqXXs4q291xIUb+Y9gZOA
kYrZM2v2j0kDLLxUkbhAfRCwl9D/jatvexgIbXVwtg7eHgQ/mLGrji61eIG5vdzA2eYFW002ojuM
mozE7xEXQwKzg0wmwTwgp6PktduLvowimmV6MckvKc08mcwvy50g0OqqyNwHtwJDlz57yu6tPilh
ZZDp6fCiSS8dE/Q2HvBL4LDR3EsFL3XZ+Ne6bmxYbp+lQUnL2vykLad0u3OCyrtsToA/oVuGcbt6
C5xH8WwEbOF0T32OMnWhWuOVOeTOZ10MugnMLGjrD1Ad0+6XECRQmBu4aFV2xlMOC1dUgiJUyMr2
C62oUEDdWg5jOzKoXcBh1KdBYunTp5Mv9+Q7QUELGv0+LTdwE/19DxzbO6rj/8UEiR2f82u4M0kY
CtInNsZkoi5CjWVFEgg5POyuHrZaaTxZU8658U0iLzRtvsWxwdE1o4eATefIGR3/snxLsFR9qrOB
gT08vsxPnqrjIXAoWxc5rNDiXSERHc5DKJR2i2+LmjtYLCRkdb9oemKQme3I0PKASXK0uuanWcKQ
4ZcciOyQQ03bfne/Gg+6QOlvvrNaGOeSoBkLpwIEv6idMq5gJ1AMxAIBnX+IAkcQSZlPbulX38DP
9IcM/ASokF0fJMGE6iuQ59WGpzhP2hCnrW1IhC7sWupb4CH1EQXkBRbqq7iyEPpbtu+CzHXz95nn
vxxyUXOrO1hmv45V+d8NeV1gtSMwfneE/3sGrBtV6tT9i6LhqAoQ2WzFMKPO5AkfAc1Gm86OHM5y
romZ7xvhXzjP7/uL2g8r3Xsk9w/OSKzlTxHzB6iTu5v2fM80Fpvse4Hv3ACnx8N3b3DoVPar77DO
eW170ABgupbNewRBhqH6zmtl6JLRohvhoZx7Azz0bRK+2+GN/IzyBpqz9sqf91UQIGzSC2XNzqbA
eum1xlxI/jppVs4zzxtHEnFufEkdYo51EEcJgcDPFDXxboFm42G6LdJCA9JOYYwghBoSONiA8oOI
F8k923v2HB+WY0EP2R9HCKLvRwI6/uplP9NZX7uSGELtlzonZG7H4/CrrmGsZUu8LBVWBv5hOaoW
FTurWUKUQAgGHYoAIxBKfjJLr8hI4iKR8r9IL4UFHH9jqO+xKd7KQIhLI9D1wXKHiEvP4Gm1inLM
+QN4tb/h/8g6ERbs51ZRCIA3XAcFaOcBWiIqy5/7D7bM5clHGWE4aWL3BpiK+vp4IXS7/9b2UAeT
15f9tPJrArGx/V2Bb1JdO4OuoZ4mGdLw/XBafFxe2o1Pt4f7dB2IhghHubLr3pXj8ApwwaoMX1GD
OwWVAs++eEOsAxWJYVIzp5FUP68XcPkK90nQ6Q1g0JWgNZ4/3sod95cEzmk8QyNrNp0w0U0NoQDC
Nj6lyvzwxLqTtlPxMXGbdzRSQyzB4dBF5Xa/xKoXq2FTu7Sa9LXIcIqH6VjtI71SPvOr5eS8Z7tO
cH8PW8ikXPu/TxKnIdwfoX48H0blVGimK4A+p8WiPk5+8D58SqxFpM+YBcwSgFEq1xOYfn8VyHil
9Bx7HVvxxZq9Ptt6MmrkmSz4PUiXc+EiAFtPhyFRG3J38YAclsG+BU3u7CG6S/FyU8Xu9uzbesVS
zw1GMMpiUYYesVaQjoL6M7wznIYb0s539vymuiT1cyJAXkE0J1q3opb8SD8GWgnv5sJ348h6ntcM
kC6IRzzGthKuVX5dB0ps4Eyvr9eQowfdl2sDjZiKc4izlxcYi9wxC78EmrNxdmxLPcytHUxfKQBn
A36G6ZRMVtOyhdXHvGQCzQXsq6UYGR/nBON3Y0ZDTGx41zwg/3GqTM1Ru35GoyAGMpCe5oVhb7Nk
0ONkrflQoBlU5JtpATrPKDQN9NMEICoEevnrpUCAf8EuwBeu33I4UL/1goWY3+dcE7okVaTE6TyA
rK+ZybCbQj1hELGqLvo7Rj7wP7a6S/1SlUJZN26sPRFm1N3l20QYXF3utA4tHyRfeAA73sqC6YtO
fl81qA4CcYdrswF2Zzgz7XCbI11qHZIwp0F812DvxcxwoaftfGtK5RNHx8SeUQyOlJrvdyqIGFOh
S6tEMklZtw+MYkhtElempP2p+qtCaSvIrfj38upAU85A9WjKywlUsYSdtK6oIAzNA4ivTA1kYfQx
AizjxP/S0MsTV1v4R9j6EslO0W1QfpNcOdksm8vKYsd0S7s+B3W2kS4mE9+OGwLwCZ18jxrtlZLr
OylsUFS8ThMhJDj/B0vKpSUCX3TjoYosxexM2OwUTY2C1WcTJytsDGM0OpFLlH6tFRmAE9lKniz8
Y+ThrdJz5xTh+XUnDhihRot/cm/G7E5eBbQxFSHL79Hy/CliHRMPxIro/Z81O1x8cMtakBIYekm1
GB8rwwQb9ryBu2CxLmYU2vvpV+IZ2DmfJdFv4tO4AH4rEnv+3KjT+1QWc9r0INQNBmHu+36abMiL
pJ/swpEyyTYiijLYPtGvxVw1ZhWlth4Rr02H6HNbD23QxbyHt1P5hKkXLfT/ipUYMi5RjmaeJZ8e
OPTmzinhF+IrRkUecGtXvkyUxHqynu3hH/QgB3g46SQK0jHkkn+BL2WkDJpeYg2QwMzbbu7DoIk3
4yG84qsRHKQGpdJ+l3XQ3bnSV8nA8PHjvwnWpIrqWW5VCxk/Mol4PIkbHXfoFhPyiz7AsX9xkgoH
LaTy1YgNEKMRjPn6LD4Ex6kgXUyZYwXJqaHxE9nWMIHwjdsEJaSsi6VktNE9NJuXKDiaTywfEOnB
YwMGdG9v1k8C1QC5MVYx7qTwsXEzTOmZSpcqUAI3GHMN4ZG8Cik9GD5rZP9rbaags9EM8bG77fr0
uWXCAKq0dgy14yBbA6U+r9u7P7A5TUuxSyb2xzrayIIgBYZ35OlcSgot3kp6+jDzd7TnWd3uxWW6
EmlYcQmcMdpUlfrNyDaKRJ3/X1Qo0o+isegkyt6Rb76OdSej6anWk5N89PvnyMkzZBskFf+SBngV
P9CMqBw+3mWNp6gntD6gMhaa2Vt1MesWFFeHuabRJbEnOVWAqgphM7TnPKfCcYP097zn/M52/ZXC
T+dtHLb55KfBCSx9+3Yr8asg/mpRAnYm5Ijy9jGj/pYk3Uik/vTg1rBtqdrhtksGZWAvuAGF0iRR
ut7YaXM4jg2sVMzbOaEyxH8a7quM46+LneddqbG6aarFDsnvb7jrkjnAw/gykL8or0h2fx/Cj84u
pNkA6NP83mgB86nPNSf4swMHyILHZIFLKyfby2Lk88E8VTjIQHCT5IKJTs4f38n1pjBFSdNzgSzz
AphGb3WsmhUbPEADcFX5euz7L/IXK2ArmvfVKoV+gYJKXHXrd97cL+s89CpDoD6Sp9GXngZpjzA0
9pGQZ8TnoYeWQS5oCOJGfWAm8U7zBo4eZaDWC1uy8cU6QPVE0rpkwICExdlR7xl8xEVd4MUcdLE8
A0yqEGiqbpAOzhzrGFygRA4YgZKRYQ20fV7LwwI6mjHUzQa+/vi+EQ/wvirKn2S0j+f8zjzZxQw/
lGUj+5hL9eMSHinZCiA8tS1JPL+eyLKmYgfEr15vgF3YhDBNRS3YOenqAVvKnbHXKEIHnsHnvVBb
Sx3gmpGukZRoivaFCIEg4FXkgdV0htNVG5+8PS3w0N2O6i173XF+QTfHkIbQnOP9EZYxFDGs1ot4
2QJctRAVPDYNPdL0r46iMY+13k6v9SnIcJPG1Vnb+Uj9vMHG7Ig1TDDi22Nlgm2+rNFKa2kt6F2E
Y3reGv3bh5hVi4whVDVGekOuaNvU+lrUhIZn3BvjCFNQNML7FpYXeC+prlpmG3ncma7HBNswkFJ+
uq8K9mTd2Tc/Q4FCxebkQAclXysisJQhZZ5hgYLPwfrg/RmIZo1KucwffJGPPeFTStauEO9qlUvW
FZ7+jlsQ/8J3VXlQQQu1RuQcZGlmuRVj3MOGpotF5fhs2FKg3nDGfDipJBD65PIemIUJc5vOGF3v
ZJGxmGDLabPwWX2g2+AKdneZaVo45r4YF5BfEhpqA9cMhp4/42eW2e78RIYFk181WX4455Io7gJb
hcfsIYN5BSbLpk+enDS+2onaFmMlWhpmO1FOKsq/W12aKFQhyXfLzrxd3nieMDCk2Tanakr9fX62
vKhNqjzlDDqSnNl4tl6ouLnjFnsZtpvUthT3h/+3dZbHHBOFw8wiorjQukdbKOa1Z2Y4PKwech3c
QzYkeIxVLRqIE3NsCfTA4A0GeXke3BRt4GeWTDsbdGhmIWQFDrq6WqDAMsKgmXScFxBAg5G0nSOS
VfjKRkTif/yO2pV3raGwHm7cxNySY5+/PmFFNjH+GV44CIxF8nUYD75ZxFTdBegz32sMLT+TRI5g
sEe0r32ZKVE8+VK9dq7vtGEFJrok1VXvABoqfOGlUd6287g4p8C60Q/64Y9jU2blzn25eslZ3ZfJ
ct1QZ1ApSz3ulwgetj3KJUrenUsTlu02xOZnxMD0piz0+gWM9QgqcGX3P/eRJTHYyQAwWTSiu7dE
WtpSKY7Z135CYhE7eUVQM1I8cFkGDi8cyvJh5kRxe2Ct/9FGLapDVvQR5TwBFai2IAEJ3upJ5dIl
4Qq7DY0ODWrvpBbO4jQRiQZ8c3Zp5EXasV51WfgLE3Bhc3nhlznj47GmRN1ojI7m4iDqcbrkBX/d
PT0w3xUlJVPp6iOpdLdwtXFhqs4/Lv64Nnc+OLYESGZTxvqUdi3JEZQ2twB0XRm3g4aMpm8LWNOO
qjEXVXOarW6VJoFZV36awh7Cpmmj5OEZB4mOFnLwiqd827GfvnJNLJBjbB13JoLgv8nFeioRDVBN
8L49DkKmu22nAYj+RGmOyr08F5ifZOupHic/iuOoPPQof0lfBq644ZMDHmOI1mOibhlWVVEjE/Bg
yRUYno0TqY6q/4E5fA/PfiyoK8e+a9PFVKdTuCj/5i+75uVue6nOpovIZdT+B6Jg3uxcIhjTaJgS
X7e+9cv6op+WWPRTqcxgZ6A3RBHhm22gbsz9JgCEdxlrLxDB1qx03OOFoTGwWwwxGfM2Sy8GMJzc
nCqTAfMGt/bJlFwbWh76SH1Fgzbvs4HIzMU8UvBSyhz7Wlryh7xGBYHW/N51fD2M190iWI8+bE+q
UD54xO2pok51OKCj4ko6htShghHBYAI7A0Qc92OTwNoShBKauRR0M6FSjV3p5jWpRv5DTeBa3m5b
rMS0R22UDXTroVLaFm7GXU+4o7ckK6Kz8GCLG/GR6csijE/ngZ/gzBKfnFthVGqGRh+k/+fmTDEh
ywmbgCyFFkwqqO04KUDRqPMyjTNfkL+SBRLR3ZmmskE06r8gSCnRIZv9/gKrZS2T2+vgAGzpO2sZ
bkBMOmbkJ0pRyn1PcK64vrGrm1NxVoMEf3SNpMR3iBoXMUVqTzN1Cvcku7BHOVzC0OhxbXD7uDQn
7dLgy0XRLeC6wW1OMAK3/gQjNCWtgXVnypmR/DRrKszJRgeSnYGFfMzAfW6UbCK4TwznXeefpH7l
dQunedFOEjuPu1QlBJrRn76rB2/GtyYbEJ8MZkfHjxUuDwOLdjNmXXqPvY0Bp7a8V5xxRo2Z6DjW
a6iRwUelTKkd6g5rP5ciMJvLC7nXoQ4z5nLfzJT2I8MyrNWwkuXiTcXHZKL3NPjS16orqb8LONE8
iBclf4EjAihgywF1fVfcJgPmq+UcefDb6rcG7Itw7nvpmRgIwqRZGFwBTD6GF5bMAOr348sYtq48
1QJruNvoc7dg3VvYixDQuP3XZs1cTq7DcijRQqEznvCOe3EubkeSs5NMnhUJckLCweG8qYii2/Jr
vU7e13Ge+xDsKzxvkAb+BgcHYDokEu+Aad7RFFCSs05HrTEuR8+/Il7E2gRSefpHvCet+BZRrMBw
8uHYUKurEPTVy50JNf/g6Y/g6R+CvklTWf48cf2TMQ5WrL7WFyKbt7ryII+Bc5yshke5cMo09WYk
W2VF+k14QNEnwtYBXURuorBbISKeJTlWpEZiqZ6bmocjLi4mNOoFdByasj/aZ01dH4M0vH2ecnfh
EDsEPiKXnQzoM9XH6rffa9jHHh1sIfewc4t+lS9o1ZxKc+tWPpE9QxhAfXMpCWzvaMmgGd+rfDez
A27tOnc8BhTdIvmgyPvOpE7E69JoLspF2+yCc1i7KGKRMfiTCo0bKj/GBgnMhgJIMkxQGgQoLSxw
wysak0I5W2DB5t4WV165RqcPHD/w0Q5ZdB2a0T0ZFexE+O1xE4rmYQaY9hsQTOQ91FjaqY6OSAzT
qb7npOnLIREBZcdAKfcvpkC46CZNR1EXiPpJh4zxd5MNltLRFAGrMYj3z/hW+kbC8gOmxFrCMtHp
JSlNzjhcR1wIY9zSq/c7Q4aDQGjmYXzZPaL53KUiySr7thj5yXUXdMCArKCAbZn7lvZUW6hAVumk
mI7m2rBvP880XLFNgz/d7oYLb3wm2pTuwHV81LkK1c1C64JVQ5fUdGD41B2s0cL5PopwK3lO5lww
o3g3DSkLIA5c5dErxzJL+hJseN5dHJDtDxIq3aMLnvxqQmoFk9tIL7F9FkpqPRAgfaSdzZssPa4N
IHpAw1eTS0rNisgtU6WL/ZfEk41icRqBU1jlsx2CkvesL/lJq5muW1nO9GFAGl4mbT/AgscL2iVR
BceoY4ZzgJNm2LBmV64MA82895npPkEBoLwqUqStbycBplPPt0vqPYrmBWd4wcGRpJpfuSGAoEyL
1iio0zXsWQ8emPuCGsMn5G7OBOWbmEPLs10sCcJ3UjkPMdaN5cJR5rSE68Y75vNgj/2d6XigVrl9
IKd4/957vr0FGULnGQthueS+9Ou6Kb7I2rKwKsFqOhQGqskxZIYEcz4qsQqbvf1LqaPmZvosRgCJ
Kr/5TWXNRS0L/7C3nZwf8ibu5+vn8W4ornvXJwJi9+UUZdPKZ7KziFb3rAz+/vOBX2DeC7RLnNJ2
UPMgv3db5n3cyYoHu/KxZQrgGx6jTMIFpxA5Xn2sF/jOnR5/U2XY2aSGnAyc2n9L674jNwx1t88L
leD+LnbcUjn8y3Xbjw7rKu2I9HJ5Wz98qZZJjUzeHDlRrfvZru1EmpmoWVLrUTSn5lam/i6+mFhY
LrIpkUzuZ3Ua9paXnQ0Anqt7KdeYVnTqmGHetQ5MqJxpIE3TQVFAYNFV+FDR2RGLeU97GFdEcHYJ
OZ1eiBXgL4qHUuh6Ks+sol2cxJMU3eECG/j8OW6qdpT6PUiE88s7SA++GACkXMz+/+CXiaB2VF7z
GOaZwIBUiO/hOpSFp/eexd40tDaQN2B5am9SHgY8Y2rli1d19az+6NDHlEgdNZ0RIBNdycdZ4Jya
3OAMUgcqybm6RVb3kCHil1Dj3dNAyjT0R3joKISEjZvBYzaQCl4Zcrg/SsIQBaCU17GT/VZsv/Zy
lAKqpWJu61bfsXPtex9t7TTnMjqH3VkTUoPjinEdI7DdTHcydux1+P9M0OA4NSPVLfosFvLKGOc1
SIq1TiPAwnPW8Dr7pAXZjs3qs02x0513YvqguW5BsU5i9oaHDyEGwXGx3ZH8uX5NDASxOBjDioW7
FuFMSUNX6SBeXoAoYE91JHvQgmhX6hQywtcXrgQVkdE5aTw79tDIj1tucR56GVLV55z5Y4ijXFvz
wCt1v1gGxhUQy/FaiGhGtE8NRZFF0tLvY6BQLWBSSwm3hLG9BEskMG3+vY0zCnIDq3ZfyU9shSUg
Gio09n4DkuJf+U7P4fOfGbFOMJg73dtd4MYg1zKrF5jjozaVNgpio7T0z5knfp0TaBhszXlgOG+m
yImB3Fwvw212okn+qtivUWK9qATF0/VtPgZshitchFVsriFF8T7b0Pvxrj5NHKqf4dIuUkLPFX2z
ZXmMr3/9lSkwzPWAw9bWyRv1MYeyrNS8p34pzxVeMSRez1T7zDzTpGLbaIdljV6FpfOnoM0uImBO
fEwhEc10EMdWkxLUwIiV3WKXBKZoO35YWwZp95GWmoVgZD9FjOtnxgi9NfusHRRBcSMRm9xvCLP4
x5guJ8LYbrzI53pbSpq+wj2fmDwdTndkXxUY9aHaDNTE1/BCZVvs5siZs9eSBmbWia1f3a69syLZ
o3EzQzLk9RYpelFEHzKN2lMVr8UXjyV6PqI9lJ2JFj9rNU161CWFAn5BE0c5xYelIWOZK0MUXVm8
9gATn5D9TDi62OQvj8gcobrq7sjQJzcc4+87Q1q0Bdqs86rgL6yVroA6Bmu9B8o3vAi+yHsAoU5e
rAL1vyeJ84a7BbAAiYV1gaeW6ocafVbHl/AdfR9P7lDrB6228IVbH4Ub5gCUYYInzCt7cmyIhVwS
mgDFgN4eU7JXCXqe1/yOCDd6FgP8glaL+fH4LGYmsmAjQw6ST0Hk4BCjyqNVGMszy5bT8TcPICAO
z8zWRLaXUIvbWzI8hiLm12TXIQGH/8iwCqoj0ltSm6EMdqPuE2paf4fNWG2px3xnl4ZoNQ28mZiU
wjQP+HT3jxt3b+e1e/z65pUfkb0xPCgeAQRmUejnA9ProsuhTQ1L4DmuNw8WK5w+qz7NVlQlYuRA
2xGMpsCVWFL9aRvbZzjPo8opoWJ5nj6RZkdAJAbgKOGTrXE7R3e0gRByryjgZLqd6E8zGnkBPuoT
GsMGhIvmR+oEamxaH+LrCLmZ5e9/39lp72X78m9GXBwb/y2yLRs26yaFcJw5KK8yJnlJbbyR4THp
WB/KU6Ey4sZIVdNxvnz993/lc+dsHIUqukwSR9cTsZuuWE87vdA8J4EdW3VOPgFHMfSZcMIlCwTk
w4ln6I3YUnH9VQS+vzV3G1vuZ9jrUljLXXFGf3ZBqZl0DkfpRH6ktfZxBEu3EMxVK5ylC4qv7qsU
3lR8Y0prkLtSvx3bJyGJBL1631o4D8hpBnUSe6Fxv4plahSgrmF9DPzCB+PCsAkWlf6A7XGq4ZGg
kKTC8llBX6QCComqw3JWAvTNGaCmhfpwk3S6lVY3GQLhVkN3K5BFYC7ho/EE+czqtH6n9ZnWhrFV
jJevOcgaUUZBVE5BauK9/Dlv56WCQS5thcTVfEeCqSdCrkz59bWbmJHFQWhj6uNgG14U9N46TSlN
eP2LZWxgCS6wpKfqYpuUsL9HUra2e9p2bTaIDnVztLZ+9WobsMxzcTqGMjmUCAKuiivF7Iarkm3Q
h2tSvF0JX6p9/rv/U694L01U0B9qcFM35+JD2wwLc6ystfWvVAhGazqaC470gP+RD7MKkoxo7/MR
x2nxfTanaS8NcpQqYMa2ebJuvzr7vUXD/dghm2yIUpYtma2KYjaN/vj7Yv0vazabBt3rgyq/LFiX
TEbsabSog7xVEzWxpvmZ/C/+DTS7i06tY2kg/YCpdBvaBwWY0H4yY9eOooLnkdqTTLsUAVPr7xor
6ou9QHEeu6Czix0NCEJvvW/hy+SfaJOCjRJV6K90shpmHmumrPsqKnFjAkaMfEkM4GxG+ewDJZPr
H0aLkYZUFTZg1LMnZq996koBn36FU4iho3NvgU2gmYRAog3NvsTzFa8xGa0zd4jk3wo5EE4+Ce9q
ndIxsnfCMn+Ci8ftcM87khiCoDgBNr7P3IRqPGEirsSAo8emgc625ubkxFh9izqAbKt2XzW/p3FW
sRjc4DMXbtQyLbYLuXw8XEa2ELJvI2oIVOXeNjoCNgA3kk2Phrhle8Qtcr3upQEI/wtp1VHb3YO8
815CpIkeEVU4VzssYASzKtlmMd0vCFiTU2Hd07VqhF+Qiem+IraOycdv5MgrXy1IPa6h+TL7XKMv
47obPVy8hOYGS5Mfj+cJklTkbANtgfrmqAF/oLVlBfo1BEfClu9Gn/dtKnTIcePLfsSLgm3r43XE
cMHFv3coEoW7b+LURyUAsSVd/9FW4QdOy13esbxPQTxnH9ppY8WAq6wupZigLTTENa+pO06ljozP
bCpOi2SxOUjWm904YBQUmARUIsj9qXzXdZotipBVXAcU/sVuBX+kW24yAULW6ztrwKZGC9WVsliO
tAY/pIWh8qltyyBvaKRpLY0vCC9cBViVvKUTu9QU4jAHZcjsuCKKUlQBk+F9twz3Fp8qCVYD5b5z
+6BPu65nDAEccOPHnJE1brBdy8H+XQXq9X+v/xYiuILVgfIes9xfM45qLwcKvBwTFsT/rD5xUeIg
kw9dhDh2yhDy7tSlaa7DSmMdC8BTdxI2y8IpLA7F1npfVjUMypexN8nGT/rIVkNgg1YDye5UvkOD
onYfTmAjo33HpOFtewrVyLI2jO1NmH4uCGjej5NIHo59LKWu7ER4zvMKRp/eZ+e926ZWVbAtLRtO
dSyy4VzhYCuBoMbQHzbsbi3YzF99ADIVKUsFpZRAqV7gHJ668/kma4mqq1XEHQDqa9mcCiXiBSUc
uiplpJJZyE8/yV3e62VGmjjXGNqR+7Nmes90zEgmk+IeGoUrUEPgMJg+rXqXEYaFeUjYHnkj8hKt
Vu/hOUitQv8q7HDFpMb8H3ZYXVDaSpLSCNJE/G+4WKnmW+A0VyHvM6jBXZH1Ky0mJC5mRr7yZTW1
rVFHbC5nfAi/jQybnlAodzcnA9BHVNbQB6nTs0THnf90xxYyrdN4Zoj9yoMfQvCfYQdpVPlSJj/6
MPjkWPS+Buo0uNu4VPvFDNqORr+o8zQAUBc0rx5C1yRkVHWDsDbMSQMt/59uw18pbhWKDHt9AEXk
KAQSeWuEWCJth9NT97OB8c8hiqJhtEU4pQowdCzKa8iUMx8ZGYa95lG4O0jifOIlrNJkKqTVgi7B
CZgookWXx1QDTLvKLfP+dx3WKXFMkSbaYcUun0wc8Y3ZtKsQtASqRXThUTT0U8EcNoYbzQ5kH1Zl
hl5wn/sdUPDfAP+/PkfdOTo7qc00Qi9aBCDOsohZ2sSkSM1U4avbs+X5W4dOsyIz/vq7pHRg4Cov
JSgJG3dXumVxaqm2RrC8KJLxDa4DBkPmd4cMZHcsOu9L0OuhIW1X5o4yWTYYSI3OgN43HASLeU1Q
HCjkzlVHH+Wu7y8gNEE9FCPl14BweRwDEfwb5/Hs5HbtQgHROIwXZN+CCH7R/JccR7ZhfG46FsCn
y6UhzcVi5wNv0s1blQ88dHYUphr3gIJ8XrEOlCJqWvKepDroa3DXqFxuMhMWgpbytcKI9bJspQjB
SGRI7JYVbvQHZPL64n0vlU5UqmmhpgePG8eitoOtgnT2OBr56qGzAyLvvd85L3JQd13vvdzr/OBF
lBVXNM9xhWHjH0BnKXrBIKxS95JlYysWPxLk1ZIAg45E4i8kYx92zuWDpBaEkq7SOsBhyo/1ynq7
YHwuV0qqDoMu/q/hV8d4zweo8St2m/B1SPSCpH5GmCYDm2LKmH0urRUqTjIHWZwzOnLxZ8s2rFeE
YL03mpGGVJUX5RbJYxEfooozhcm8t/ffnh5pTmVa1kRqj8kLDPmNkZoLbtg/+6H8B96s8q2LYmfY
L8eo3cw44sTQ+lxhgQ80jMXS+VUvxUdreN28MzFkTJTcsCs0F4znI2pq1qlg0IeTf4HeuzqgfT+4
HVeyErjiX8cAFcb2PKZCPEJ2WixDuioghBkZSwNXSlR0EK77caICzGBhWt5359Bbv0QQhX8kZIiZ
9nRCDZmulOM+I7bVG8jop5v3SX8WXfTbkQQqZ16feyzQmMueAFoSidPNhff7Xyd4XzwduSOeL33S
PGoFaU3F+8luDgm9WwyYhZJkwtAnIRiQM36gM7M1Yg/4rQ95yhNrgvAFstfdS664q3WNXsfRFLeT
ajcNUsbuLOLawyWqCB7W3twEgZciJ618kcigw2lBzon1pkTjB964INkmQB+pWURjHxGxj0bCwI+D
1RlyhK9g7NUdszd9ojYDomtS2t+wOJPzEntIehdGhA2IBHlSFaoOrlO+R1PDrOSaN8GOcAsZDaYN
XlCbREXkRq8NHcOqa+85t1rGdPlk8aInKM98WnP0E9hXbFXtFS2NddyXshzdXx+ePHT8OMz09pQs
2jIUR5dyWxn6Zd/IPFWOgN1IifleqNvk/TpTCOK8STzxjX51GIplLSomUcp9yrUSGWVXLlYnaNzQ
M478J2zXgMTMAf00Th4YbPn2ncaK5WG2hSmS6ytZfiS3IR1kRw==
`protect end_protected
