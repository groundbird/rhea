`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GVR3tpUqP1D9tNDew5iD61F86qRypPsSkj5QVYxZA/F1uzAofhHK1aXv0F6vKNSsS6JPghF88I1H
rM1nqgXQww==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mmm1Pq3qArHf/jIhaCq6mqdek4tqRoxjIXwmX/UwoGHa0kgpqw9xmrl1KZCzzLLJydmwjSDgTFlV
mr589U9bh+EmmLK9uqWO/NVl3pja8a8GEocGg4gm+VJMOskyZ2EnWaHVrG6IUp/EQzrlM0FDQbu2
EZq/a05s7D8woIGR3HM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jD5U6zH8NXmm+3dRqg3oV5ujJMbmxbS2TpKG8Z4Pqp2UnDZ4+V2I5JI2pz9X36W3TI7rI/jZSsDT
V6eAewp+Z9ggYdBGMLrp3vS/4hY+An/aTBrZAX2bt7Q1iDIR5cbNaqzn+NSKYGRjzzx3uFlpdRkM
FCqyqM5RKYzUJqsR05Nz23j1McD02w71bAqQID33x+z4NzPlz0PG0w7hQcxGYUEPw1ZuIxAXQchm
FimO7dOAtsKoY7WmmGlZAEtta2h1IvtCdqnm2oq/gVSOjgPF4FwJuRwD9/Z3EUHnOqresSk18k8q
nO3FuUThLWCb1Yrbc/+nCHDlDDi0s6eYVQ37/w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Wi6cKNdp3k34AFvSYKkcflCpfKrpDHlpa74x8+mfVoq1S1+O3D+wL3HL156n26x56Wc3MmsQ1WoT
M3+k5XRVb51ydqZ6LUEySwxE7y/dTTYuYkUm0qgS6T+e36P1LQId/LYZhr+aA13PyJNWFlWqxNY8
U0To7NHmCqx/UDwcrcg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aPYILVcRPSju9bzFnAdELiQgmB1nypc6O+VPeNMM/iWt4nceR+1cl1DvGV2rukOC7tegbT4g9NRa
+jXFqyE+jdj0NLejps13j1RpuR78w5WER8LhNHlZChP9bYZeraPUfLuQp6nfQ1iAuB1ChKCW5YKL
yROQmn/uQMh+Uwdvz8uO9gSj2M8xjNpkkkYqGDISnej7Jtnty4fm7zZ82E088kee2doQc9W4DvEj
8T9IbPQLyAQULvB3cIZHVBhxH4WJaoVzfo+3Gj6qlpNR6uL9HFIk9VYCKJhL53buJ2rLPiweOPgm
Wf4akPPkSo5tphBvbcKEDKNOLxq8HrfHpcY7WQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1540512)
`protect data_block
X40EzPOy0DTCJSMgwe8juTw2MjNjeFdyJVsRJnwB3KZcMz64cxIRp6XoZlt6CkPXlIAD32LDZLGg
skybSz7tQMcUmWwcZsSpRKqphxtFZsmS8egOS31+k2j2Z7W99FXEdLIBgFwTnRXaY5Os48d//Wy7
o8WIldnrLE5dFSfolNIkt9/HVlYS+2ks7kU2nfhAxIuXpWGdmNqpNexr8AyNTlqz42txVPnlu8rs
vJ6Nkp+jct9WaSmYEsmtaFFNzbP77LhPEqUaB36PFoR7lAxOrfu33o1j/W7Z62BuInDEbIN3DfnM
p7xb6+0OXJsbl0sX3UjteI0jvhrQ+XFiZKOkQDHZHYJ6bY5fm+L3RurPQnq0UbMZbHhy6SP3UY2M
/qKwmOibaxMbq2gx5evN6sv0TKKpnaHw2Km6OxxDgiTB9QCC1hkRtCSsj+N7cCnbQZNmCLXs/zte
UWJQHxjYRXsALOmnvZ4Vu8CcMdhUtHRkIVawPStmbpeiMEPqX4HmqVCZSqxo450nWb4wqjqLTpY3
Gr/yER8bjDp2FDYJ18mcMuv4xwzoqRJZK1OPv6GWzqC4ZF6mBUFvhWNriR4zQiS5T1ucimnlTc6h
/F2yys4uSK1lBqpt9OYWklj7FM+4gzSFb+TsZSrACSjWYu8XV8ApdImA/Tqqxwewzr3wG8EaaK2g
ApPLLhpbgR15ChJ+uyRE9Dk67L2B2i6lLOZUX4pISVLL2qYEkMR03q7uLMTmu9i4XFILHxBc3S90
Z3CrANzJPcVscxEmmyI2q8s8CBSQmDnaiOuuqaiyA2WJroxEKePon86GnPCZuAX8hXbEqbw/Hcxy
aY1aU/GOiL+oFg2Ku0Q5QRJxSq7wgJggblGjQZyVeK25/zzLpkmt8mIQz8C8KiJ9YX/o+oEzTPpw
1mJdx+KzD9YrSlX70puRQiLisRWd4v+yjo/PgCtsECOTJBkU82OVlmSlg7rJF9Wf/lOtx4Cb6BEi
3w1VcEySkJnsynsRca759/3eRQxXm6PvSLL9UoHPOgWEPqo9VocGir4MXBQwE0Xfl20yaWLoQC0Y
fhfyp1sA+kFeBDLvRlbPSTEOOxzrycuSWk4+rpAKJnzRcAjnZBc5MFe9pWZ3O8PnxheENqExA7Nr
BAWrbahOMCg2vSgXG72L/YGv3cUIfJpn9DkclwavEmcD60uxIYjThB3XGLEr65TTPqzMVrW2IL6a
EyhmACbL2PLVHCaONsx6R8txQxM4LHJju6KG6mc9Am2L3uwWc9hWVcQcF5F0tob5lwqYtcIPP04J
0r4TrMlzhqu/BxZQKh7OAvAfwkta0GNgbIvGMwYoKiLuNTyR9NxDNXcZ4uXjCSVrAHKk/j6j2FiV
lvYJ/LU+UctlpxpgWV5uolagFyKxvU2ZSFNnjw8/7eHRvWfiIIlLy/Xc2DA7PLJLLjVkVPj21z0x
UTfhGb4t2jmqo+4QzR2OC3jcTGWPrU8kPTEgguWvTnrwCFtj72Rz7bxI+2NbgRMc9q9QMVXg2xd+
d8aLLSr/UhDp0QKvtmjGqmMBQiWGc7uYpWw/2vsbeOwr0H0js2dBwLBNvu+gxhoVYSmVncsj4sil
yeKRhw6vUCPjxIGqBPoC71L/a9z9LU/pHjW1AM+NrBAvsunqskcsxgg64vTR0qZP/EvmNrnOTDPy
93fvPbWIYz2ZaJh4bZowCUv5h9k/pnpIYDfXOK/M8oz3vCHUuk59niXpf5dqyugs82W4QV66GhXF
ZUfyEuSkTuFCrIGUzTiERGFXulnBM+mYJtV+jt5nuE6i9RQBBymQvnuxtf1P7objVs3iSPSZz3m6
MIOtZaWIvp4eTmZQ8ig9GgoOHzlAV/mbAYhTmLgAocnxnmARX1bj3Te4wNnqdQANu3783kvLq7XB
4ZflbVujpVK29OlDw4xKJllMXkSNo2Vuus35FO+WKSQALaBXS44JuX4IuaSFZ3rIN5WPREfXnsY8
vBkkzeR8Yfk2uNrS07/xhFrv6SOZxLw2BZ6gu5Z2lUbYgmxI86tz1oas8thdn96SLuAP7DGEdO+E
TTZcl2sKr35C59OP81ccPgir20PFUgp7Pa8o/NGCoNYd6Bajdxpv5Adw3MkABTUO93YJZg3ttddZ
Y5Ad/Iw0Xai6WMiAV7TRLY8d/rc69EGu2Xak5DnDIAHq0bPbbuioZKdlZX3rJnJv9Ziz6cAd4Jkp
W8ZZsT2FgnYF2vYqmLOlXKC6wIqGNdxIhG9+Q5faPljrRAl5mDUd2p4I+koScY3roERK1fDbeSWr
uD1BSAmcf5thi7RvyxPDgKaHpGHS7cVjHCYY2101mUq1a/9wPOVuZGceYN1TzHk9iY6/6tP5jqqu
968PA8NaAZVUuAI1JaXynVM60QJ2ddGz1MWM8L1S7zGsy8e8qwt/fzPfmfL46pjTmC13TajAyHAv
RinH0kdnqNc3KlPpr+p1BbTDpCD9LMqwA7uQ5GQNhxp9ryz99/4+WMhPZwjzv1AAcmfHOPveWo0r
h35rXj4MXyKEuCtHld+4shCjydU+GXL68uo8apDyqO4gY8jrsBiYZtDhWuwqrV5okgpl1NqloWHw
zgD26gNfUMfVR9TYTHpom5+SICxwW0zif10yee+cw1SQOEU8lZI9/LngnrBx/kB4NWn1RBcEuh9b
g1yI2JNm5i2LnbJ1ck7CVEknwuOKVmEzc+99vd0X/NzGDzu9RZCXqUWyaThPCO3IVfvysLgAs5iA
yTCvqiOOS4utPncqygXQ2MLaNz2eMziL+AvX6xRp4VDbBRzFYs+KmX7cSEd1+A5zrI1aJvDFQ0Mt
tYu8EPEgXPwDDgeXl8Lqc+jyq263l1RfJLiMmSB7Io9Nb9dEO5WkQvmAJAGyB7CQmBau0HG1zDJL
ASNOZtRtCHLfk0YQU6tGLA7L8h/lt5lGxkrWk/JlMi0ZRyHWGmPsRrtqrSVf8ia1kAPtoS3mdsob
cXF0hXpkcpUndKz7V6WN81abnxEsFdb7+rWdTqny9M5hzllA8P3LvTS9GVvuU54Ssc02GGNEgCi+
EcRuGSCGx4QNUoBrAnW13oh8HB7ntZyy9YEQ0n37XXXBXTCo5R0gEt4jY1c5oinMnN5VnChZNioW
Ds+N/7vwqYNRA2qLQHo6MW69XjQL/WP40/BBXSi2xMgdeUkiw6JJ5BVjWKt6x/xb8zNFxg1p3Nar
8AlYI/vlXTGQYILPYMT4z8R2NblQngAk/i7Ig0LcQSfx+8CNAtT3xJyxGaYyoGn4rOtJGSIKnKsZ
G318aUr+3GF49dKBhUbprSwWYGHEUX0pPkD3+2BAX/1N+y+YB5bSH4cMHkiI8HW4p3OdRVWaRDzF
mwEydxQQIVqwHfKEoZL/859ptiMYaIrk/fmEX2ppoKLrazdfvFWQHg9iKNsp2NUpsxvjK8is0Jjf
omqMVdhKAdCHdTTO7MI0yrCUxTY86cT8Dyrz6Bmj5b3G90zGs3F7oTaJOyqxmOhRuNdzbmi1DS9G
TxkqqNrMfQZGKZfDWnO/xWnKqQJWH3PpGn+LZJN+hZQ8HQH2udSEZaJhmJNnd5Fb3qMUmC5tU7wI
rj9WouBznCDn4fNfnVEq87OszwRiWT2f6q6GM9DY0H3V/d4pBtjs12kXcbUgvTyzgO+/j+THiFVL
3TXG2VDTZWCybcYtDIIFC5qr24LDDmw3mDVHtqR7G7d2JjHhwsPwm2xGF7Ytnk5j2IFDwy0WmDDT
9yvP1d1/JqojVn8hQzyiXyeZbJAWBK5eFOj5j08sq3cJE7P9X/VjNDnUE2bD1ZWRV1KXVGR8gW1x
4x1NTudXWZLtLVGHXTv2og6xu/IQmLXf1a3KaaFcdm6rM51riTur4cChnwwQU81dmQAFLB9hLrvu
nYMvtUfXRkzhUjgqZzTm/S9uXZ+NSvuP1TurIkOyEJA95XqePGvT8QokaOE+KbypM49vCY88Vd0X
fG56mgn0pCBYAT+JRiI68K0YsI8G0um2gK46f/weXeL+Z3GrX4hJdvRt5VYtNhnAb6uRQ/XYHINC
6qTrspjkgr8k0FRWtBbGvinzbr/VXq5LimlCBjAUEk3OUgdOIx0beEEv0xpHvk+vT1GJpTzUW0lz
4dvSJuKgQi6VOicWlvpa9tkavpGPaAaNQvIcTmbVcVPfo1KUv5fM7GWgEEgAWwOuVNIwUc9sK/n2
WuZ1swSbg+0PrkU+JEu7kFcw4KnKeQFQeyrAuQWkVDHAfHMfuXNzOKBUNPLf0kOl5PsExhpvgSeH
9344Ceahqn71oxUliCh8qcgxm0iyp5uzFfzNaJ1XlqUd6+vlGbvpc7RKTYJjkIfqjsAL0tGw6hsF
SmwKTcJaV9umip0F06ZZTcDJtN8tmzFHLEPspwxFvDiYVcDgIuqoYxDxq0bWAAhDysc00q+mIZ1H
OyhqWCh1xP1Yq/syun/m9r1aOWzRtNBcRXhYZSLwgMmRbAp4EhxmY6dCa53jCWwJap2pN6dOkQtj
rV66rHiNDYoBqTZdskYsgL6xKVP7f3dthdPeJxXwgGUWy2woxjxa2fPslSbo83x25RtnrywSnk4T
fTjYTvdBfEz4nJ9uBNL6DadaAp5E9TBjsmRPhcvM0cuyapYH+wvdXG5HtW0l+J3Mk7OHcW1Yb72G
i8lmxVXXZYdKx6ZhSbl8vf45I5RYDziUPB7b6xnCzbeAyIRWwF4QnZJP+eNgT1Bp2V1uWMJ97HWo
Q6sHkmaExxlwqBZzfO1CQtbcs2X+9MdwLRwwice0rlgspTSzNOxz0q1p6UyAUPrJIexTntgHvj/B
Nd0t9pHSrKhCdFzI3NOx9GAuPTF0yEnqHqefTTHXs86HRIkl7A8eocPc6Nzfcscax4mQztaKzwMz
sqgveZhfk/CRcdQY5oRkpNv4Zar3vP64hEAAhDCoLWzjBEGtods8HazRAcDLHUfrsxePD86+DL0t
99RQMdu7nbHzlkO0DNPWo5JigHxCw4X3wG1m2EaaHnTsRWiqaH3JgSg+KB+WcMpt2pj+FLzbFylk
Ucd30h1s/z/aV6OXPOShO9bdXOl1U1yvma5H4QKkTauQoMeWphGxgkWNE/N8EIbPcB2tPhX/WUOi
1WFUQEWqOxuEtaWmxMjVW823Alzme8kb3ZQwVHRN/KxO9E9EaumbmdAsXsqJfV8DMRan7ZWIet1A
OQUmYvc5Vu1GsJjb4kTgFOcb75x0BPbQEvyVMJLTO3UNd6pkPBVBQWBXhI9LNDWafwtCQ4jg1wQy
U0Xo3UCFJCUEi/9P58CIvrdAx10TgPgoOpUILM8xxkUaDjC5M49IOeMzBHjO23QW2nqdj8J52bpl
byc9wpYAwfStcwR33aEeQgzk943cNkomxlWTJJkTBr75SpiBs6CBxdbRTpc5RD0LLXuNd0rFLzVu
oqQmAzw9Q7D5DD2uWuQ/0MK0pv3JqYebgQno2HkyxBqb/8eoMw2fKZa2YKZbPv6qa61NjWsRsNyC
HpYXGp/8ECsVbrMSPXFZCkYmUUf5ERZymoWMT6oCZ4XHpsfPSWic0E96PxC87/826XnPSnj4wKOB
AoLzCI9m2ggzzVxHxNXCBaSWJaP7bZVWRbsSRdlUZqhXzpSI+pnXqpwtNjlKsT5RwzJ7aOYmmFBx
NGgOZtoI9yk+tqq27RkbHIwzwjLLvACJ83DdKcP/ECODgTOQEdwArPF3+sn+YcroR+gY3CO6yAAt
GtKRioQsz/31IFrmEeHNP4OOvsYRhAlS1ahyeMi7RH0q4G2NgKBAo4ZapoQ2/4TnRLnBVqx4wKjR
6B3ji92r40qAy57hmwAOZxHGWRxzNOT2+Ep0g80/bue4eQqaB8u7D/HfiSU/cAt5itPtP6EtN870
+b9csD9VzmHanm8IarJnrdTi+8IdfJSb16UFqrY/g05/o8vZEEULC8+9FBmdXZdTfZ1WahxX3U68
68yGHFgWjPbCDdQa//mnazpVfOM/A9qCLTOUraKOFfeVnyTVGeIAGBbPWkCgq/TJXwzP3IKtzgsJ
Q2xpxdcmfLS43u+4SgkwcpYySmvadFiWmj1/8QW+B2JP6iblu5LJB48YKQ/U07yJzWT+7SL1Reyh
inshMpleQ0ikHxs6RuuYM5OPos3s4aN2pmTVlNBQm1bBBexi/kixNMDqxGT7xl6SeW+AB8cGEiMh
CIlwiKU98HJmHTM4DCZPtI4mzb3k7Z2V4802XbH1skiwwZZz/WcSk0lgJ34/oclLtkJvLZ6atg2w
T3wA+K7j+N/uZQ2uJg7SiXS8lUmtlNrXnehl0//c4gnpfeD2QA9B/a17iU1ZLHmp87VgzbXlk1aP
WmSlBl+I66oTko2G2upUZZUVTsT0QpxiwkJCYaCbtKNcdfmzwcP4ZBJT5+0QM5UkqQmXcHX3E9X1
3a/H+QveiOfNbm41CcaQgS7b3LLeyB+n9QxtvDKQ+zr6S4VyvtpKJHEM63kC1rgKgkbgSNNtlp5g
F5ScKNhEIJhBGcXbcSeuFfz8bTgpwYSRuR1kPo7HiXtpRv+AvXS4C41Uvo8lo89MiYzdkh5l2BZ4
orLwPCfMMR/AY1oyKn8LhcFtDF2G8osqPuqTqbvXN0sZxFEKLxatjAaKXFugJkmzrPiC3LxlNytj
+s0IJuYY8tdrB2I2J0rucHq9Ub6onu1Abt01Ah3hAQEeQsnAlw+Uu46rQmLrsYOT2nHE79hWjqrH
sCPcu0w5s8hjzrCH4mHagSL7MUmUnWZtdxS+USwAEcR6yLCKz3CFLviaKnAObWpJseQDAhGPyNSr
sOszG+Sg2b3JNKs293dXH0xZJ5s26SbTLUlgSCnRvkBYsQKn+5wmbQTXRMq6tFf0ZlbJzfjxkm7i
ufKB8yAHoNlbbnuqNEuhZWwcQWGa0wqt+ft+MNpyEaDx7WJKw2q8XaLQMBXI19G75UFCBb9iUVS7
zrSHpY/YH9vN5EZNHbJjLntnD/DWt20ynFkyBUNVLacwNHtFGCrkRDSxq7Zyi3qPZgCTQSoD7ch5
xuGQer5e57sDEc/nijhGtcwFQJtTg+7s6iVtNpjO2UMj1OXTcqwYRVc9eibpFIGYrmkvYpafzkIA
uFG0mTLhspq09OrLCtRkvrA3s/H1K1mTxG52OpPbcIvIYfbWyP7fmgym6x7x5KmClYN2c3wr/4RE
tyBqaGITJEr0nRUg7jSusnoh9viNJUEWNeCnVqDRfDyVO3CWjO+LFFf+keueLWnat3zmmGy3HIXb
7hux+eH2JiRE885Z95mQ+WKPK4q2FLFO6Ldkumh+XmMEq3nDiM/27Uv1eTG51QEcyE0wwuFmavEH
gLE181+jr4rrUSpuBOPQzkpXnDWLpmImkXR7tIE7NqTXZtgEgE8fWMyPQjTarisqgI4isTyt8TcB
Zv64p0XFoSdeYPmFW4P/mF8Cojar4fqrPefoAyu9dYsxdS5RtgGfoeR4SkExgVjScSDLdnPELeNR
eSQ+46k9OrMC9yf+7iVvPrfwWT0WuPXUKKJDtXQM9Icp7RBKG/XSk2juRsE/ol6dekDGQ68HVrb/
fWhcTaCxSCVCjvxLVGUy7HC1C7IKSpobeSDNNGTxIikGZP56gmoSB2GDrxMhrwQPf++Tam/QDx0v
hDVA5+ss/19lOIcFwG1U9TExujkMkRWjCGLbpOYoX3gQqZzPrmVdpNY9fFE4oRDdT9+Xv3AjkFG1
//UZvOTsvrjhIu6qQF+rXQZk4fpb0gskHlh5w0ls1fQV1gXxkwXuayK47jVylPzZS8q/W36qUxsK
NTCYhJah6BCOkDF98xNB17P/JI6yctP7B0l2ZM+qOBE6AhpsYy2UoVnIF3rrGMIzZBzPEiSeH774
YuMYuFrdgObuJ6ZaqqCOEn25zIJ606n5ixn50O+Ejh7HJUMwKTTtUZsOVRteNKerKw1m6BDIky1b
W5OQY84ldKANaVegC7ETaDPRpTpuaHNketjw+j0O3l+b5Q+/Y7dPZKoW6ELyCHRcl3OQUf/tDAia
MICGQfbgLrAoph3ev+uQNGoTd4vnC4RWMQDw/oZfZrJtJm1HOC45i9DZv8J+1OIgbtALvV8bSXEO
SFt2Z/jNLY9FR+L8I6xPyzqDRqY/yFqRQ9uYYJXv71OuON2LnEJwhhJjUwLFzR4u4feoQI59F95g
D7oY2QCZMYaNVvigmWAp6SQ59Cv5XmWs5CfvgYsTgDtyGeuAFFuJ/pj6ujtsY8mRVtLvxhdZozCP
8gT18NCxmlEetxDjahd5/w+H6opAaR4a43JjPZ7atjRKTwCBu+k8TrSH9GI/L5CvYxstIWYmDIea
qehgizLgvvGyzKaeqO6gh/uHSZjm5N7GB1uaetYcfTs1FTzX30AVG0zo520ag3t6gtKJMfPWWGlX
71efGoM6dQgduk9zw4vZHKPmtatFTUzYFTPsPEB3Ekpn0HfY/8MVdnV5EU9t5G8WCYhaS/FB1zUo
9QoyhZ0u1E8tghB7aXnmtw7uQQfbyGBJU8lp3V0awHkNDc3LgvFpG4Ncikfnj3w00JN7qYtdOlFF
bfh5XK2u824k5kBWTdLb7obQcr+DHYFkG/ALizCg/yT6Z39qGzs3Kx2+AKMYofQyV5p1piL8zky5
8xJyWTuEObMmEb2F+BIrGycbaXmZaJW6w0PQdNcyaUxrwEvOJfYOXXhd7bSdGTh0siO34Xo0lhnP
a5OFu0CQ3oSQVrEfwM+Q9oPXyfOEc4QQhGOzS1fRkaZaOX9OVlglIY2kNRT1JmZtt7ydk6J7YZcs
d2gj4og0uhjdu3JToM9UJAqfoyykdH9vYCjL1Wg/i00P+UBogCRlKhFZI0xvfGmHO18Uxp3VNawS
HKI8na0mvroAzpd8C01esmEXeLLevlm+hVeI4ZWsjOCVgI4VXOyxg5Olxxn3E69+aqlh3XIpCNov
LuRGqRh8h9mmkDkCx0LhUuZibxw0RXtQssoGFQCOAv7kLm17VFZ1VhWs2RiEC3H6TDrI3v+oegvi
7SHdohoxv5QRC+Z00qXd3QSY3WmnaEsGocbwXot80jpTf/z9apQ5FQIsltvknAlP8p9OwfpKT/vs
4izTftPd2thqfHew4G8MCu2vqJXamHleeJ2IReELTRtYgHe4rxQj7vA3+CjewgTxAieuDakTRN7M
O1TVfhHTSsSIAbOBCAHNSicqcqBorvdc8E3mNEThOzDC7VZdyg+fXZyKyeXWdmtmYS4Mp8mRP5Jw
l2UzD3H+5f2F19ROY85NFYMH9bVGeyD/hNwtb2GMskafIp6B+bszeATSpTariQfE2f5XNJjbIDUa
C/ZfTW0laV33ve4b+7q30b4NXhFWB9zUMcA5+v4j6a8IM7UaQp7KwHHsHKf8OZXqadb3FDeFna0l
CebfW3rzV91LwBo9zt3lgVb4PbDxc8a88bBU3UAZyJs99zB8LPAq8tbu6tVYqv/IeCVYyvY/kzD3
Dpr+ljq3yG76xdvVeaoelArUiCQxYs7fRMw4btN/U1QnsaWzzs90Paua2VCaDETgQW3l4N7lIZLL
Isx3SEIJETLDTg5ARu4zHvy66hywRDKf/Av5Cu3N7pQyxAXME9afI7S1FzKTSdp6oCJi9IJozbAY
rZNjDrZlXycYfkHBzmU+ghMxG2y7n+V2+8Kvfw2XEkmFqiVYz2c6ZdKugKG5FuaAOX95Xv3jOveT
NWcrY/+Ix+k4zQ2Bh9ye3zPyKII80HcHDrtVYDcNn4CpGTkQTIeQOr6etLhidH8YrQ5BuuMOtFsm
lOi8hDie2foXl9KFK2x/66q5c71J+K0bWQMmqCj+w2hrPAyjsTKq8N7HrQ3ljLy5Fn9XWcM/D/d1
KMHHuXjLSw4Qp0qHpGfysPlSxuPk6wTSVKu7h/yiKTgUs0AjxsK/YSudUgnaZF3V4M6qkjjPg/f9
udSRYYGAuo2XKan5GY2BaJpMsDe/BzxT7ZIhheLQ32pHYfDbZRf33OBdIKOoB3aCpaYt8qFihaOr
0C1qOKhLXQzVnMemre5V5iOvVOUmS0MAxfQnmwS/0vfey7Njs4LkGgLkKMmInLciOHzoAu+vg7gr
oIjzqoqas2bWJyjFkU33Ccx3NCUfQCkRwsHVRmKqj7AwqCQeRqQn4hvym3GsnTndWRG6oi+y14fz
IRmX58/XPC2yEYHPgKZc37Mj8/YvrAD6gxrCfL/oDX0mjJL29TwqpNEJhW7yEeVudlO4uGFpEbSX
10h45CWrnn0uaTh/f+CF6sLKFXET/X/spKMEFZ2SDsOWaaRuVqLhdr9IoKUPjdfz3egoA6x6fnGr
Epd2NbD/CEWR3voKgyD/VXlKPO2lPQTevoiFG03fUF1/DmqFul/O7/CxuJ3WEJs4lCpltN93I44O
zo1O/rQD8eQX2+7rJ/XH6LEgBFm6ozSwnDcTkH15Ire7dP6p5yLpLtK5njUJ1fc5fRJFEZZl/ziI
jq7AOqvG4BdLr7sfgTBIaTQhfyGYLpfdl4RjqMQJMnuHptp4rZoIO4rbxfZ2OlG9y+HmExu0muWx
a5tDcnZNkvvXR+xdIjKPSF4lgyLp8N0kXRfcWQf19MI05MsvY8eyeggkxzlYr4/dwOsiP7jcuHYx
4pAHmE4i70Ma3hyBE0EyMx1l6I7N93joyeUg1uHxGVAVopIFuQp9biFzhcLynAVw3svELcfpWA53
hl9RuiVOyaNAt8/CHYzdnI1Oiuk9isVJG6X5xBl03anIN9S5hZzOPuW6zzj83sujieM+OQf9iNPV
MaLc7/AOIylMNN1zCOGbUClxfwX+caOuTewTGJL+wX5c933gEWN4NSTsgCFRNZzAW6wxXspLqCxl
mDNNWL86n22lMTo1OwfWxiUSOdMijIcTMV+/FYX5M6HjKf+j9j39TK2ZqXPNEZ0yfKaxYWJG4mOj
c6p2/AKHMtTnu1nVWMwzOC5K3AtiDAa5f3m6lkTTba76SMWk0pRw+kQRXi1sunXZeYmNEzXTvBMR
bjbUkjgdNexXckAD3vbPd1avb+TGu7k2eGdLa1xZIYwEzWkkbcUVj7d/8vNHM/itRIk9r43/L+p6
L1wKiyBJFNmzzIOB49cHVXRnmSN5MsyXeJEkGplNMytgs2EKSTJO4NOgnujZVyID996ky2vqhiCJ
6EiZoNJXHW2BeYx56JIEuiofnqHq/ypDgcgjszm5JpZnlbN+1yej885zzfQU3uiOmAqHWMJYEYk4
hu9tB7a6tUUXrKCrx8tuJOUNaLxgnzsvrN3N0rwLzKsYnbeN4MIziVTXFqssZvXZNXtgGRSN/K8B
Ej4kXYNMPBoOkd8e/w0MBi2sa197DjtGd1vdr/9U4DmdFJVzXNE0pASMe8vsl0tZR/weFPhAt3Kh
3OqL165ICy931EPDj/GcUZjVZuQMkK+0Qhk0OS45lCtv9trykd6tOOEB9eTLCeNarZBfavJmB9sa
llbGuIoBb2/GcBOQTM+TSf/ZJjJ+SuS+LBxeEvN97HQZpYQI+yxasEkwYrV/mmjzDZJ3Ie3/kgHh
ukMwfhYUSQ/ruzpcA3gMGHAAEIQ3aukh6oWJ69vS8w8nIVPec5bMT/eJ87DOhjOtyZ3UYx7WUeF5
nIMzpAvQ6IwakuOUb+CeiwX6matgiEw2qi0oGZkvbmTQhyndR0BNnca4hStdxN3KdjF+HHlAVEbD
Cbsb0YD4ICY8WXX4mh1Oh4vgqq/5kDBG6yXPb6/uuLbBd9VJFLcTrCjYzWLgZ/RzzfHqe5hBJ5M7
cM+fdlNYpcYbQytc1SLCNLwzkH+MYzDr/Nzcmln5QzWn2nLLqyU5lh8zfuP5x41S5HTvEqJEOZnp
xvCx/fgpL2nK/tWlDk1/BXpB0TJxxH+jcBekEsXG9kO4/YY5GQON3H4QNgQiGqU2EG4lyKwdY8LR
60XUri6DkcDjaPRDU+Hw9wpNzy7nVUxuQBJzxTqqiRG68WOq2mtYenM+fs9E93QA1h7kmmgokTcN
zYQCE9LeeU4WWQIN5TAuZiBLQkr78H5SWEkvyGwk7rSYdeb2fwdeMK/VFukyq9CZChw9FP5VCyg8
HnCuWAwMuvIDRDrvj8fF8cPbqI7eGJa3uxd/oGikbPN09IbrL1ccSCPUfKB70nxhR8D6A1saOya6
zTkrT1shr5Iztu4GOzAZo6u+1QYZq9SGB7iyp5b16dquctrcfy1pXDm39A4CCxuJROADH2eOxSum
6ygP5i+lKeFAz9mYnBJEraeP1BQX+bwVPygweO9YdFDtv4JUpCKKyaMx8fi3w0msl/TCdmCHmxqO
welKLAji/BfLgsN+SxfmyCh+lGVtutpuahNJrJbz51DJd1xhyHFgW3+C9y5unVWXpBk+kt25HLba
GMQugpJedQTWQs262Ql5GmjyKbF8nvjBA1oiA9kDe4D/sNW9U+QMLxe6cFuf2rqztzRlV4/Utt2o
vnEihmU/OnFpUpPCxJmaaxRtOMRcjTsX6E1fIhsWAoKbO1dm3/mMKzIRdcd/sTP+L3w0iFp7V85C
JD8Sp/7dVK0c/ty+W9qW2/uxpPks2EJ/Z+yf1bEojgqmpGUWzxjxUcv/1ntwoB+n4fTOsaeAe9MB
3xs6PpQJJQ9KhjLL87IjBHZXNZfWUCoE4w/MocjcuVCu5yiYd/VHIHVryNMcDPI9rp/WqmNt5/Qa
AvUT4iudqc2x7/Q36ke4PxbYeJMaMXINC9/10uuo9F6FRHKEQEYArKyL8ncC3wKkt5VTyTkVy1fg
Bkwri4kfzXClpeAYoKW6HG266mYXhbOJ11qb3LYagIAzFgck10rqVO1u6UJitBefeZGSj8pAR4tI
tGMCbnV68KxTPJXrn1nTGsXMsEc7kYwObkf2siwrW0cuRW4Drn4uXN1q5kpbYrNRM57fzirqOuCd
hY8INIVXYldxJe7701xmqDp5nycV8fLXBVbyWvI/Xv2WdDbm2d9MmcKuVUnP3hvW7Q2qBrXBpJi/
fe5yHPhHPM1nX9I4nfg+uq19Oc+vFGIHNe4HRwGdEca+A27xq9IzxbFSNyeWtnyOY2EUhJA/Q9vs
KF12JWy1J6jdMLfI2WdZ3BF8YY96MsUZ/A21CStetQy2B8fPPeLFrJ+V7GESJiD2lRFOnmOkjJON
VWsM1ZfqVKOg+leY1efvyCALEqNowijrAUwZTTjHXmlgG6ad5LaUR+4W/wU+8Lzt0dua+ALSAZYA
GM6iO8k1gD+LVt4gpNUfHbcRJqZpWvjbg2F8AEufyQ/yBfY5TJH5ZRJ5//8Oa8EqQWNm7rYKhSN3
GtZQqi0vwpEjoZ+ICsctKKYcCJWkPpma238nlXlPzUwXO/rujR2Z39YnToU+t6iA+QYfonLJV9y0
+IPsQC2N2351TiFLr9UU+nsuDSWop4YLjD9cvvl1iFi6UjSyXWC8bQUK1VbVbaTi8wCru/kjr47w
a3qb0VY8l9tXM+8x8hVAIV/aBEjXb36mckdSU20CsawItvO8KwOGS6MoWkXeknpbYlrcQckYyG6p
YreX5/ix/z+x69sZK4KODVmzmXU55PF8dsx+WQhKcqe6NSFjNbTUMJl8qQxFsjjztKWMPdmRQToN
eqMZg+cfsflzmZJb9ACjIIqbJWn9ti7zJPL7FA9ZPM/j5QGANc7d+FYKFlUHSrciyrAwABjyATiP
NfjurmVKGccajL/N+fxDEii78tRde1yrK7fiDnBDpT1WYwK8xKrMnT4jTEG2Ct2IYV9MwJVFcNgy
HryxxH+aNyZM+s3YJ9DyqWPDW/SSXZTjfj8iZzhQ4cKMWCoAU686msk31uHs/PFHW46jntYlCQfv
xsBW3TpUST52ItmipMxu+tTRa0MKVIb+4gFUYwLwIWHas+Jv/Zu4rcvr3NwalXBBpkNm5XYSyuKz
U3QfQLHWbE32EYbqoFkZF4lkVTXfYmPSzWWumwUnertZEJEB296Ou/cYjfBKgTzFmT75D3MQNm3p
26p6Bi9GGLlpcf/QlykeX5WxSdbJCsVWS7hP3dTbsSrybrKcQdrkJrfqIWvfdU1809cRjAUVhrag
rVSJ/bQBfL3oSms+ErJL6OQsRhxPL3poJhFn7DEteXXVn+35dJrJxMlCSl6TwvHZybsVOJpK8aMX
n7Q+219koQ+I7nLZtNK1Ze7S1ZtpbZVYwFLyxyYQS9RKjiFnaKgFaUMR1+q5fggJ24mFktUY9PMr
AT46DgGRUhoumKtaeIUN6LSkA7ooVcnmIdEaYFTW24SrRbmqbSKioXWQpCHcB82Gy7R78tTuWFre
sdh20sNcuRH6kq0Yva2+mzOqc/iCoIX3a9OjaTMqSfzJMNpJ8jjxjwAyKf3B08zb7c4Qk5P3txWn
1MKYgvlUIJwiA5Ih9xSZHEp5JEjiCnSPnXxRV6qb/dnJQk9UY7wptRFM1vTaTJo/tk4FKzN1jevj
isQJyubbpJVwBJ23hn9CBcsSgQqgx1UAjMtvPs1rLLG4/KlVGb42j5EPED6J1ZA5KJSu1f1m/z1j
YXooK+DtIhBZ0t4DRkSzYk2+/vL1ohoO6CMTJCpl42ES+kc9FQCufSrn9EaGLBhbWzptNNkRTrzt
JuDL7mZSOxjPqiiEJPLw0dkDtGDqJqNgMGkPM8GULOzlzByhOJVOw8g2OxuFEWlmzi4RL0Nc1Fmi
kYSxezDaDxjbVSWF5WNyAbADpVAMT04QesWJ01KXB+CQql+xg22/zgJlqq7VnlOR4H/YHDNexp8g
6+4tBLTXnjtF1NowX7zaGjI2Vg9C2dravFPrUchy7H7NuOCsol3psvDhV03bl8rhh6x9jrDPg5HW
Oik3e7CPnEVcRDOf4U5ZggZvE3vpEcbJKxw/u4edmlBYMsQ8KUXRLHGlMv68SHYG8RlModffepcJ
3whYRduSgBeSwqFQ/kPNYYuaYFK3tw30ls87X4lDU74EnJBV7OaptMRf0tY2Uj86zlE6qLpGstrJ
ojIDWXUpGak+MVBp70L7f6bGygL9RrTtM9KMZo/11timbvbmp1pLf/GoLNeu8rz0QSrUY3yvDC/A
DVZP4aoQKxPOXYcobrOCFLa3ZJpjWi1c3zSJYjygAmoZBHiRQkgan0FPeJ2n3SeTqrBkKmt/jb58
Kl7ujwb6mF1LjM9QvjctCd6pLCCMIoVVZNd/P4pdQFBViY1A//hhFF4cIwSzdOBJIXiDqrTxjZQU
/9jfIoHdAcVUq33L1IoPxZslcNez9gNovCqfD74ycuv0yAfOX1tmTv1Z6V8haq6GRe20BHG+v0rS
A4ytty1++3YrhiBXRETJGejO4iXpboBFMc6fTxHMmjBerkgZZR4eisBVVzvHilRfMGkDLdrU2BaZ
5aRwS3gcOywOOp0C10htkz9wHanToLMlhUGQBZCln4TNPmUQA+ZBi4yir15syo0ikW4tPh6Hg6zU
Cn0Da9bblbSuGSpboXo7paS3gXQokhX00PBlYzacgXhGnFfJnWslMOkkCj1qBNpQeZX2E9i1+ltJ
MexDwO43xXadkWeKxq3Z6vKhPF3ah6qjHKes178CsvLsU5op5g+0NRnS1Xr9g0qs4gM7kL93OUiE
PiSQxWs4zQL1vo4xoyf/I6wW66XFYdaGboynheNr8o1rxn/WKDCPEww964CWd1hIFacvE1vwO+WV
dhsg+L7qIgQb+xjWw3TjaJbADNRM0QPXeli2CEmEJrqjl8+EH6NjBzdSmz3qc2E3GDJ+PmHq8D+h
Fc16TaaarMyAjp7WQ37L1xGnq4YkBVmcwWuqYnT00W64DI9AFfyCXGAFSP9+qz07tUX0+wAuEk26
Iy+SRU8e67FTeAZsGIoPH5YTZDhJ9o/3MknBHG3U0w0VABcCnYjdAbQwwbQi6ku4rRllvKzRZgcu
2erpdM2hSrBhjDsgqRpz8dtBIeRcRSQBmhI5VFTOtk8FkcCnRVWXWjq9DIzsFm4EPPKHzEjP7ADM
fvynEpm32xkNEH4H489O23jTLxDv24KOoWsC8o7eTOzJ7AtECdYJXo4tZADKBuhakrSFYkGFADIo
GWERlCEEAXjBIEyAmAXGvJoNvWgRr8YD1yiaT3FxmFK7G3Pd1BMid12HiYnjlviguUQm1fYcsFuO
tvrMNwmat2c9n+XYBob50A0cX1mzZ9t7z7ccWvfAQSZZr0LE/qSk9M0rCesaPA1zS8wOvU/uj3M8
UywBrOaes6kEpm4z4MI98WthkERVF92fR6qxNecZTqMf5pruk4A0z8wlT0gm8Eo48+N2+JXw1+jP
mGBPBwxwvi0ykvaqrV2yZ2g2Fnd5dA3lxfPGk8wyuWh3VZSeVjZOA81QsnRSsaN4OtGyFTaMqvWN
xU2nSnc0zH1yuJO7y8qK+EWwazEjwnyWZvEr2tG45GdCqz7Zd8UP6/4poonZNLl2GoyM9+rCkA2D
ljUTi/r5SAOo+pi7eAVzKyDqfR3HYB4Ih4UQQHMBRHMBA1g1TAwIsGbWPYcYFX9xnvZPLoqtqCrh
Orbtb7OIrn/gCJWXKFHZ6cc5JLueHzxfymxBIkEGOHGGsOWf4zF8EUQq1r/JM9WqSBqgZwHTIKOg
PTHKGFZzpWQLCJAQhIPyohsQt1nl90ZiyXi43ie5ZJspApgTjAZvMbir9CHa0/YNHOddNh7xF42p
wgtYBdCCc+cjpA4h0kdoBZE3cQqPKlHBDVvi6ieD351sepSFA2WqbXw8cIhJEvuA6zoK+agZ23d9
/6ksjc/MrDEYtqXCEuDCgt1Ugw6w0ViFLxcrSS5B4royU2dR4F8IKOQiprOnw7spsIdNoZfyQgtc
xLSuZVb1i3BIE9/nT9Hp6yNXsMhD7j+pNKRLxWlLbvwvsmJJrdIzEh0LUrDnxKOf4LZySEsEII0z
z0NAGgU0cOVVSmYcs/NtBGzeu9ChP6s+6KgFzAfd3i2cJBmqGopYIbakKTmHYze+oEA3OwyN79G5
25efgRC9ZzJtUaSqFcw8+uW15UmU6slli2M0jyW7mY+Y2cyhRhg8WRB1+yfF6A/lHHM13xCGXKde
8FVDIhhRJ0xCXij7mODrrBEbm43b+zN6/gsXbCtp6eMAv+yOV2rtHd8zhZitDXffihT07zwBrbM/
+VAMc9kAGNiJpZEHXKBNWo6Le46o0ZRPLsTXJ1KMDK4UrN7C98biNQz8LUBhDhuSt5emFMF3Hm4u
xk1h2eYyNn8RxYI+HoU+y8RZOC+Ton4dpsPYkCEcJR8b34ftRaS3EAyVgi2/4sBIMTBlf32NmQf7
ERFiaQIdBE2damlA/8Xu74ZqZ7Si2gmVswyAfS6DNeK8bfA0qUidcjRVkiDlJl8JQk7cplb3EzLc
j9sfq6dgOL6ASla/BF8p6qgwWDamadEfVKUhsbhuxxH0wiLpdXq5w86XybzT694Sk5DyvgUXv09X
Uthhk30unlcZYOu0QYnsJjwnU5Loumhf7J40uGDaU3e2WDx54tZ2mQsjusznASW/+dwgp6pbUoTB
/wJrV/KOpNTT6RYHfBo3zga1LvC4ewTfE9V1+d+w1SqvJ6Bb2m3vx7fZIWXvi1dgT5ksQZxcVkog
CwwW2swJonuS2lu47yAD3vS9hvNAvv4PJHKGcjLH6sj9Za0ULSu4qER2scQ0n1+caijBgQZxOjvs
4HUUPx0x/lFMmFT5u3gc1fDWJz7rfqKEFHHOlxH9nelfZH4ICU1ZkV6RPbtOg4J+BLOgD/L+LKx+
x9OMfeGUn20Cu2Mb7rxijeTE/Y7EREERbIlZmbb18cem7t/y44aKv54CKchtSK136TTHTV2bMOVb
lGlnzoCNEImAuzq9RiJQ5iBGJqvhGseQtj3O/MC+lPvN5bpHZUosIdnsrtqrdObOQtywx/ZCyp1/
tdYEnzPQrth/sbt6DibiNHe2CrWLzJwnyGchRtp6JC6Z2BdxyMFLVsqnUhZVrxMEzRPbHii6xKVc
289J8hnQTYTNDW5r1jp9gi9rT84tkufynww3NkCQuVbcYZPJg1vIwXRMrJiPqnMBoscI1e9wGmBH
Opp90fTKDvaK76KWZdrn9DLoR7iKF19WR1RithbYnvsMel+qmtGQSinEp2T4WQYxLcAcYefOVolV
8LiAQ6yuYRoOQRF5wb72L0zdcBngE8EU57YeyLCwJYwaGwKxM0gt5hDddRfiar5dHTtpgFuPjjJW
UAZfROzw3hw9Mdb/oqzS0hH8cOPhmm3f5pRC53/P2JYBqAQb4f0cwtAtzAv5Hg1xh2gkkkTL+pN3
73NFf1g6ozWjEPnVUPdep0WDiBN54/vjNtLAtEoAPxUf+f8qk/lPs3UD9E9SlCn1MzAf7kixApwh
LsdRVq0c14MV3+xeQ6z4/p0qV5ufC20nK9juRwWzzizurwHTMh+uaxUOfoBkG520vr1rGPoDqYt3
xM5HXKyguILlLhAs6H2aZrqu97nuk68tyHWciZLQj+FnzQRD08f6vxCBHvFLQjOOIkUabjH+Tdre
Bt4guYAz3VmII7ObgzAUUCQ5Zq6OgXeHULXtS1YQk4fWjzQMmg9ordH6C8mapxYoIyktyeC8e9LE
HZC5TYmx4NIrMkObb/80c/Cg0YBriySa/y7V8ObaTVQIM5TEnHaDyR+cLSc/hFmT9sH5fTbVY+P7
dbq5N5usWUKlY/K3+2M8lg2ci4rQZkbqiKbwEUlhKHvZVcCghzOiGBSW57qbvH7gp4NxopILyR1Y
dl6qRZiGwPpXCn5Yd36j8VbLfwdl2In/Fu37gfmfs1/ECF54UlZ1pmm5pUgKEhXFbIRUtQO1P4Sn
Fo7JAOPvCXnaRs2Pb+azUMw+7PmUdvOCcBj5qa2YvYgibM6QXC6yEF/HLdLDsry/elR/p/cQ0FTE
9coXW20R0SE0KklXM9O0Ue9V9nhdXxqjFcoYLJhVwa8qBBAn6NxWpx79dw9HADBO2seSUmWKffww
rMC4IfU2eTProXKYsVsLLq1U3j4WTfi3OQgwgbNBLgeoyVSv4tXSnjNlR9hKze9aCCgvHnZf3Rdp
8DrG0S6+HJiuBSQP7nzmUxSyz0qFLDSUmlR/Ba1j3wyAXwfQMilcVGyFy3xySHyus9xFmbTDeAxu
wRUl1R0rxtZo7eLJcZRweQK0N2zgfMBoag4mnid5vitdAqJFOfnKSEtf3jAjwmOKdRirJsaTRTpb
NPy9JQQ6J/LFzByS+d3Lrvb6Ijnu80fTW3U3H9nXHZefhAHqLHbQPbht4yGkce6LD7lKXx3qmfED
C8K76tb7IPpExE+EGQJ0dbEb5WmZEmZhaQlz8sLEm3s79NEITQJ92xPweUQ9/c5/3ZkZbIjIQuHk
1tvKu6SpqWQOO3UZXriKtSyO+hcqmpwWZI7v0CL9+HlzPImGayuQHlUd4+81o+1xFxkbUOoUSOrK
s9zEnXyaCsvpr2avdaQFyWYQ8nK4MG1pXQ1P+h9cJX+viLENqD2wqnUYR+KHlbvYP4TeMiVmNCon
tOFlrYMwQPwrO58VWAALQBYTsGUU1YHDuGQYCQO9xX5p4Gq+0+JxGik71Qs4z4BuQJn5uQoyRzt4
dPsX1EU+ngJ0mCyOa5VPYocXdKbrOmFc4zjdrZI+KD2lXzs/AM/WNvTq+kbZ9NuqXut+aZjNlfFl
0LKpHhqr3uhQRYU1Q5Ib5ZttkjQDkz2MxpaGvFF9fd/bmKIoOKEhNLJJ44bG/PkAIBP1mF+RECsj
/fvKQHY5fdpFY0HJy41ZmEzsXR5ZrXWlwnFvRPTWEdwOdtkengD+UaFn2nF1g6Vllz0NZ8m3svyz
RTP+YekYIoy+vzoccGFahYueoe4G71hpJuL0/tCwPP81KsHSO74hCUf7p5WVGyV9vr4LX3aNaKww
YDifPRmTVlqZNMsj2+xNBE29NivvMcWItvpwmR5G0Yxt7m3hvWH3GyIbN7NusiIO6NWN5r85/c8G
NrQzzJBI+CuE4xGq7DMlHbBjGoWEcv1CiNj0mDWrK8+YEw6vjlrvxj5++6FlVFH4PxVfSWuy/JJ4
V3nrAMExmHHgATU//GWfC4U4ZfRYJObvQJJdeS36Qr4sLTjP0w63QCJSP3nebgCo0lbKMvMbnWR4
/dzBh+p6c7tzBg4ToXiW2ovfaIs/kqNCHw1lfGTN5AlJ10ufp+LPy5Mdg4nw5L4XKZu/uwoi7A/t
zATUJX0ustAIG+KGsuqxAUamodVCN4fmInEnsLOwi3SlG1akLcTdm4mBcnuqtd8L0XAwze5+6iBs
Lryhpoxp2LIoTaJqler/1XVXmgcSRBl3QvADgHnwJ2ZxUYApkQN2r4QNzvrLWeJuG8kvnm/o5Yac
MgQhtPVnuixHP54bxkJDxLpgzuIqti07Zwwx98oA8p2M2BC1HZOeHd5KTB4uMuogWik/p1qB0d4H
SdVoSUo3BDwI4AdaL5F9q/tWDFPGay42hrGvgO9ofhw4T6zItj+e9rbW/cPJatcorZbygtMaGLPX
indt20JvEMlCx2BrUKF7gBAuvfwTW9iX1j403xxOrU4EQiOo1IObr21ta4PIv0BsIfRENDR+Nzy8
Gd+7clFgc2GyeS1gzRzKTg3QDy8VWHnx7Tb9KIsJaMbz1miudQqMgWotcF6kBOUjpmVEWE11Wd7N
TAIV75GxZBuBEOD9+uO9oix3WY14DgLu2hgmCXBMgZz3U5FwMdrxhSASVSBjOqGSKtMjuyIW72sc
NCTDKeZ6E0NyyEo+h8ulCaQFQ6UpZL9CIFARHkDWLDrmyT57bCnvIIYPCy/LlcelHc4YJvj/wEPA
Eg663SfaeIiEW2DJyNCGUl9aazmvrs5fkt5KabSzQrFpnrEjvT0ZVCDmFo7XEQkCTmrpEupWytyu
NyuzB4LzD1D+b6DbB0MRx8bPV2MONL6Df/8MhdOfT4AucZGRYH5YVr4inNzlkrh7Jj1yzolSgMbF
g3KxBJDcQk7cKxYsBS+SggXGnfjXTPj4DUWkB2GaaWSUJCaUb03cI7zwpwlSHdb14KPU2JwPzHVl
W/W4zZiQm/8Qm9OGiQMo7h0S/AUjulc8MI4ejLtdEBR8taEWSS4653EnORz1P7Nlow1ZSmGlFiy6
jOXZA3m3XLow5BJ7zlgdM9r9mOg1/egFQOp/dTND2nd5g0/7+/H0VIVs7ztg2b9VWsnyhwiMKDco
VGC6xFc4GwSpyQax5VmVeFFo0592mNXUJgmOek54+VPd0vljOw1ZBH2J3N8fW7OT8xVUKvcp9b2i
bx/oknXLk/BHFMKoYzYm1N2nw3UIH7SpeQaXS1zO46w8ObZSkoOUoWyGCmNTl70rite6GlEg4ooy
b96rlQJklfG87l0/1s26OKfA8o3v4lQS5OWn3yk21LrZONfY9WRmVVGMkvhQvAiPrKpXAJT5LwvP
TD4aY4ACv+ezwKLcK/CKvMD3OuBk/pg6kNNcVpNcrfNFNIkbEHGXKDntYWjfEToBayQrKayiipbt
u9p7WbiGqX1C43ysOb8WHG3SR+fRQLzECJyibayzqI0cKCt5EUAIwEnJy/0ORTWP+n+N56/x2v7D
ezNPk+CYNCtjhg4Bbhhgc8xUf55h2FgA0N8RGzAKBcbKMWTycwBaQZdIrf+lJ7LGwaTUB5QvYQRy
6wKRPu52nPR9i57DzYCbt7etW8WaZkbgVyEKUIRIs+822VwE6iZdrUBsxxgKBQgvYZDvX1Krnh8g
tmljOnII9Iyg7YwZlnc2RsDarr4fTuntizzHoMviu+XXZCY7sf/swjJQ54CfMbiQRTQGoqbFXzEy
8snukzr3q9IexEoaawdM6DlccpaoKpzmrqmN/AJ8PHrmy+jbfFB3Kovgt4bb2/XcOs2QLwgnRwfS
0zC/E+59ymEVvDZZEI6IejPs1YahvDGWRH4L5sn2B1OCFgB5NCrjG0mdbyYvvx2UEfTMfFAJ19Uw
MxvXUeOdNzI35DpPqQZVAUbS0FAYZ5pZcWyoqTpu331QqehQzZnCfZLCAN6dModgGQNz5ZVa7CMi
8YHZ/dfvAf3+IRE3HWGIpo/b5Dlf2HosIFJLnRmq92j8BpvL59lNWWQ8DjKmsHHy0kV+PjmIXqZS
+WpEJOQz8txeQj0noYhyp9wE5bdE4zt3XC9EqOjszLUZjd0IeIfa2dYsU+FPkLG6Ch8yGMLAyPtK
7zuV3Wo11F3zbhab6G2sd5S5cwXYTJEE2D428oYebOFGeR9ta88Y8KCOUyDrbbrt/xTrR9sVRhXn
M3aT9DAYO7ThNWm++6vT9OGc0UsT+WD8xZf4qBB4PLS9yF7dd0dwI9S8r1n2mZkQUE9ean9brsfu
oO1E133wpuG1hn5uP+LGuY8BUXppKcp3iW5rY/h3OUUoG+gPIko6HU5y/iqEXCkR5ARoWqRAuvFa
ESQ5eVbRlQhmWvb0XylVqYUpavsVwiQ7YBwW7tQ1pzR8tV01rIUpqPWmQ5TQgPIecxcG7P5ywUH0
61n/dGiqF7XsGluy3LjeI28K/+J2/6HXGHDNsF+/N0txbZJopzoC9eNghIZqTNctGpILL8X0v+S9
Nkwi0w4/wLE94uwQqvAV42zuvLRziriRcV11JB3KT/ndRlocWYqP+9VWxVkilPFXCdKMmMPeFfhf
4x1qDpdd7tJYLhvPOcMriQw4Ytr1qSB7bEeL6orJcF/zzOKGjrg+mUGR48UrehVrnc7eZ4L+vvuM
hzgk9L5ew9VUBTC1IS2P8+lBgmS6Y4jZy3RJisOrxwrFHgQFh9UDA/jMPTmrQepc/6yErpNAfhAP
I6wzK6lEe1VMJt2o8cpfmxO8jl4gcmlO7mvKsbEH2vr10CuV2uaAwxoMORWne8013cYWOcPvV3SB
gf4Or9AE+EmVY2iBA/xWGEJh/fRtQrMBLN8vMIBvFv41d0elEV/fb6g/u+UfQJhYHQPTLMxFj3Wq
aFsehqV6vvvuMfAZgHHnk53mhZCHXNNR/fHWInfsaWjwjyKHIiFvCU9H3ejt7GETOy2X9Zjr3K+p
p5VmMGPXD5Uh1D/fFB94lNMBnJFSIJ/uh+KGG5m6+i4YR25t1q9WMo4x+oAP9xSRxstkUTBI3UxS
FTRwkV+kqPfknimwX99lV9meCDcgLd2hyY6m2mOCD5uDVKjklSBCah7ienTjctIWDtqVHSqXP424
NXJz0SV47x1N+1ot5P7mWnBb+RWrnr1eSppOjNEg8uqC+6l/pWhnutyHlHAnr52WYe6JwboGz/3z
w6RnNO04k8VtwpXQcPpaJOjzXVm5AsvNYAVSyW3JTVtp1Eh5OXkLeeeETn1cLYctdpIPPzAwWak/
yyP3sqtFg2iMqxaWeF3DV+DsN+EJ3wpeqTHePG/8VnpnBpejTcbKfmxgIYq86iElEGyNi8gEsKA6
t7uEU4iOObShZj14j7V27zuN0fBobNZAosT4xKIUE1EJq4/Jgm89pyxu0jbPh/N3wiE7pZWQq0OS
uUF2KqeMYfbsUXyQIXF4uTls6nqeXY8ivMarJ2q+T9yE1p3di8VtV5InCfzlpbwpY3fOR1lWIQsF
mYgWbRftOvjk0j98ytQeqnU/Y27cMQD0y366AZiI9Q+UqPFe/cbI5gpGp3Z84l6UPBJ9+7X/CAQa
Us73o0t5b+8By0o3DWbuGnGrejbeXyVQJYH9b+kEuQHAqR5KgeYkQ34paXItj+NYW8NdUpWMOV7d
Qap3HyFyTJQc75RQET2uT2WuQ6gs5iO4LSntuXxwsZ/QsJuTOOgcdPlSLstktoHT3GQpTHeEwfky
FtvQaydpTBKUP7KeQGkGTAArNN70LgOgx6AYelPBDDsXnlwZbqJfSTyDNAx7+BWlksBMU1WMtmgv
SS7cFb/r3H4PSQVADTCTcCA4PSil5q5HbmRRZsHaZJt4JiQf9GSTqgQvQKyv6Lf794miA+vi63S9
r2Ym+zEPsH8VP+Rp1cQzz4WcRpJdSAyJmacVAy/zjWazeAsJ82fhlKTYDgjFiSilupFV4VmbcDAL
ciz/8/8ThzSA97bmhT6FanlC1H4q1t3Ch8MfgvhFy6CO0g6/tAfbICN4xKU6mRsStWCsB0SNmp3b
Xj0e0BMxm89V610Zfqupm98jMWL1/TXIA+Uyi48xlNV260vUKqChtiz5cZe6iFChh39lT4HEq+uo
qm6s3f2gz3zb9c3TJkWxuEQgFZS+/PsvK/IQkU8Vk/f9ERg6vYdJlfTrES0HqW3uAaqALL6XXm+t
xw3YKEuExuj9aPbOUqM/Sdzd9yNVhadadpIwOJn/09O0FS3Gd3/mUgFPeswrWyJw7/j4HP5Bn+Nx
AaohrNaD6sG39Ga6xYxB5RQrQ8GgXaM71T6MCm+t8y6zwpfdTLc/ooqXOx3BXiTCRIm4lHJWEuCv
YTnTBFP2o/uc/b8wFd4MRONkrJK7PTcxIHCYyxt8ybAP4DOaQtDLvAYJktpN+/bzKmpKX5dXekMu
fF776h39VwHVCdXMK+2sr43MUTw5EN0+7/n6fMQs6YRtEZONZ2tnLgE+4WRD9wAME7TN3ybr9mIp
Qh6m9R8llEKrqWuoQgXE9pdHg/LiPz9gp62kPrphTKlnGXUB9bnlPYyv7szt1sd7QeORwYaGdYbi
5TcYqWxkbjT82AT2rDIuVzKdEPG99PlMkTW/IExOXug9t1B3ifG6Hb12Xzzr9eYz1rhvT/qDrANg
aaHvAT1FMiV2XLH14RmFXUDXqnEELr3gTHct5JNOEEVeerL4rIR2G6d8AwjQhl8CpEudyd3aLhhl
gwYSvRgeU8uX9HR8Q9+/vJ50+DACiNgNOUkyaybMR/UMOzQI3sy81KyZhgogDw9WZHPfmKvrjqQJ
NHDOpQqTEacPBBmSRtiNdOJBBRbqeynXSDFYYVnd6LPobv7Jom8SlFwXIznQJBimf2cTRfc02LkJ
Ndm3J22PZjceeiLEWsD5XsogU8hPDucLzsfln2iaOwU1CjsEb3AjAbeVIZaD1I88Ea7Uh+boDDLu
1fTiT9o1nNh1x5xZuXtwFJfjCBfnnA9v3JX6rFqTRcDJRwaFGaj7rjsHh4Dngij0nKSSAqSZXEK4
ETRCyVRTVZpcud3DLt7VJpEwg7kvLm3n7gP7DKXS5pLo9+5G0R2K2sUTHofZJRPdclfE/tAOn+uS
4NwAvR5zkaWkFOdMRLWPvtC9aKA/EmWY88hr9P+VMfiyj3yUY3LP1r/Hykb5eK5DcSu5v8/QoFYH
gjdIQg4+H4DEFZXL4bgLKdisnOAxZz/TvBKJrPI6e7I4+apFU5aeu1F5doAUI7LZZb9mV08SSI0j
qJt8ZUZ5P3XVDYWqUIWv5cPiLq1ezoSzz/+/DaRWoavkzVhkKgUoa66oh9jepSYz14GKPBCyHrti
sit1qY7oWBkRGBEBK71J2Eb7abG0iHEuQBGacuJMMRDxPFRiDj8/X+bkCE1nbVrM3PGuM/KsgfEF
pJCZgOkp3YG7duH7Sp3nwfbTkWdPwZyXjnIWC8VtkYUN4UyriO3yLSedbmBPjZag8kXprWGdl+45
NXSHO47Dk/ti8M5uXbwTopPdYFPiz7I2AHnAYb0zwnxnEZmGTMI4gXpwhEifQa/FeT8qwxOc/GKG
Cvi+4o4nvK2K3cQS7E8nV5A8zNw6l4OGZUyfjsfdeoLcU0oKmIcZZqajxa7plCMnujawMZGlUWpq
itr2ZAeL2a+1S14l77h0xfFNqauNVXz8M6+It286Y2ujaV67DHN/wXBWIc76uamy/hrZr/XVY6WU
RCW5sizZaPKtP2UDj3rsr54C0mTeuTUknwWG1CUz8tYXvg/yOvNg8qGaRhqzpbdCjzw8i1xx+oo4
ucqKn6T8zcmywYS1NqM9vLtgHaASnpegtLvBkW4kHcfUibs/5qGUTKI2txkMy+MIgRmqFIq2nRLc
/2S+wBBCPiY5v1Gbyba3ByK8cd/aqED7ewOWgujdwdVa/ezwonH/RFCMiIVGKRyI7hWqd4Q3hXXo
YItU9QZUKdCIDIrUUKE84DLyH3CM0l033d4tPGAoo8CY720CMDSFmTkVhvwldaEPVv3v7dP8I9+9
PzKhygcpkiJ3MjLTavuszimGLvVKJKHWYbb7+Yiz0cL7xg/XIhR6KDMR2aAXlnj941oIDswHi6cJ
p47GulcqNj72g8JtyPg68dfOq1AqCJoOasRR2ladnrRtm6tTVQmXxYiOeSvP5MmeQRZTPNnqxXf5
9FEUaJwLM4MpNMuHUqKYriRydhBJfhiuG1aUd38fjJU3VNH+Br1Z75QhaGt8TP+ZZIeGFKWUT3n9
FQmSHQoggSU5aiUsFn1gF2jRXx9EG4I9Ako/Wm6L5Ex7m1ECdSkere1cPrSpL7n+x+GqjM0aU31+
25nI27FWgxznsZgA4SSB682t/5oiI+DIBmdRfFKRv2F8O6ICwKB4RdqmWaAMezsvh4Vr/7DoLEx6
8qKVoxP1Ey7m9ROAR2Vlu61WMaYDDfy+TBRohSS77WEWXn+G0aI1lMfVJ6XUQuSK0VnksjRNs6fa
1uIJRV9Qb+PD8AABCMOpdvQ7uSDObf9lZow1DKh+YMXHSAW5aSlUkYnzt9eHbUILYmQKcKFRRahf
Fk4FkFj1rkgW8HcgLiwsYlQKA4N8xvFEo9IeEZsGZ9c56SQs85REALtiSH5JA8uH5q+4eg80gAz7
ssY/80Xn7aPe8gmc/sAKwPeIeHTomIKWLcF6tIBLwGHmL9IXsK/aFPmvc6YQsvBEcK7dU7d0py5b
SVOVLYOGTB6b3WIchkZdBlP02EYeLQOihe86I3uWg8N+rAtzT584BI13cQ6hrdJNGcuP6KvtnDjW
1/mYnnlEdbV56HtzvEfQS/I6xGUez32w2GU0I/LLNiPHsMQesC0T2GBWXAEH0u15qYbDQptco5PX
w5CesZLX3wkAaqE5YQtuW5RTFfHVoCEhl/HWv2AtMyzr9XU4puL26HmRT6JS+XH9b039CZESmjQr
Ni5Hsf9GNeTsODoMzzejCgeTGDwzo18E5HHni5ZCO8h7+I9eTr9MRwArG5BBJtAo/o2fWPb6+eAp
z7ww5AZm20zkKGU/KAP3f5lWu8pBWRnuPb6BvP1GUzg5JWv2q38sOk8wEZT81vNnB97iwgncFAuC
EiK12f2p6ulQ5iC9z5dUd3xYRl3JI382oRxxoxf+8HvpwNID16wCB3vaBLwNE3Q30zpdlfnBUGDu
zWqY/vD+DUnvhCmA1I2K6HzlRVx8nFQXSMnlBXiOVfn5H3UC60C7dzqh0q4u0gxqEli8WFfuSqfz
D9SW2Pr5BDgBSCM6iaeof4SL6JRiOTS4vKCGZYEspYZv8V7gzIWO7DjOwJH6QTm7q9LhvKvrn8aw
G+S++wK5lST2sC8UZD/TY54XVLZ6lxNhYUxWdrt+4DSHxcdn2ZaFvXptOk2XubziSYYyA3nf5TMa
oEEaLodDa5X20Qt98smkrDn1sRaFkvItSsTv1RNhYUEryf4xdJ1X1ufTOvZKFm0yu4M8kX5xM6qB
97N7OzaTqhXz379a9B+83FCKmU0Js0SaI57IcdEpTPp2IkXf5pjzlAKTM0a+r5MUlaYXRLtk5WTm
7uUnX92T3qnhNQLu7Txw4+ZT8WtoAexr4BPEogFaiivIT/w1/PHen5Duqrh3pA2fpCS1RlwjvHCv
vs2TT34Wp8megdQhe9jkt1bg1F6rBRIxYYb3ZG7Zs42VAYpNtWoX8jAJdnvTTE3vVH20l/zvTQ2L
4tvNOTRwSrzCgfGKML8HCsfyMxSNnpRPfwm2OkbwsLXVIUhtuCcxdDKLlkxsEx5FIO/dnAFpk5zN
kWCxlHlnUShppQzvW0ASqcBIrMgHRig3FOhQ97dt9IyFDrkj2tWf3U24/4YNwF/uJne2sVrByjQ2
Owu0qt0iYT7lDOZLNT8r28eezoVpxg/E2qSyX86VuI1TiwGfWxMi5waoZku8ReBl0YEjqn+9Tp0c
rk4KynTyZy51bTFZYgvOFa3vzPyq1s3wYHfC+rFaPfVFOd60gbxjpU5Y4FltynStELw21MKcbcBz
oui1e7S1Apcf6p42XLzLlKwwHBcAVot/WTrJse3oA4CU2TT71V0FIjSjDgWDH5rEcFTNBNR6P4vF
0tuBWUMBOGrBogwr8LEW+0quk50p1G1o82fhPuli7ceDhhvnHCxOnGIeMYhC07TrwtZeH5kpVc4n
siGwlaqksAjrBurbvJBK8hG7FOsYuQ6FgTpHBU7Cum4QJqmjxFlvkO1BrZfSa+NPWAT/oMbHsUZN
bQaF0RhQ7y51WbcVnIqQE3vtgmyNMouvi4CLL8np91bo36QMaRzqpbpZBBtt+hOKCN5s6/P/Ewvo
wR8zzKu3/nBKB/D/LzDtexDvhzi1zoXvMcBmpqlt7Nl4rV9EZe7EjKbEOBZNfwBmtFceG/+QcZmT
IFahOIZugwFM0WDiMwY2TBjstznXmULEtTgpBAtGRFHNAMX2NBwx90ivBCDai4XOBlHnkNT5OxTJ
44EOwR3wS6nFJjz2djxS5Jw3LADS1NNBEZace41An4vDhx2pV+HI0CVHCAJEWyo4/YvxIAhFKM1p
cRcesotv81Z1KSMZoazR1GuJqDNTi6eJiHymVba09mHWr88U/ZFgh7xtbCLTk4tiQTOHapIsMRiM
Xd4umUkp/DzHNvytCcfNXGuCqjnlEwE9h2roNva1I/HRTMjPP/knBV0U2VJR9j4y6GHeQTnbSZj3
yhYhCOyYqSW+nLJmLRY26ZMnOyrwJAo0lqhyVdILkm9p2WaGshwlAM3XP8UnVVojDVmYOv/cVeG+
j5lmAzS2hxIvSZbqE0735V+62UvsunUpqysl5vsjd5w4d5JipxqbE/sE3Vhz6NfcMLO49K0FXIbA
l80vL/PYXzuIY5vaSzFBHAdzQmVNR+OYRgrzctiDmX6JlqJ+zuc9c3KNCMLBrHCxUaCdMNsadwS0
vKLc46s4obzxL1e/P7N33PMKqnU6TnFFWBvQiC7q/91RiU1sk0CCidZ9yjrCSuAueD8mo7HjRk8L
euywrfvjbaXs9ukpGHE0mY2N7P6Oup/ifPPO9Cs6mMCnQ6fTeD581XaRSsxe/JDCiWdeU9jAuE6k
Eb+CPr5BVVhcDogwuUVlpRSMOga8mvJwgtQhFm6xX2COmuTwhC3UZaeOUH9GMo8psrgYXvAL15uE
DN9wlU0eTGJwgRgpA5hdZo6LFXDPbLTKRLcZX+bFV4/o+W3XloFm9Szg6RIxcCv3YFf+48fz7cYs
XEQwrHdQHsj/KKfvMZJLx/26hFlfOinHZmAcN8m2/HyQqvzNTldmJmCgmQd3EK+nqY0TeOKwbMLE
l6PM5xkHD+TZMowUHg/TAgrCeqyDhDiDUXMQBC06J70lB7nYkObb7luAztfKs3SYV/qg5Qo3YNWo
Uej+JRBFV5DNy3PLyotclt3lXFYQJKLTGD8fyatF5pG6NRFtzN5lD0AE/PGfKLxQj/0L01ahYeLJ
B037NY2I1f4MYByrTG6O6hCwfU79YePw3Nl2ydSAl5liQmswko58m3NrRx0kCathXzezw3giXsAg
Z2oJIwkbi7b2kAkMXk97+qV6Xg0oTgaU5ucWufbFr3+LmFnWNZYGwZwyHVGfoWG3QLwIMFNrTkZ6
yRCIs7Nb07fJEzbwj2WMKuaDLApYEMH1w6I2kbqgieGIoJ2zw/Ghvin9D924zsdbYk/513yDjPd8
OPPM3Hx5PCGPbyYT5t9wTnLzyEm6ZmOl86rOjOa4/ETrSr47NmFQAHahRMo+JS3N7kgwGhvzNHdj
fl/3YdMy+pIilYUlDF1EG6xc8fEUB9TWe5fhzpQE3ZQxVV6L/vy2xJG9slGyqcSs+G61LSEB7DkL
0kjrdeQBeetzqE5Y1wdynlqqtroG79J3yDDDsmw6195dyeMtHthd5pvJj9Jqv6S+rRP/a6/tp96/
yj+4WO8cJece0gYjGa0I39kTrcXab3K+LZhNIEqWHpbXloNQUpcrPbe00TTDniiVXmdAV97Io7kz
0d5SIBXKAslot+K1ebAMKLubEcGNUTrfQiexdMQ/igmDNCRrM00Y6sGsCZ6jSUcZ+S/8KQzxzFpI
LuQatM+NyzEQ9JO961Gb7iQ5rEpmcPOTk5M/svYf4MLBJUtg+RCi29cLUcSldmN2mqlRIEuRJciH
iR37/WEdEkx8KHTPeqhVZ+EAlNFKMG7Rn2jCO4O4RVLXU3TYJMRlR/gTRAhJgz4CRC/u6Y403th/
v+l5TZwN4j+R11wyDTnFGbZiuYSp95MwiJK2AjIEHorW5x3didEJ6spu5fXWnbiTJU4Rqv1SFYHj
gchuNU4rD8ATgKjcGhRc3/+u+CMXL+0pCBJvOH2YjqIOaYYkePxREnzHlYJ1bfil0GrQpPLhjS0u
SOIeP5y61A9C9Y2ute9XNcZgZqG6JEZz97GCANiWiCORmxp9cdIwfeOjgm7wl7laUxZv7gv7gehK
I2jjZ8w3qH5NlL2g+JZnLK1mbTxnxakQfVuiWVghRjMEHfcBqNN+xgu9SGO3MZLtBjVDubMVpJgV
yrYefxqxVvRptOSztcuZA2ZDb9YSzyzvcWNoq9cy30SuABhjZWiYyVrOPYRR0z1En2cOk62JmCUD
nbEKUibiFBUQAFofujQ27eTZWpOJH6qSy+4GWAxOE3DQiXbHHzXGCcjWJBlbt6/s88mgS1Rkcrlb
NaLt0NNtdHvk2x524bMxVpGGEsENz74+ejltWfVK6YqJNx3TiLeP0UAVsFesLYsqS44AkdoQFxoY
ahnCORMDcVmdzu55DtMX8fBSrRnbKp3lL6BH1fh5gBeGFfttCVbbDbW19NLzLZOU9D6YQryraa7S
30ZkoGvBTbDoJqdLFJ/yIsQg2kkgaQIV9Pl47AoAB++kcFX6ox+wS8QloY9HObZ4YglfKuUwOC7N
7vywk2ltHmsLaHbV9neE9uzwrNzU+Rorc/ofLE71PyeOcdaeLWkdA8JD6H4m+HmnbNhqC420bizB
l+Muib6k7QceysSMHnwF1KHZmVF8u29N3HIc4IayS2AAQ8j8L1IZ9cbpdk2AvdKirwR+mSl8yJ2W
YtzrTgYg0hNoNXtW+wMOHiznCzLaK0OtOLRp8NaZWPF/mimSg/KpWUNdMAqvL6tXhLj8vR++xlDj
5tdFoajDvS0kM0cRVhqiFhaAK2+7RtVT5LdZgVlDbHCRM5er5mx6T88It/kU18kCVP6Fp9SinmhO
B6TgAoaQslWg6I0/ve6lOhfMHh8Ofn6q9jtbUC5ghf3xkgZ6wG1lWauoH3zXmuGKQ1yblR2H81Vd
uYWLeRgHtPtwWNu80zrLT9eMpylx7sQyxX95+N+kGVwH3CjOPQNF2TbEZ6Sqd8winE5YA4RCJFDJ
AocyW3zNQu+azrZfdOwE5fRX91BKDPTdZ3I1y/OCPDMUSxvnK8h5L7YT4PpU2ghSR7nNOTzrHHQq
XQSSfiM6ZRcZHyHyMfuG2NZ6XLjltrr4nntZrzsAgL4uG8vv9kUgX/x29nxEiflOMn6x9WpgydqT
Mj2G9lkntItmNhn9q4nP7kldGLo1aYO0XCHmV0I3Z9JX9UbibjUXceDbkCbAmDrHy15rEIKjY1NX
R6APZ9IBf6OmZ6a6LWABwLNX7xbQfnp4bH3CuOED3c+61VcWIGvEiYbgQs9S6l55nwJN8jCi7iPh
y3PxVsVISJZyNdkvYUqURMBVSJDV6JoyqjCjcdC5XnYai4wnoh6k57qY5m4DPqR7azRnlZUglzGG
CfBWa7t+uDpRTW2HFxuPPXBw4gXD+nsSv/tGmPcEa6HG/wSFcbUKVf5gGArkyquI5cZw6FAOdnO+
06khd43HjO6O7AO1c+y2IfN28CA2znn9mhQ7NLP20Hi3DjjGXk9WhF7Yx8t/HaGAU/zzJhTl1BsX
/joDKL9dQlR9BzYn90etRhk3oTk1DzvT/pJLt1peBJ15JB9cdAWen7ZA5gTS8JGVLwjlJq4ygqZA
eRZH1ip5xxjUYRoCPJtsjS2OlHmQGmSZ6E23lE6yh+NK98vJg0zErSc33F6lGxxTL+Q1SdIkCcUA
Vt6jKqCitvt66UlkNC+vtycLF0Zm2zR23FCXDsmFOV0Lri9zEIiQ1TIWAolg2Ark03QSeNgkkQpF
V/TOtVy8xHL1QfvD8ayA+fZhCWABQtYr7I2OQhaOgY72rTRhJP86RwnYCbzo7rARTcMJk6d2wCPN
AwIsIdpZjD0qyvHElCRDmBZZsgs5S/nGJK39ia8Ujocdu0uRiNx/r7Xk/JQTcZYCgoR3MX6PzoD3
RmCYIYxphdmPVweilpUs2MCiJC5kibxG2TtJgaZ7bD0jgYOyJY4HpftnHyhJ6mGgPnioBRAgNcft
fIz0+aV8DmrIbhA9H94l/FkhNO9kzBBTauBqEUR7wQrdZlM8pEC6wVeegn2J6Xpbyc4qWlh0G3la
FXaADdGV2c4MyC6MX3eeaST2O5FIf88sBmskC3zxm+gvsdAfWg97f08FcKvsO9pRmfuFge9lO5q4
Yfk0MigVDUNS+NOyZsX+rMe9ZNfbsBWkmBXX9/te/AiFVzacYnmQe0o0reXSFaFpfJeGVgmSTPGp
pnCIZ8Yus1BQLBel5ZDM/RKfqpe4v1QRBHHwBSjbq/ePRinjDWftS6BXdXEC9b++Kd3kedtyzOeQ
dL9pNZNzqmAVkqC+TBBm54HEWfYGuXQAGzRB8X2BFmru0ILjW1DRj2sFvhwVxgz9u4R9UVcrKRym
iuMChfhImzFptbK+MM+b5e73QTqk7MiB8GIipzCkyiRFaEiQ0B7XMKX0/vt6+qNjbeaJ2fKCjt1a
0fR/A0WnV2zF12yqAOtXaoOAMlpfndNhNOUB4UG8fmhb1TR1tS1hkZyP6MhzZMxSg83dEdHlrFK0
9dfezz7vnwfk6K0sND5/E15zqfZdL/E9kUzA0X8CvplmWWVLu7d7/awDBVgHgeGTBJ+N7kDLuaPH
EqAoy4/HRx4YHtvlgKy9ftAqcQr0MRLoKj4JKEMZqpLgDb8HeV87rCL5um4BZuf9e8kDYJ6Xgxns
g6w+/pW5/kM+8bVUOf20KSuULH5viXXxnUCChqgLpTUdKjah8XzSgcIURtIqy9lRZzVliXYE29KV
kXEB3yKzWOms+tZUystfLo9TP2iVDd9vZdsfPfPA68O5/8bPNb/wVzjZFGkC3LHjtpr8YzPEWJE2
NBkoI9yjVF8PRyrlaUaxoyLTIv4aHbs8wUHkD9haLC5l74zZlyBHAVG9vOAIpq0gc2v3jLGpKZB3
bZ6HPRBcU5CKa6loqPQauVMnxZ7lMJNavlsmW5il1PDW563aG2GGCWV79NO9Tzd/oeaDxERSfdG7
+CVDsbGQo7gU783hfMDW9bzU0/fc96PIgTRDUi3guWalHJGpW3TUngPhHs2NeZoxNVJpB3w69u8m
zSFBx5mcEwsRatLk2fgltdPmgW1vLum9v6Fven71FdzMuCajahBt3oEyHQAETtZA1Yb+U41gT+bl
KuB3y1YCcODbOVjpFHbhrkYq11o7BDwNcKZhrv4Kt5KMHCo0YPoGXOgoo9WGW7TGaPfJHhbxb0Zj
IXHo9qsUzTS2FJhu/dvTE9jEXUn5ltYNtUy2D8X7+a6JEdSGIOMm6pwn175O9diKfABfDJVymW6c
WYRxyqwXx125FUN/806cI93UeyOUI4gvHH1c/+4ujjM9LdYeDqEGqR8D/KnsB87zU+gF06InnvB8
qYqeoWOyUOGnYwFI+iSHanin0B58Cy8OTm32ySQdeML5mrpxP0iFQC6SJlGaw6ifkbVD8Mggy2ez
ssyq3p9DG1fYrxfZzH+nQ6RgLRmATlJfKk1kpv278sxYnAP7evxV7997mnS8h1mzvd+J5wNRqkE/
yvuwdWnXsKTOrPZKzSBYf/pKxmk/mhs3slfVCtG3MWU5Bb6DOQoBk/sgzhH5ArrNWp8jl/W3f0T4
vcqO3Zi6LgyWkdxca1r7AjB/7/GnjQa1+XGDnQnGcdArp8WHdShAN7NKiEE8OOXU+USGUA90G4E1
KIFz11l9nn8i+R9AbktC1bPj1gia+Jx4Abmw/bDCeyni5xp4laXNwymChgHlI3VAoNQYqNDAHC9P
79AbRdsQZ1SGO853LW7Q/LmYop/RStoispL2+pCuI7WFuWiXKOLeNCcSyFuu3t0+CoEJk4zX99Qa
obAF9N7sJwFrLFWvYG8mOiTqSXypq8hH+mr0GgbdkzHnmnPRADSsiqFKJXuVCB6Wbcz63wVr0gQn
CO2u7B8UGPDFCDs0Orw4IE36cgcGdpu5roFq3jSm5VLPD4T0K7ysEj1qV+b1rR61L9X6P0hVNVEc
7W8XbmIGNNJFjUocDCk5/wwFvzsCwuXAN3BsvJ8RyRB1jPyusV4bkDdlWOfpiJ6FruTwMxgskN7z
jFIs7rwVaAlQfz+c9MBwKfFG2zGG8DNs10yG/HN9fcTzpji3mJUE30ApVUFi4U8dqvLuixsJOqeK
LmB/5ZD+rdciD7+uzrieC+Hsk7cQk/FQ6FNQsUe7R8RAn//Rx1cbWpEsREy7DwT8OSBiinvHY41R
LtURNXwKKOIZyeoKWjPh/N22WM3LZrBgnv7Y3RbCgymY4U7ZxRVJeBLBHi3itaTIXIxPPm6ReyM+
B8RvfYt5hjhnb0H1ENDZPO5ER0yHta3CTxaSKRMFvZVec2JwwxALusWAGAVLiqLGsyBr6SLZQ9ED
uTbnOidP1C7XzfbDYBHwz/5VxTDX/GZpoM1YiTwsh7qiCoXf8hLzCf4SjXVrPZtWktzJpo1YRJ10
khB/RMPN9FLFwLwJmHYNxd38KJFPczDSVt+2hSUL2BVc6vHWDirec5QvzSZjO6dtKYWVOgpLECiF
KlgCFmZo8ndkiNpQjpXZi1prX8IpmWYI2xhS3ry1FxN17vsr/DT1h0iSIbMmgpVelleFxGTF6ILh
OiuoAF+vUPCRtOcrj2xXAFvnWS4+MSJWo4eKfWdO6Y4aKRQy4gpPiMV+rDBxAxUZgdLHpMzT9F5M
v3YFAP7qjrrdaNK2ezof4HTCcN94OVa6d3jTYeD6udHEbWzKN0AQTR5zgN5PvCcZePgTVsNy0sDB
3Xe5fKvTmod+wkV+4SzejKb1VDQV84W1KXzql7AYasnGU+bDo69NfZvKG4y78p81X+p/WOvB/uTJ
qxZcO8DCXLo942Y/NJkhSXNlyTbMY0qzCVVN/kU5lFtGK3zg4TPr7iTenY+2ufRJ3uLvdMSrSume
T95E8MQtkXD0VO685aTcblhbeEm8CaAaEahqGujLcZm4JDY+hYft8gn6CUGI/tGJlt7yMoP5tpQt
AyI/zcTMvPNaAFpVYmlgs6THs+9blqyCUEUGzD5dC7ZZYc85J3vSlXsSVBi9h7xWvzq5QiKygUQm
FsI0qO/IhoFYy+E+VTsjdwQGFRUgyS69FUUOe07ZS/qvTtPRB7G4LhSyc/GPmTmdIQe4yTqYTu73
nVTE5Ogq3dFuRWqZi0ERkngndSubCh4kNMWPJVfBjH9KS+tcgW0vwDFswcz+VOt4YrorGE4WOtvi
q2+9H9xMa5jQY7QbT9+W16v5EqYrlkivIPfpgpHqDAgMxFx049frBNVIrEc8sPJysO1tk8UoC15v
9ACTcoM1PBA6BO4u2SIGTBBRq87ryHAegxmpLL4pdIhG7JjpcFzTbRKcnyoERaq4er4JzdXFJqUe
EtiCASmBkeJdP70uDOtDtm087DvY4yEMXpvCjvT+AZqAW8gxvOE4ZbJA2NY3qVK8y/WxYvdrr+/6
PVSC263hSUPA2EfY5UHgVjGrXXtav09qwoCRoE8RamfwUyW5TpPGibjJb0z7gfL/xuXwcLme0WAF
Gba8i9FRCy8qvZAK1f6LR6JRy2OXGZcQRhlamBTc+Jwbt7Ld/LaG05/CamQq1Vr0fdkFDIBbCnjk
+GZp3OKNIBP4tcPYkPQSCgoYez4hNOHIJhDArDsQS0Mj9L5TGz/tBIB3KnFmArFD04bhr79q2i9t
XwR7rPh/Z0UWZ4FKC65rC2ky/lFHFRdDYvYz3wn1fTpX+WvmG44ljOtwrSWH4ANm3Z6w/bQbDRjx
nQ/hwTj7VdDalm3F01EY1ekGem+a3MP+g9s/xPt4GToqo65ONZQ3XnCew+pTtssNpqj9CGvOMLEz
h4J5m0viFCRemltbtGbMAacO0HjG4LEP77fPB6K0WZO0QbjcH/v/K7cK0bhr1YpLjvMD75yGGb2d
DHQQ9KhjJeXlAKuk/NAODOhQYzU/ArZsVxdq6dtZbbjU+Yfs8s1cPPNThv22j5yRliobM8F7Tdds
uk4wDW+MWv+nFA9752NxQUmDeqxjUfuTRj0nd71F8p+aLs4qQYZzrquMokSR9Lrthw0tEQWmOAiU
8NF83agB3izfL/Yj00F46rrjX/NxFoTmx65nGoRDg0W9GmXafke3g4p9I9utGOHBzYV+PBPfFdDb
IahDxffW4bC4JlMMCd9kQe/QuFEEzjBp82AwDm5Fvq3BXFXdDY5jOI0NCOCgpBNEgewVfHrvFhH/
MQ27rZuYk8U3SimLAN9v2U0dGDXIHpPkPTt8TDHFhqUTPJPD75o+gzBGnIYdNR1pBCB+DVL4GhC9
m3b8I83MTm/9CXtI6fFY0cUHKzRMveTmLYE5aayFpK6OvWXcmf0K/AwqSq5Tk5lBm+mOvJiYcZds
RKr1KCGJLEirEZLwl/nG7qE7vschPawSGBvZGQG9kU2+g0ZceDCbGr2peej9LzBOFFa0x6umLC96
48ZUcbXJI0vXwBlj6Nwk+shkOf6uEKAMuV1zMmSEtJp6hF/ULlK0GkxRFLmnI+M/pqu9HOIjWXSN
ZO+Py7AhUYMsrF5Zv2lWtlMOQ13Trxs0WGgWEA6GzUgdx1XauBT4CZdqtRNagBHyme7YgfaQSx1b
vxturWU03cUo+ZlhVgyh03iNngPenDzr66CbmYgXN/Ema6Zv+FmaFc8JAdDx6m2Ce2DkSwvbC4gK
BEP0aEcwpatmoUGUdIF9dCvhLO865KsY43mbxbAJdJxI+8MoRSD2BJIHDK2guheoWssURihiVTry
mDGPVU3+foTMgRyWq/7H92DaTI1P14rC37L3UwXaEoMNufeuBwnxjnVyfrikPxtP8M7QUCtuyGZe
P6yA2DbD/8SuSqRSUSCIOTftAr/n4Wec3F781EmctHjnNOkwccRZ80Nz2eCktv+xDC7QWQvOeKsU
c83le6hWxiIhAQA5jJ5yxLOOJxGQmOg4iGmh3LVWxSsQ5SI2t7aWD8oFZzuUh9snBaOow7g82qvG
c0TGkRYNT+GXGRNRGA0hBpUmDr/sSUKFENYmO6f+3VYl76PsQi5yttQBDVr535d60RS73HaU+POK
RsHZtjHfHSVoA65V8fc6hVbWfcY1MLr9eCcl/bDMXnaHnSGVh5b18o5uBDvQaMTfX1VV5Jpzhkae
1GNhy/GoIZ0F95bHTNW6tCh1j8XraQg3H3JRuGuRz04LrmrCOttawgoyLCxEcrfmqsfOMgiKNl6b
heUp/kCLhx2ienT/n53lY2i3HT5aYgfdHEZQIktwRHF2y9HDQqMCsQh55ZRFapW83cPoq8EhUpL7
ZefMHqaSu9fbCex1hzqTjqnvea4fAH/QjAzzTPSJoOUzQOt+SkI/+K4zOYpvq8Com8lnFfQ6907y
UkUWzNHQFoXZjXcpD9rcMliyMsmLhVGfmBWTlo6QH2O7Odsej0qaF3QrHNgsxU1J2BZIxz5GRPry
GROcqK9p9IW7JKRs3XuA+Od68V3T+jY5wniSLLc6WBJ/X14poj5OQR/dMgA0MeOhJI25u+IM8jFU
EARFviw/VIv3TpFYBBeSX6jCjhOTRZS4UofnBU84gctHJlqzAfVFOq4OVmRTV07WsXiVjlJ9KbEM
Jv7Y+IWkpyzOsvqQtarN7ESQI10BJcT0rc6E+Ed3SuoYN5rGcB6bZVDIBxBU4hpGelEONjqJqF73
sCSZJousVnbF46VUh+QlR0SuszPR8SG8JEjmHeY9EghUegVUg+haU72ISpgJ2AJvpUmgFYX2SrOD
n40W4f2PI+YGIplz6fasMFlsx2mbdAXb0LmhMI+zZlDWnSEoNvCokGPsWO4vPS/MRcrsK22Nh+CV
op74sNj9nr34ZDrPEsygrMwZ7SRdcnVxMamIrpBZmGg30NI3hy1dXAiSEWs0zykXKlTT0Ddt0K+g
LRgM3F+uYuLB0b7wcFa1IcbxlgAvuYO2ZLan98E2SAsgT0t6gmfN6d+g4i3Iniu7+nM20LvISMWo
2YbRlpprnexG9dunaDy+iD5nfkUQllEGNlFwJNjxCQZKZiXcidbuu1eBOcXCtiUhzzb5aTObfAsp
r80DTKvg4g3C/9XaDo92izcoO6VqnDjgCvrzE5w95sDtX2VU3o9XiF2pFm3dCY3dBeLCUd9Y6dJ0
OywdBo0yFeDLPRAJQqQyc+wqtPE//zvMHk3CXuZoGmPSDxptSCDQYcxf84KoaAo9A0FWuQxqdIiN
lbAoXBwLSJ0+GGCOnew8qZOHouFhrVKhlYlK4Ns/x1GlvqL1VIAquDOy/UOdNT7cQCoTiAu0BSUy
MsamGZrkGVdX/Sdabr1T64Tg+pgH0OgYV0NwuH00mGFEcLlG6eslceD82Il6zW8Bq7eL6uog4nxK
3epNUoCmj73HdgFMjNWMIzVWqiqkFcvV7wjxCyM/uM4UtgKK3ng9u//y2KeGKWn8Shgnn5HorwxY
gekCo7XiLMNImhfLsp6Gbo6qui3hvzHwpaTU0McQ7eUBod3hDxOL1bhOJUfYC140BoPJO541/a1/
XzUF/BGq6etnQ8yEfkWVYxE0jNtzTEeu1+yDZQQAo11UQJaWRs3/KvZD7FWlzGnUDAztlDn/E9xg
AZ3pZdHdW0GkMt0SUjSV1OZWOp/P6qnafxS6LDm/Q9dfnUAA+SN3ywatVZXwls2vCH5/jvYxPyqo
htboXkX3n5ggQQ+0FZb5lPUvlr0M67L1y6y05PBeZTHdwrLSyESJbk5mFh90IX0rQfwJ2+IhqvhE
P8nLlfloAX4brr7lzs7c6VCeM7nkiiAz7TnjX9dz3tLwXmMdTWq4wnfVOowCc5zZeoho5XROugVU
Oi3mrRJ1z3EfJ8Ru4wEZQb4SWU1JvCvH+hzwbg5snJeekrx32Ad0q3pRktB5c4HwuX6jWNVkP/r0
FUeBsPOTG0+3kyl7FWZdsAzWRis5E1kRUNpNYMlYY24QuSKDKJaiOECPyZYkyrVmZrGVGDAhjbjd
dG57uBfUY31dnqd/lEgtZs7qt83xpbH8rVP266g4wifHEk8PeCZ3znreV9cEwZPm1CTyyQN8kNGv
nDcDD5lZruzUGU5+vIfg5qyCm7t0nWhsdImGb5N2sOoEI4Z5JQE/tNgoqXeE0+y4E54lOaHsvRgj
Z4oAXD22i96HOeJgy19jCEG2tppUOBAwYtBgtjJnCkc620kZre2TcjqHmzfuy2G+PDwU5dH9iXCR
+vCLNbUAP8w5AGy9m1OSLXo4tJye+wjMrUjU+uN+jk0PSNI2MDwd056FCkX51zSYYiiKIwrlch+w
x3OpW9Y2k459xVzXljDnP9WBqXUSPc3YqobZr00lNTYKWntLt8O6Jzk41y6CLGjkJ8dRiDjsBRwr
qTqN3+BdG7W2pcUPRjZDP4h6Lh7Oe9UDCV5GdD77AosTIDVcsH2jOUenYcDANNuQ7wA6Y3fkXS23
crn9ohQossdBO10VgHD44NATlVRKkNJ//rbFwAT1E7v9SeVKrEZQ11MdNHuT4aU6b9T9UJ/ULyBe
TT4TTs3YWmZMyldhf3t+uhGUzu3TCauEGxDx2gzXy92t+s/LvxKn37VHEVlrzU0rJGGJV4h+7UbX
iZ6Xo3D858WWkE7qfNr12kl7z55TNaFWG747LHkOApvk/FFTlkmKRT0OS811WiBDwLkjXPSE/LiS
j7gZ+rtVHVnHkcWXKNinJav37vvoXQcRLHU/bGiDtrGiMP5QQDll1H93W0qlC9GWS2p0IIwLQBuk
+vxqzCICjWiW0vFgt904DA+wc9exhznLDPQrVe6wyZ0U+bDdQnCKpPFJ/bXVcOC3qJV4BjjfSv/Z
llykxb7RZ+Ll16GGRgI0nBz1EUhnc/g3W7jYpjcEknlY8179zvQ0N1ACWomLlPBtOlIrgouEx2wF
W85iONsvxXem3VTNsPjMvxk7B6lR/IZmXa2MSrbGd6rKzjO601EwDSlx2L7kXlq+g+gHdLcgRIif
flCRomDqWXLrvGkejwAMW90yjeeImhWYV1tytZkYgNUOJ45i/QcxdbvqwhezBJz6ught8bkuIddr
8exXBPEly2ndEN+8SBUlbaOodeqxr0daDX2paKMywZGu9RdlCh9d0ck/zlUZsItBiNgyteRue5Oy
0EMh3JhSaVLpVmqltYgeYyKWqk0Z5MdhmUFIzv0jVYScVwWG5s8weYLdlq0KMhZEIhGdG20blxsR
4GLF57XVCLCSwDGYpYawwB+o4Cu8cSWEbP4rUD6K2Pb2ocg+pSVPdx1gsmsF5Us2SfKiklf65Coo
O7sOzCr1ghmtRFILe8gDHUp5adP1nQP19126ZFI3AlNZvUuF9obZ11He5oWs1wuJibWH5sAXRD73
dy6W4/OGQb6KCCstA97suwN0x2pn/Y+NrRsTEMmYso7TIzS6vW0ItWeooTj5OuUT/2LaMHQRp68G
JAbK9ZYnQMgbqK8OhH8casrhQ/1gKowc1PMwmqY0bGVgHdOUlcoNZZ8BWtgHma+8lYqIt7MtmQtA
RBNl0xVttyysH4eIZIAt577MsExZtNg09jbTmnjPNrf3thh4KS+MACVxBO4cAvoVw1q/gwRh2gKc
fPf2OYGCvDZ7DGcfPMZHkbOD+bvDPXmeQ4/MVSc3kgaXEXA68mdc41IXZXwsbQq83BSnJEW0Be3M
mIqMFwo9nAASjG+GEJ+JOkZq3rPTl8ItpDplkqXdU/Gs/sOnZ8Y083xB8roTXI06zxJtggxMJXbU
dm8UwUZ+FHp+Ve3umzBy/JR7dNrr1prB9hINwSIkttz9+ziAvjUwv9+6aM2Y00kippWONS2RPgcU
wjjClzr2LWG3HIhtAizQtZrhjB9hmPtksG4ihi4L2a6lJmmhKRoBxWPFdITNjItrhQfMnCeUH7cu
+vYS/3OxMQWzSzVdk6mXeZnqHseMRDPRdAgZfrbu6LDaHBiYh5TtRFjkuPTTkAxHesQeCr8uQfUt
o20GfDzywKTBj/wBLWKQ8QXwZcj+La4E7ABS9nvxF6vcscBIY4tBywLUd0zXmUs90LnwtAJGIaR6
Q89q56WqX8aGeayS//Iihuh8NpqhftFz7hsze37VoywJ0x31xJJOFghi+uly1Gfm4I3XzIqre9mY
nSpzfKekcCStI4XUyd5zpVoh3Dx00eR0ucVuszTFoQcJmVqmw6RULYrIwO7H4EwrJxHD/yf4cD/1
oFlgcnn2zvgFeEQ2IKrdzBIKUzMLC7yTlinhdmM3ppHjxxDUxj0ya6AIOle3ndxYCD1l1oZ5+KYC
+7P6a5lGYPjGxsLj1aTOuX/qvhwbwXvNVW9qy7kA+79JxlKeC6bCGL/rFc4g087hHTpkSrbdAFRQ
ocaJs9Dv3ar2pioHrIyCJKyi8wOuGrsob8dHVBKpQ3B+Dj3isNwqpSfwLBEOzJxIEl2zPYZgzG2x
/gfgLP0vHqEek3F26JZ/HBGKTcH9puM75/Ps87TLbFF1zh3CfhaT3qGx7AFmRtLapbwkm7lkh8OU
XvZsXILYOO6oA52N5h7uRwp9McO9AdGdCGMI6BaDZL1EzyXJlkBT1o83TuRH4aYpRYoeC6F43ZGn
xd0sXFJSVaHRXjccXkLngi56bFoZDcoMVJ/yPymBfosGgFwLV7/g/txZnjNsikpm8iRaLGxfl7fa
kIbd4m9xb7s6wOb1A1IibpqkIcMxg5FZCs+NaiYwFVSlKODwztYq+fnRVqARLAOXjXW9hgu6Z9bX
u5SKXlPTAnlPaPRrbNR+iZ6IUjRuMOtvoXQPplwvFkWSfpJUlcuxYnBMZ9yka1AVrzaCPk7zkti+
OwXRZ0tPT5uRVnASWOrmeNUjPouxVl+G8yWvABkPbB4uiKmGPQ2gqrZltaXhxXz6gkIsoe5K1UCA
bB9kex9mWFY6VwhmOX629QGf3/iqBBKX4l4pZK1K04b31VwXurHPlF0XpotfezT+QM3k3tJFpvoW
o7glPwSW7IXdmXvFchYnGtoX/mzfaTy703Sn4kJKyzlH3zEO/04bSrB6HLBxEYc4Lm+LgDpnOSOA
jFMzjHI6K4NIiopQUnzFMhBu/YyCM0/NVSkMSXQ0mynBPwG3oNSlORcUq1XHUabouonna8SYWp59
eaabgH9JsaaqklS3SzspZAUSlN8clekISeAtM4evUwdRoGjWvy/1rzNTELnzaxPLbml6N9srxMAu
PFklA0xx5SdI3izeNZvyVqDEy/zhAWUcsSHXzCByRmCY/GmjQbBbpzU7boKwcK35LEgbU4tBbjKa
rmF/FkiU3J9hcx9uZ9WmSj48QuNZ4MVdfx6kFzB+ZwA3J4fn5bHYbl26/6UTjJIzsr4a+gDHSzlq
iJr8jPJpfOgT7B/Ofc4hJx8e5c3TfB0ijM35vV3KEdgMQZmXp1L149gTEoA3afGLHAjmG375K0JA
m+054v3/b6ZrqA41G+jSWFhFxZAkYY6V56bNPD1KItvW+uOvBfqjxTa0lANJMY3YwH70WF9BYXd8
MzwDFbJbBoBXdY0WcJXnSMq6FD/+xdZ7yXbfnd18K/g7qH+o8uxI3bHiwrLZJez55jmu3NYOExIo
b825bESkymY0G7ilvBmfoh4vkEl+R71PYi1ukx89Bx/+8SKbczXj+gfhyFOUPxu78YrbYZQxGA9l
qDNHexfJssgDbvdsmKEVGvnAJVCqKk8TCRLg/+FNNJOCq808HERSb+8wiTi8Kpw5TXXztiVA7MSK
YuA6odpfpJjYz+flzHhTuHtNY3h2oyzBEX9eqf7mWDB8Qcp4n4WnDdTBnTqJLjgh95faHudRJCiC
Q+neRP6fjYYKZt7JPhQjNDWiAjiiCLuFBkHd2VK8d/JCf2ptNOJQbx3gg9hKmuAcir6I7rErWIKU
jKEN8vo+GbBhui8+h85bmGgRJDXFDjQ7LS8cnGPRxFpq41cMX4ucUyHa57+bY9QLweI+jDUJAPGt
nNqOVFyyogv8icC9Bhy8yfP9jP5Ay+EdEzKbYvPzxx8AjKFlfQFhv6Mk8IzvOeBVtndRf786v5kx
yg1JiEQgzOjkogCEAt+nNuWnQZoLv5qDDqZvq/3853BNkLKWcQqf3lxMQX3/1FQx0B/d4zv1Uvtg
mT+5Q0qK1/CN4XqhecACaS3hznoskoZwjHPrmR1K+JuqodzNzLp54pWKITkkZV8B7i73AfJj7m3J
DTo/F43hpi+xFpOvcBe6cdNM/H5EO64c84r7Tn27RTy6sOQtw0QqpjCr+i7DbveWJsXJ/v8PxSwv
ydJoCjZhkpvNCOCeqOuZa15H6aRonJpRF0+Bnm6Ph3jIwnMxqWeQZbU/gNSHQhlYNXLASZ7PTKjf
c/qBjpHdthQTIb3cHGGxkczQZxSV+mT+/2X9ZpH2DXo+7CcoTIAuGJ/XRGbKjjpE0Gh8HHZ9h8XF
YZKA9B9AEUX00p10B89z5sYeNAvriVWNQ2GYLNrdF3x6qejcE6sTkfIEWBDhs0CMvdTcgaZoO9F6
6pXq5aiDcvFVQR76MR/NSuWr7LIKrTiC7tHEqQfNHDFAPE3nUJ3xGMqY0dHOAh1UrXrtfLbNFrCG
gU1jmERyuJ7YO2+4Sbpk4htpRxFBwjJzefK015BdrjjO6/e3ij4kUzgd1woquvv+jTTU6EGIQm+R
9V8Skviz0wfo8BbEpn0liPn0PyQ7WTzTQJBl251kPJCuJHEiUq+coyj85jQMBzIsombqSAPDaogY
vUGnHpXf09wg0KpyRYz2Lwo6hCGr50FsksKI0b6GnI2m/R/QwijbICppMJPS9WEkBnuyFWfH9eGb
DvcSY2aCnNjLwX73r4oyohfKLfwbF3pG+CBWPal2WD8/V9DUFyfeRUf2tcuK7tzu7SDUJqAq63Y/
kxIH9yJSyV2bo5b4VMHhx6QgdYjYteKIhqWyp06rBRvT+wX7dlb6sH52mwC8v+V1YS+niSGippK9
vpXBKISsoc8V6PxvjPC/mIYe3O3nHxH9xiiVXzCxAwivS1C4Ug0pPVzo5SYoEth+G+EMYjSVWgXv
frGC2sZn7wOw5DhmVhk6E/AEUS+CnSmqad8X8Wv0BZbh4axi4lb8GnijUtOJy3wL+zNSOsciK+9N
7w5ngb3PHJgM+MKmCkUtL29P3cn7RQx3x/2f1+/sk85/pMOJCLnZobiXlwO+1T9B6slT6poU6VlP
4zPzwDR6104LeoeC3ABeQcZnT1uw/jaW0xlHu99yY8AXbZ63sgDEVAsMMsooE0IWI9vyplLiNDEq
9NRllQ8VxKmVmK5IsBBK6LYTbI2glwYG4Zo5QkE7O2vw7AZBMUOk9WYPuruEgs3oJcPt8M3464PB
7MyL8gxF/pks3BSqAYth/sPFjmRZHSIUkOOMhAbydTtgZpaxTusjHO0fTZwKlbHzMcawK92Svy1a
vCicie/qbLE7g/cVuGMr5jIN9y0gXYI+PCrNFq5myDxe1prBetvTFcfY/gNms20Lu5+JAbC+3dWy
54rBXHa25mkAFSYV9wKLJEMoBKBLi/yWXiiM/COnKtbtGQXMJdpHt16kirOJslJQoIDibs8x+oQj
pkUKp1F60zWIVG8WI17HffQTiqaeKs1o9jMfI2PrERACnGD6dS8Wlu8dcK4xNrXUh8pBXECw2UET
8Fp5kD7UhDzyCtDvYU3wokriXlorKg/RS3UaNNymskJMQLL3FX5UlPSwkGj2xPqeZ4AWa17GNBPw
GYdJAe3GJ4r6lscWxxrgm0FlVWSRkhbYPKy6scDFzLE9WgOWWQwWeHdT9oxDX9pqGrVbfXwMwsGx
yFMoXH3TB/mRAXtrzKlG8BrcpgZ0VEO2grF+1XQxxp31CumzYY/BCgURVv7GJ+8Qp9k/BD3FUjs5
IOFUh8Jx/visdQTXQOYiH6QAPJn8k88l9/qxFQ9+oEHSEWC2ezgm6ukykNS1in8otwEuoi1J3WO8
BWP3HTG87Co0ICjTQyFJiihDoLtXgSzgxuW+zOhUntKaUwLWtkbyT1RuR0jOgWnwfSI8SYRGoGGP
D8X82T6a1ak2nBJ2OAiEdwJBEU/Qx2MFj+rjhaoJWAsA2NuQmBygdmG3m+zg9Oi2x35UkIgYb5BL
1WLanA2shm5LfU3UhxaYjQhK1NtiRRo5dxP2KY1OVglKIb1oQzCcc3Mg/Pwl8uDIn81T6C0P3tKp
VIjz+/r9x7Tkm1kvAkWGHl2VZYMGeeT0QU55pL16Cs1TDe2QbBcwRL3k791xdppvwpCZ3E0t/lMt
yW06Bp6h8VusO9vyBOOcYh2IabofDWyDHBAElg8DgncBneW9oVN27XcyJsDlurNANpNNSr6JcXkv
LZjrYyrGezGTYYG9fURbHeEN0HnvOBFK9+YDz2Dg4vhsMZTAYGG6wNrTZ9dDsB3w54fYWK6Q6QZS
ep+AjsOnuZozLmRzU3qNvvZdPkAMwlKT1J3I1xUrqeA0cKTlioFZqemGDXm9Jxf5fwEwEdbGCZP9
WJJKqdmoNrgrqDDe7+XHOn8zTRlIL8j2rvoLrrzpmJxlxeoEnHDf9qsK/Ps+3IcBvEIOSoEkOezi
XKE9BFXQNAafGFsBkvypftKpwJvW7KOaMnfTeSf4MC7LTTWLTcqmGTzMxpq1nYipUtAJA6IjT+jp
aAtutxR79fmd9Jjrv3v5fqlec+HcAO2fy+XApnHIQWtVBZa9tNViIuLEgEB0VpqelblcGmoQ5OQR
+zi9DbxlOn10v45wFx4enjYqzaaVvXzBVsYdNDXa7dlWjIzoopvio1lvDx3rbAagls1GyM+g8d3D
3CCQ012KuietTzQ5uhuqzAdPigzHI8f4t73pvSbYa7LgRs4Y0l7qsO89V7m/IH/XxiAU+NDc03Yt
6MPnf+gwC+H4ceCQe0yiuz2ZwR+MQZCekScMms7q0PMwEz7FDAVctSx5iyD37WT70jZhBjLH0l66
Uv7N2pS6aIUnX5kPJxcBr22gsX5dpQmkZiBZPUCwz/C/RnK75WWr19qaNCCZzUds5puuPN6Zm3Me
vt3CvnuRNnwt1o6X81qdgo6a23RVry1148SHL8WpLPWCzSvsHBNlbLcfn76k/Xr69QTiK4Imb4H4
sxEMtKliioE1twxKNUyKna6bpYM0KdMTyAiiruEGIf2uwn4kiMmXG8eB9wi3ZZwvMNTXyjb/GNz6
jXQEhhAx0akWZpYrBH3SQq/qQuz1bD2v2bK8JFZqMauAO/HJidAb4QrlTFL6ZiLtNbGghvVhGeV4
IqD+4Obny2cCqga2WoUs1EviB+USZbWMKVKuwtrOG/K7HTKTqHuqLDF6XntVP7fUKj8W8c24JItL
I3ke7n4QErpnglXd06C290O9qYDnhqusoadJqhr4dnTb6djizdeO/mHmxTaJQyayfqlQJ0px/a/n
3UOz5vUvek/5aD3fCGiqvvDuhpI6LLa78FX56YQV2Rc1mHtE4oOYl7h/ULxC1z4iGwigZuEPF1K5
ilZSD/mcx4+TMtTDwX/+CcZ//wJYh2AuJNKbsrwNLjJUpW41WxAGZXeidVWm0jPhTNzY1vgLxnKg
Apg/Jwl2ijEGAgeqjJ7uO6vkhX88Cm1lzXpTFhd2TFTsCLArjslkYV/ohZSWyb2zzXhTdXe06XJS
GyfmMtPAfikFaJ+tjSZfnu7eh9rHR/hfh2aKa1vke6GHxqS7XYz0cVd3xkPUH4LeebhUYj6UF/wi
h4ErbbCNrXxWVX8i/4T1B2Idif8tCJLthUPcUugoZx4hOjGlBURnYlFw1Db1DWKGnTsBfnhKxWxR
fXEZbQmlDGTyecYwsrLHZsseU6BEiSRJf3Z46GRkcD43U417XN1q/kq3xPFsqvyIT9+qZOefkphM
2TLAxMHHUIJAtm0xQcHvyI1Nd6EePyWE57QTZ0CLjJI/3rRrdP3JHS3Q9dK2jnWWQWBrxXlpHKTp
ISfyybu0NhMp02/wLDLYqT3awjx80hKo9N5HL2dFs3+0mf2Vtnpo8hjytkypTWaVUvkAPunopT/E
UKd6gRvoLi8OTI2o9qYUPhm0pE4GI5WdVjA1JxJiK9pRZ4eYXz2zM8bXh+6PTUc6cbuH8R6h3mec
7NGTaxz2mcSiwrZ9IZNC8+d/O/3sKnLF872x3HNJuPk2P5LPxP2jRXFlMriw71AdSQR23V4ZwbCn
6tS9GzMbjoXojMbEOuAagT0cbN1KoJoSXqPKOmBhjK0Q3q4T882BkfpbTELSapAc2hJ8UhfMWeiz
oGX4GuRne99pGGHCduK871CJ9TPnr9ltzWj19YQuhQ2Uzscbp3hl6WOAy6g/4m/ICO/0y1KwtBt6
XQ16p/jU5dFuP+96iHBV9b26rSir69anOXHt9Eho/L5ievx3mqg4/FmFDi4AI1OIbw0FJ6Y43Msh
+R4asxX7snKK3ajOHW03bHc7N3BOvUCKknigq1u40cUNAGO6vb8BeESWa8ABrpLATK1bz3OBRfSX
vkw53cDziFp3HYNeGiigJS252ttlwjNLrjDJHaYH/T5UfB2AMapjKyBse62flvqwHIgOBCPAqQj3
Oh5RxFZUMroFNx6mlRTlugSQdUkXbHoY9Ymx9HW5GZRK3w8I2wwvywjkF+94calr7R97v8qovf9C
TFSsUEgBWqs/+dN/meTr3kjCuixqaz4LPTEht6bJ1CIgvy4e27USpQz3MQpufon5Y7TEvqNchp+E
FjK2OdIpq41d9MiCEq3vKhv7MVawziH2I6xD946hvOweGDRt4I4gkllk2DXsW9iP5cLEZdetAVww
lq6Sn3qgjVxS2CeYUStswa9olVCc5UNQpBwwgJExx+FhZ4WRgCXyTPa/WCFM5M/YAhoxieFQ8p0Z
M1BxtXGqxaZnjvXshnyOmw+G7XggKhDF931s9ePAoJeAZ8RZItbBX7q+9FRLi84NM180HWdEPYvr
N/IRE0d9LEgEFCozKkysL1AfZtUzhSkJMHbcxbd1XmQBqE2GHer24jZL4TrzDAmCrkPSplf3VtCE
hArfrE/fVYtZ45CCbKt3+LHB6wZz+VPeFQ9564QqC9MOZiNjnjwi4chI3DcyYewQfqP9W3T7pW7R
doBOjLtZ10GMDVLLV4u5GMuQIiazKzRPllQKNaBK/WwDpCJp1yds9rMV+/pRPTGB2jteWWD8hipj
Z2+SxA7MXknCi+vTPpPErC5amrEkaRjU5t/0xaiLJZQ0o2FFs9w95cevEhjEqikbvlOQqFxxEkBY
HeRYxk/0VFpeEaU5t+LTkrfltYiFR4AbThnCJqLtHrThL6il4o0ZTOmYJHIHsxZ8wN+QWL4RIoFo
h0Fp2SCPoeDLgPyGNiiGCnHfVShUQtoRi9R+m98ARbikH4ruQtbSebfFfmtoHFyYZPMfP9TeLWiK
niopfeihQRG167Uws/PK//NN7nAn0HEGp5835B/9fcyWhk/kVOp1P0pu98ZtODjumgDiDNbqLi45
igmVykqUkqPFC4puNRgSvvkqtoASkSU6/JCDahpMoLTEI0zuscNkO6i3GZci6f4U0CEOok04orM1
Y2C0vpIrE+DU9bDqKNGPGB31C5vOUGbhACv38+mqFpIirfB9uRTW51gwQD20rNNNmLj39dgVIPFN
zx8wuFRRr0R2jqhpce4YyzRPHOuoG/wWPKEc+oAZH0KmBEoTvEdEdQBwD64rFluETdAq4MzdyAGU
ARP6RD97R8To+DYCQHouktWzbu7O18S+Qx67Y9tWZMEXCcBVeW9Zsc2UFFQm4wa6B3EKZ03GH3LJ
iUcHjQIWUbcYau7W21tAqWDIgBT6Sal+RHthxW37tTYfKKmaFWcljT76AfNUpvSsx4CRhP53Ph1+
1KJvYB4Dr6y6K4r4nC+20J+G+dwgmBeYsGyrg3pN7masjVQl5KgD8agXD0tSjGthCztZM481p1iH
k7/nvAdClNWx6ScpZzhhptGGqBxL9c8JROVmKzrupf/5Kg5OOzBsTCr9Gd0X809sRNdT3He/LtVH
NHcCW2pkj0TjcScCsen2lTv1ne5/4Iko7QJ8dzqZsjXcIIGm2mtn7vVSQ9180ub9gwj7fKRbRq2+
esYW5t6kygz3USpB2es2LeE34fS813+6qaGwLJ9LdCK/cB9nHi5Myemxo4pVGe8/ovqC3B/P1ErY
cdDvuZ3FNboxvSb2I/pW2dw1LFeemp4Us+/m8yQ9K5v9Pl8YPSDnwkjq4sFnXjGL2NQGJASpwkZd
x3EbW5h8ARbrKMAaYrkgcf5tY0pNX8xbf5yZwUdzULWaGZV40AWb4KJJOAvxV6SBIkb2TgmkCbAy
f3dFAxPUW1vJpt5i9BbnpP00ZaQ9D77PBbmHiaP5/vOyPFW+FNK25nZG4Et3gOVyTUGflfTrh8kB
An8mTeSjqRE7v7rUeq+5mDvguh0dfsWrt0A7ed+L+51IJlp71aT8+iYP9rMhcdnjcCbplRPj8Cxc
1fJDum2CU4kvzZEAV/pIOJ1VrlclYRjWlU/MH2jrV1ycXKDBTx8VaJWINFnNfALSIRJGb2sME07E
JHxCHmVIrh1tpfGaYbkOTKMHTWQyTDICuKv6u+nMN2LSw2xn1WYvGpg+JgpPARB5gB8Pyzz4/+9G
F85KblNQ4iGbx8Z2D8OJ0hycB9is1IvafS3R/qGq2fqOY176AWxaog6B0HoOu+lr8j/mVTv6nMYn
W5zPWevusbCRRyjHgfyfhngsL540Usy5mN4Qx7lVbLoF93Y6xeQNrRIn2czCodCHINz1T5Fug91+
TuXp3Unf/gXNDxVijlN9xpvESyLcg+nqs2BOCHbcAV3q24BnEPbrDxt7nJmB2ZUg8ILZkLwRCAVu
WewxV4iM32+t7vpe/5w5LU6BjGxrbHbUjI5SgcqTq+yOX4O0QMUIWkfyZAywjrjpsli+G2T+H4QO
PHliaazr9cr4QeKxjiPJ+CFpro8rm5DFWPDOD3ap2dSVO51OOl8nmDLblfEOVVGq/711BFCAsubv
e3MNCW3lxLlZ46pH0Ei2xVEVIaQbbhdSED8wxKxJGH+33y4v4LsINwr8pIFIOPC7CEJO/APwwjSz
FDYVzXh5dgCHfKfEOurMVPW5XkqcGoLtMcQf/oNZ6qR5uGCSBh3PYmNP7/Xz/PTZLxxIAMRwWSnB
K8TaHHbRZJ1WsAGbxbNYcVAzaxfBQxCQNK5besKoutRBtQeNPiEwORWZuw/W/pb076voG8VHGAQl
DLTUOnrUO5neYJbsdV4EKtpPiRCApHZ3fxMYG9hIzP1fZ86nl89+Maw5+Jjc7jQvpJSXLvzHrcZO
vVTLqHKuOgRfPn6wQO6HQoCe9PIaoSPthJTXcbPxqRukzmqEIE9SMYbisSfD3nLDphtxdCqmvYlx
dkwrObNoncrrjzeyucw3mlBui+PYQ22BYBRScVjc2xBGapW3CPO+AsuB1WU/sHBjwQpYT82YhFg0
Dnl4dA7g3zubc8K/efTJ/L39EJ4lTTtNNSYRN/Dbe3/bJEIYg7JZ9mRTaz4u2DVd4VW8dIaEzpuX
2NlmQQSYqb0rCDW0ErUrJU7JPqboBCyKxWo1uoFSn6HWcAYipp7VCxCmHQMUM/AOrq/GqP/pnEmH
nkMgHyxqg1eIDTHpGUc/Ce4/u+j6NdQS7bPh6BZYC+ySMWFRfor4T2/mP/kNSWjiFPXXZfw0Umst
AnVl83LuanlLUJq/XqPeXKygeFpL7h0n92PL+xadt94ejGXOl8rhW/3FH8v4UADR/Nwq9IqL+hXh
PttjQMMz2wurtUAhtAUUTfaY+DjM4mYntenNee/tmZAPEQQTd+a8u0zKR7st9LBxHWzoHtSk21ZT
PDvtcxAQhuShYe3rC6+sFRTwprnkcdz6RFRtuGTnPmfxJoxSLz9c/+qNolx75kUb96DBNqw0dtCu
wxCmBgfooalfNN1xW6rg1DFBf7rcolrbksah9kIgIt8gM39xsRRyK7yfEhXBbtNXQSvSmV7vAAcg
E9+1UBLcgzUMqURa3bfxhrDnAxarsa1ISJ5msLQLEFb9Hir+PwRyjZKxzmj+8tKXZWWRA3+5rEX3
9G7ycjBu1xed19mDi8+WAB3uxkPb0tbbFFWfxp88jDpNHYO6byK/WFYaWL3DSpRDeI/EO5vgSJkT
7Gb0G9ltqJMhhrT6BuV8qGU6owUwtPV510qYIU/BMsgBM55yrOOyfSEdfFSEi/MJtDcZq88RQFtX
TZazbjuqGsmPUWK/QekbaLPeDYk/DbW7HOALRLbNLrqAdyQAYdVzU8nmr+DyicIDQAQWI5vafYrj
CHZoMLfeBBwy7xFIfWA5eMwYUYC7W8ka7br8vl+Uz4Dc3nV2B2XKf52R+T3TeWU2HXlOS+VJxn/0
TP0gW3d1/yMpA5pJR0kTzww3l9y90dHMMtbchogfH8eyCYVDj3EhCcj91LSsUJiw8HOaotUF2Vgc
huc6zTNzCTckE/QUQ3CBYrkZDCmyZiJMZJMWguv06QlwV7Nv1QpWvBOKWALtx9wrOgWUEZqHaCH0
+nkfAt1rL2Jyc2IOrmgauo3G5VqLDQ6d42Oaa/u+R49Ytzn4qvUnzntOj2b9CrFHIHcaqq/WfWFj
40Syq5ETj369PVyqHadGHAoJ/7MLCIHI9Q2NKtwXzJBF7GleKGqfeCTvuvzPVWCFl9dDYeveUxmt
jRgKp67JoQpdC/iPaOfOls4ySsmGsKlRrxAlZ4Rch1MZf0ex2H1gq8Z5qwnuQXGG1hipvRhQSt8a
MiR+9bk94GU94hoZlnASb9HAy3dO875PqGruDIwOmZtC8EuMgCmh2Kw0XlnQNTZi3PkxSpNTOSah
uPtjMbJHPzvQdTbUeq/t4JB3v+LR4gZ9TuPmQFqgXQ7Ei5deN0chsaTuI/mzZlPXXERrixSRRrwi
l5BC9kDbpnYYMTXxabp1IfvakHGyAKss8CsPeibnUoW/0iJv/Z2vzx/3qp/KLXW+/Lbs6Q4f07sN
wi+If6jNg2XW+t+t8HH/26GxltqiXTuIFKPIEyJjNZQ8iv6TmJxK57ILj4QM/sUrC1HziZ7aqkbw
u+mgq+Jka9VU3UjJJ55C8kTLeyLjIcMK+rOBQrSHVItd5iR+nWQbroKHxoTqZXHdUyzEr5heZ7Kl
79yBO5YU0ycqXeuV39OeaD2Aebf80UYxaWRVN4CrSzpzkVSOLsJwOJEm0TMRtTj4y2nN1RNj4gSg
ejJ1w+rDGeI2N7cREDZyT0Xs1MtNhvhaIbkrieJKUZIENTpY/xPOh1EnRyAs/itY3YUGRX5s4EOB
UCZfVLkhcqCaWpde+CrY7WE1os88ylkXYCVF9KpDswcY1EQ7ztFUmdRXrV+GsmK5HMXoQ+aNxH2Q
AN6o8NW3RAZdVBYktaZ9Xe4SobkekH0ORDOm0GFcaVvj4mCSEi3C3Xp62O/GQX/hLmNhC75oDjOp
WW7AAZ8lCH3IqVobr25jor2bXipqYWPfvekBBmY1pLQfFtEFcJYFTG+5L03oYWkf8CX9i2UldhfW
WXjfBLVnvYaW/knbi5mXGL/gaR7TP82eckTNcjCsNx1PuUAhluU+VPw7keqOS3WQdO+jejWhNj7o
kW20+n9ADCdewwO8ez+37Cgo3tUpOiWN2kjC9SpSV/7TJ52yhkqwWk7HT9QeIMr5L/1Uk0QXQ9o7
jXpQfS8w0XYuxExhxpf88ZkyrRZCKI9d8A4i6Xnex43jmKvENVAI0UWWOVX7tRZ7pS6W/+8lJvQw
7eCKbosAlA3bqv4//jGpZYwO1rXqfRqdxTMoUBWMKvV2uVykfDasZ5iE0H2W5N+DM5X+zlUSJlVx
y84FPxUvgjSNNqneu1XWAq4D/vjG+WeCuKxLvSKLAC2+Bl1bFlAAXOeNyygiNJ/qq6uiNfKw6c5i
gan1aX027SYPeYPd/bHCwwveo+LrW9Kmxy2BXl8WIsANa3cdm6T32Sb9X+GByoF3YeVm4OvaETXa
m9LOtLOQdj5VLPx3k/MUcf4IUf6UStM/4JcVYyYHO9GCgk9piNZEtnwi5LoyErL/BAu1ZeIKNbnf
PPBMej5Q2gjJyx4YLM9BohjL5aRoW+Qg8xPlzmVCJnFExGOH1IaZ15rxpf/D7b+dki2eQetpaGbK
Y38vZGD4ZOWIhgYgY3an3L3EjiU1vx/S9WNYv0xzgH2UO2IhrXZQsb5sYTkj5aPEzQqT5j5ckvOE
SrkEH7oSlZm4zr5hBndhpmMB+bJsbKx0ZtCBlEgsVeH5KrNR10HzskGOpiBwEkiUsz0zG9vn6Mp3
UfLN1Vkyk/peSlLliouFINQ1tflDM99T+97IDinajQoYeOJ1ywRNMMz5akfTym/09vImB6gbmMlk
rHlrjtDNYUgF1Dl42ej6W7bV7G0fuAy+g4bTTPXOQjJ6YKzMaSY3mivDQRTxF3AabJtJfZgFficR
neOumG2SsFly0ig56patOPwc5PSrwa/dw/fiIUinrzQxWoOFXZ4DsSoKyF6bIrjl5KsfCcf0b0+D
FwD7/c2fZ0ZWgEbm8TxPIqrWgUPOZqF9IdKeicQAICpDXPrKUFvc/nr6OJ69abnyqSwqdhE6ZIpa
MeogcbC7uJnMWk+T8izF8A185lUSxfpgItByctMsIkumbkvGU5EziK4QLbubyNYOnTgK1LAfn8HO
gf0szKWgTgjCCC5KUEcgH/HOTO8k8JCoIWkoDQ0J+omy1Zx4ceIXvLIPTSvCYGiAL8A4q+JyOkQj
x1qJVTu+xHfkXhW02Bp1FtSxZraPHDhTHIQnW2cjF7jhayk6yeUTx6FI4EVOxifPsc8jC7uUtZDt
VYvJqle5bthdhQRGUWKghe2QyRWSuC4iOterWhLczoo92GgUvAw972tfHnBnQi64gTU16Vg4TrT5
J8UvYO0Rw6BC3tDl/D9e0l2MmuU4xl7kFATQwT2Yb+ry7+FHNwGhyp2qevkkNoHZFx7rDI9sxCVt
ierJX/8nMFVgTZwW97OcqHEX5wCPe1XWF9AczsbqETS1M2UhPkWtKU3C+TzpjFXXQms4QbuZ44qh
HJrnBa4ZyY7y3jOQLu0S6gWu/k7XhYVKdg1BihkkmTbd46TQv7DhX3QAxzIeqcIZeofmzyBfiZ4h
o1/P8bCFgi6566S83NxvbzvMJTyHzO5JTxvlT3pSZJ2vrw+029FfacOoJS7AyblHR/kOBXTs9MTb
CcyP5TLok46j5HNlGcNOuWGSSFAu8NECN9xx19zCo5J+HZZE0P+Mhp865ezo1Ht/N2diYjw+9Fgs
0DV00aXuBVcJbRwQOgWxcGHAQs+Znj72RiSA7+FyC19DXvTvkiJE3zqMVvhXgk7aZ5Axj7FbdmQn
LD5616DoLiXayvSFDxRZuhRKobr1iBoH1vxsJ4Az5TIM2Bt0PLQAmFfuXOKgwalcs4lREs5FAL7D
Ny0gUmuZH+U29oa+TtSLwJbsNoGuykT3n50sY/OA00UY/TyaJD584J1uece8zg9JbsDfJWTtsArS
FV7A2z+KVs43PP4pa2EwTNHlfp5+HGFCchXDA4j06R1e4cA+ImQR7qewBIlyoAhE4xO+Yc+ZKfvh
VVctTIGwigWYY1pvxQ1IksT208GnjDKtCnNx9hPU1SQySagToB43o+pjVsbPeyTBEmB40PFyFeOU
LtpdePms77mLWwNpi62nH0wcsRrQAvOPI9nSY/vFX7XvlYEFbEIuOOXXFPYgre8SqBVWFxVEMZfO
6Eq8QfnrcgK2H6sKiOaGr+35tdf4EiH0R2gFSL9fo/LSkrGAZgH2TWcT+ZhsYrR9Rc5lKxuyuWmS
pfXBV3Z6ZQMYXrKuHPNFrse3enMFsPYmZpLyDBZZJD0/fJk7gPzEj75A/iC/8N2uQsNhx5VCnB4J
QxKjNKPZSnmDZ7YDW5uRkJjbCoccZLP1/FhcyhhuOjBvU6yBvYJqHEO8XndbNuxDwUhBA6FLqRAO
rDsSsQS4236+RUuODLQIbYEAIosOlZTgNpppa3NTsfp16cS1Kg5+R/jXvEStU5/bTbDzsaLLrTQp
bgERb8PUNw/ihMP+ueqdQyp56V3hQiRKXdVFq8OqFKnmV0wAatdrn+r+VBVSi6OHGm+OKAjNEJk8
imTBsz9PYDkzzSVbr4pJNHzQhRlEEwRUt9t3yFNGiBQMxAstqd3PchHDt5L/GkUUx9QDMyPy90Dw
/xl/GleXuwL1QqQDTlOAieV1mvqUOOdBXii/O/MwPheEPBPVN92jCk/ekIdw3arPSeuvnkgqagW7
R4t90HTign34HmMvFXYmNdycrtpRO+RXOz/mxU7ROeqFItqHWfXRVE/+DFhxI/M+Os1ImZrjZHrH
F2eX/yUQcl52jCPZrN80TiO1GeOAMfcYZa2LbzqZl17WjF7ndRhHGv34UB/dfQpnVkrCfQMVsqFf
78JkmTfZTW8GsayOQAdZR5Re/PFh77ij39TVRfWBot75QJq59NvgcZAB2Bvq/U8rOoIrDrVuedaE
h6DDjJFtgdJPb1Fkw3EW4teT3dSDlaXNof/BM102vnVrAfWd5VSDref6oUw6UjDHYjb6THpZyPlH
Jxf1/1vFojTJoF0D2Fs4ab7btvarX96mlvsjDG0FHbodvcCIB1cq4iuRwHDFNFywuET2Vj+uMDDr
y0fmVfmLai4f+VmU+07Cv+BncG76oxD/qFN/XCF6qTqGomFTX+fWGu8f9KK9JuubEuiLf13IY0Q2
PcIU4DaUjX1pVBuxTb7kYdjMY0sR0WWH90psuzDSJD1gwFLCJWfsqkod7aTOHVTxKy+6mgVqdjuV
emTa/f766lrmL6Os/Q6E569hhe3D5qShP469lN5YXX7JFLXJA3z+EShDe1whDMPfpi+PT8CEKjk2
fwPrZ4I9mhKxIGTfH4cuJbSADh0PGD2PX5ApR/xxYzNvt2y7PNtg5HdZ5g5QfXp4WExNcu6R06dS
+RpJMtXmw2M7baJPeQokxSHraQ7Sbg+MzeA3MGY2r1OUPsAfRH3WHSQRrDQTkYVCTrnuhszzrSmj
htIYY3JdAVsl95koJ+REFuWsCw4FvkgpjmQuRviDhqIMh+W+0u7bOpM7yJeM/rNTkvxTQDJ6QBqH
JFqb9PqpSdsanxm9E4mtSNmgGAiXais4JCZo47XNW5Zv3wjt1mo8VKN9MuuJjLSOVDe6f4bN12is
wVLOMSaLuoh94jQOJK50xHDDjraTXbdnEX/EHckGwtj/w/K0lgucDYaDhdN2+43bTLnBOMXhWZTo
kZ0LvCU3m640NWYVqH6jGpURbORoU4fJhJcwZ7Gi9eVJYRDIWa8zoasM1TRXaujq9hUtc6ckreeS
hn12UgL7nbxstYyY6LxffCOtyrFP0efG9eEFrDcaWRkPcq9jji083k0UaHuXR0sbPBEOgVe/k0LF
U9aHZVeUCxjH1nTOiEBMPvtQqI28cORHgvJEP7h00CAWLNe9jFOk13xcj1U48Lj3GOyhTEtDE6UV
h1oLC46WmAF13eV7GGCeUPwwxPXuZcENi6iZC6rt2DRBIWFHLn3+LlGovvnEEFqZ+c9Atn+HAP+D
DiWxgD2VSNmerM5eOdzuP1RuJVkYiHGxPmkmIHioUbwoCmQbJvw5s/rN8L6UvlhCn91ecsY1slhU
AoH8UcgijrDQx5vn87TMoOszas4Xgqb08iBkb55HtWc3NQv8+cIKnm0MnwPiRGeIkzal5nh7srLU
H+HhMZZHQJ41nGoXZ0eVu6zS+eYUvHA77Y6I2+nlx2hx0bhJEXdOfJJIrypsGt5gzhay3A5E78fy
zlfpmmytEs1cFlHhSaMmzy5dyZHjmxL6SolDjcQsspOcsyQjv4Ei1UMpWy2a7sCbJucrWI2DqSRc
mDmdS/0zpP3ILFbLxZEckesSnP0SQZF5hhS4vo6Gnv5rWunfAoO5KZfAj2OQpVwl4jDWe2DjHOjZ
wuMveMUTc0O5cC4/bRz58jH35AgSc35Mbdg8DZQ8srHt8qnkotQW7P4t0SqLEeK75mylOPZFhFx8
KPCqct6meN/bd8WVtCZlaQuEPXR6OqNNknuY6E94oFwhOv6pw2IN8/vOs86OIB6llfmeGKYHNOPR
uFB+FACp8uFO6U7/bvrdy/fmvgP+ioARIyhBg5XGlC2jKIq45UEGK0JkyJAolDhbui1DCZgQ41YV
Ce6SR7E8hAkyx4t/iPnDg/rON6cWjoilgZlFRRKUs2txrW52sjs9IUu0u5FdDA9VpeuEAfXC8uGu
2byEnc38YFB184kWWVj/v8asszkz4nD6r0mnqX50OAWev/eIvyBWeb/SOf+ATFNXtZN3Xy6qsaIQ
U5AdUvb9v48ZuoCvZ2/LkC5Jws+McINB4xewrX5eG/4WjGB3rdMj1aJ5zy1fKqO6dfNHneh1eFwl
fKQ7VjgYy1t3bHxW5cdWg3BNJSYnHKekDuXYbAGf/s7vj7LAj2RQgkganh6WnLwyPx/GEVo1igU5
vDEQ8M1dXQfTd0zB+ciweP7Cp1ZOMX+Js59iP9p4fVumsQO2D7hEAz6zfrxtj0bpgOntvc6/9mIq
n/E60y2QHiFUFLTBMY1SGxGF0qrmu1Iai4bWKXXAtdR4UqGw9CCJ+SpRXmye6iStcHTZ7mbRubSG
DxWkDR+4AtG4w34CYDRx6/HLdqlLdYBQeZjC0e8v9sdAzIEEfqMOpPumgOj4wrE0/zYjX1TUpujd
ygIUC3rvIuTLuODXM9LQV5aOxgpoaDtaScEMgSbh5OE/Z7pO9zqBjm4wKG0a6j3X7qOkapQMYNAa
Ul+5JdYe/jAz7YwTSk54V0QmDhWRjZTyfGqlvns07A516QbrxJVqRiC6Yq4S6hGToDtlTSpSGVy0
ee89PWqcXkGM1+oEqu+n89kbVotAzd5wR6JaEhz0BwC5nRbXXjPtOv8zEOt8obcGGyjfh0lT7C16
mum8MU4+d2KdBPzVqzhkFUFQAaeIkhAUcqjTFe+HLWY7CrIMmEXlDLQAvJO5BwOWIqTioI07VHrq
JHR+BryVY/gKyYOIvnFvNMAPBlXIrDtJZ0dW9TuIhFGorIWMN8hVdB8BwsxijP9J0bHd9GtJSiTi
n2FocM9M1UyJUFXXUNyIPJ2P2kPeT9oeub2sxbRQpyGVnvcxwGZxW5FLgh03sKbU4sshEax1XMfz
tK2LeJeUNd6x3EKNGG9qNmUKhbmd6UZM038giKaDUBT9fxEb9VYrFDrZ/RBmpPOL9ZW98fex7JnF
ICLutTTchLtajkgNDQxg84eZOEqV7Q49Yv3RMz+UNnEEoxKP24ayM56ueHcu6rG6zA/hON6Dxbf0
Unol0NUXQPbaAvWV27jex+1zxaRhOXwEfvZrk1be937s3N9V12tX74Z1gCvl5pgitDRa4AJE0q5D
VTSx7fM2doMVOS7gtOh7yKAZWk4WfwgVEaFrJa/O1Jz8TekT/X3h5ovnzRKDt5h7Kms04InY17La
NwEh0RNlSQ8sL1pO+lUMnUGleE3MhKvX9rXHzskyhuRquMFanntS4qQhA9gDsYRxMivMLm3AcV+V
085D05NdbLkHSNnVa8wQvU8MReytkxMQNyVJUnCkWa3x6zVA5qpHZ8+jvhOphfVnXlONoSIXT+Cp
H4QMLLM3nJHmcXEoFVU+mae/RHBugMAaVHnauPSCy5H/yB9+x3ZvEj+Va++jq9THo/bZF0QZyJkQ
n9zTMcvpADdKclTZ/hL1sQ09zHLNZPa2soz5AiexjYW2vpIUNl+ZjvwGHCHGOMQYi4iFnv+/PMjR
SmCgwJPDihmf/YCTH5RH/cbLopL7+8Vd9MUCb/4rD8kBb9XNZ+7CeI1u2vAs97C4L2Vk3fp2NMt+
cIS/tGxJ038E4pqWncAKVv6HUVqAkg9G8ZSLIvmQYgCSJWpAVTtzb+ntgghYm0n0Y15BZRVYtDHt
2qamHLF44gDW5fxIc0pMzboFF3OZKo/E6CiJ6ZzxVAoZQAEZmOPeVv2u0vO233mN4HywqQIr/A+u
+ck9rXiuIuCtqa433l6Rkxlx8fWTsyab5DSbBBlfrO6Xm8N11Yiq/Nc/nlIL6TKe476/yWEGjLTD
4gvzwcBdHVwFQtKMf/d57sPDqvDjZG4SfzpxPt2+GXDEgEL2so9qjgbxwkfQ7+TfWqaELfDo4/dO
KMKRntrZ7a7X4TCF2uVVZcCHTQvFDbD75MkhzAUD5096rVRkpo243ePVe1tI2vemPsFqmFo74+4R
WSPX1cK0vGWDbNAn1l0VniZjes0F6IG0ul7NTXZ8aBvzLJr+jD/LvyH3jj5FWx2Mri2aakgKsk1U
Y1MCWIsRYSAXVYu0d2+WnEsYnm1+3DqLILQumywpa5eGQlPtD2mh5icwy/GpFCClPvBGhMF20ksl
wz6/sIM+kM8XiftOG4Q2YfMiu+e1JehJb/AbIOM+kRihZNXRHo+oX65tahggHAnawvlChUKIVJms
/oxf/7CnYR/LJPt5ehaMY4glbAdwsy+/ks5VUisVoYiLG0Zudfe6kMzM/EWmKyak/dPwihVxwOsI
2k+XD69yXxuoLyzkXbgHSB6n5gg5onyqaYhoFbHgc+FBjlyRmxBtFHP4pT8CcACzEn8X2pGnnEfy
WDDr1mfSYEahRtcpmZecLI6JFGdPFXasb+h5VrhzFoplsgwGXa76P4urpqaYcUL+zwshcoV3zmS1
04MCajXZY2Cgz1BbMN8lEJI4vj+RJ15MJodpn6c28j86hnVwKy4OYAS0brUhxLgCrwuko+ttxMYj
BqzkOh8BaicX7VZgQPesCtnizNU3wM5RQipAnUNmOSX8sdqFYanBUiSA900QBxoJgGB2WSD0UfrF
di65qOIwmRDcc/qx8KAsfrRZae+BrV7iNBASHjcgPt0aEDf3ihI9jisM+ZWWrdU2ugBsct1IYvSD
MS1WO6U5QAwV3zvtw3rDUfbLg+qyZ7q1b/0UnH78RU53w2PiSnahleW8rpkndbvcdJV0qSuTXRO3
yN7KEF+w+/pq71NNqmdf3lZDwOliC3IgCfSjtZn3GknerGpMB8ghTyK6Qu8Vhm3MPsc3sepg9LJN
5TkpoGiENVP3o3QCB1nKCufa1N5esSoIJV5pw8kWqyQRtzrBKKY+RwUUcxgiZLt+YoE1Y9VIfpeb
DQolyQkH0bfsFlLd+sL11HCY2siLT1uOqC7qhG363+imXVIalnOVnrKNRM0QsCadXn7DUiVG5pBl
lzIwKdcPyVI3nLXvV/y2oK0bA+89gpmXfI8fpO1MT3Ni2p9mYsYtIPcfIf2y2XgakV9WyrMF9jq6
hrUrtrXzKWqDxA7hgOigJ4bk3ZNplFnC9JBF8Fc36AGGOVcgTAVeKQDNxfztn/SLGf+ldb75fvdI
rnBZWF9+yZIc/3te2PWWmNFfxjqgERDehKnovLtxYwEUvHcJchJLFGZjjWsXpkVe9MTgJN7uNlDG
SQ1DfNTny6WW2o2ytTF5oRHu26Czt9Tw6ekf5l80f3ej5ipb6oIUEPfuwTqFoi/LUGd9+fgrA/ar
erSM5l1qTjAaNGKKrmUfI+vefP0qxN2G5yBcRCsmV2PGFDVfsSTKS52sC9+2LP4jtkeY/aX9KT/4
W+agcAKtacF+mX8NakAsWd11BJl7ecc24XTAyBobwfKqcNVGb281yjug16WjZ3bREjDMvJOyiWng
qShMGt7BVjmVYcAyKiMFerc/NMClyvV1ho8spaKxZUEiT95fgkVpJzigL2Q2PL/N8qBUJHK7irb1
XYznW7P7BRd8ElavXSgDVtBmsi/Cv7XrnbVSpWDLYnBxY83R8wlEb6+zAF9S+QNM83plHpjaaFUc
9buUBbXUU66RP63ixe/x+mkX5JRvCQpYOPFyASgbnMCD4RiaFd5H+wahfi7YUouNw1kV1UGm21IT
dBv/2nrRRf6ueFidwxc/gP1kS2YXfdoXFw6EthsTHXWea744DKfNi4pm0BNpWN5kJdbygzCRRRC6
q3iyDABvydAxOWHwWFj9vSM1gCVJBkDx/HmejJ42b/tqwCdV1yvEyUl5ILfQq3orC6rKcM9HOruq
h6Lzc9J+/UcxjwoqNH2Vmeocfx/EaNaw/GewLQSYfiLrR2ZkuRvEX1cRPgLJCB4Jwcfl9PsWHz0h
ELeAyB+UPA0D9bbIDaImfgi5M5YTVqm8vRtgPr45A4ivCRkbFI4lPAVdzdWcatAT1oUuJ5JuCd8C
WA/a/zYVFbVicAnnUQ8WfMnljUxy6cdT4xwpRDhU820AWZkoALuIpr+TSiM7b44rbD/h5+CZWjXj
uvQQ65oMc5KLtX6KOUZMInY0lKKIxuyLv4oRo/QwBviR6l3BVq+PKa4ylC8VpI+iLo9GczS2qNMG
xc+p9F6zjZCS6dY6mv6KQWvBhmxb9SvOhFleyFbarvAnE0MGsbkS8Ku1s+1smlwM8hUJEC78wfFh
P8lj8KOfyT+kI5dZVJNq3/RGiAm9WKXxJ3I1wBw4S9eW6pzsXZd6Rjy1JjC8mOKxQifR/FWbmdy4
XlCqjKfVm2rH6g2myA6NUVVFb5vNbnDwI78Czlrl+R8sVabpq8LKd7Df3iXrgYASOPlG91qMcCAf
vpMxSWjFDmgapogj7MTrypBvIE2oigX7mWMXGtk3VhUcghksKW2MlW7uneDHV9tQMFqNQr9h/ynu
QKAyQnFPPHmZ4kooHFKfgtJNyzVKpI68AUrZjkVYsURZ/1CM2+8gfrlcvGh5I7BRag8oRO1T4G+e
RIrwpsxfy9zvjzQtFSPyIiNt3xsXu0esL+9qHec+689DDloMeAs4I0E+DVLgRVYCMp+6M6sG4b7F
/MTcp3Ac3ceaopSmPjcuTxyis0BXQvrgz/JkTDRdCEM5mrqe6rTmb6tSTN8EiItHNY1FXN4zbfhU
nShWafH1xtNf4FqSfRHvfZS0jK+pVwCwHGcd1UuHVw+dRTsD2g57+PQMCIz7Uiq3+5vzFdlW+6dM
zmoc0LxCNssd4j1JgaYFC+ixl7eN6bdAonqiDvP45+uOMkFcUUFz8lBMFyWEvXqavCtrGXSDgtuk
qv0sdk27ZwCERpCAkqwxKkQ2dvm8ym7h4uRBht92y2rSERPMUJx5ovznoPmVbkdU5EZzNMswWF/x
VtKvvSIbdqwtqGoEvqEd9MI0Tlw6aLlHMXcoF7JMBIKytNeOL/iNRgTtrmaKtLMGcZnlyX6Uy/V+
g5ZbFxf5eoKkehQ3pFWrEVnID6e6kNco+te2ID2QER0jHQALhYcLndEtmszqvYZn0u5Pv13fk+nh
gtcBQKi7v+eF/++d23Zc0xm4nfN3cjwZlVpbMX0U0mmC6jP5Tw3hsJVvxyJ7/ZsqNMQa31xYIuhz
pPj0M9ygDWIXpG8Uhoa2u2Rti67QwNgUWNj4SFg70RScODxK+9DwMBSsYYxiOQ5VGC7ciGGMm4FR
5YK3/OEhQ0ZUpT0asZSvCIPEKkWfB/o8IE6yqkwgt6LvQYPf96cjFA4VrA0/c57yn3C3EKHzH2Qa
m4cJw0j4RU5p1TdCtFDzqxFYjec+vDVcMMOBjgZbgIKkEPSkb2x9lxWAYsbbODc27eASwRY0Y+Bi
sDxVYHBu8dkekQHfVx1t7QflCIhYiC5ys+r6D9C2cna0SHYMC0vp1wf3ahuoh32x3gazXvF+wREX
Uq6xoT4kDIMnF5VyxnGCxdOfvmxe205rKg/9ElefBOCdJNfxqwP0K/W08TCr3rVNFpqX2C4gR/as
Zjklv8tSXHsf6QH6rojmkq9W7wus1vLGVuGFtPkimH87HoZuvOIloBMk1kV5uDDm2j5o10C7L9sE
kTVNOHwkzVFbEWHilVKYuOVUfLqyfLUHpN4AetmswmxLey/g/d6IxBtELfg/OVAVyvomL+Mree5Y
bZxzEqAM0upORRDkxg3y3qpj7PcJpnktx/eERVyB8IhNNbM7rFKhQpa01jaO1oZOJg098364GpQb
uODvygDIpixRPtqL2PlGuKest4fU9nbymjKmqcQH+PgQfRQG4jfq8OysyDwtZV14ZoSXwWml0gCk
AS0idTsx93xkIy/q3rTe3yl2/q1B16sg127AthRJxy4oQoABmi8L/ZMcn2gRoUo7dnELX3FfuTNu
J0CQnUwLLVinAv0VLfnbHXQZb+RlSgL+/hwpbf8TlgY0OGeN2OBvO5YiWOexHD/Y2T+Lu0KZrTHj
nZJ/7Uh/hClyaleo3f3DHkH9XEYxyTM80ZsowyQgcFG5yNQrZtWVaz3h2SXlNtIjp9JIoBs/tBjF
XOyzrGg1nVpfosSs0mD+pbL7L3GoHCb9Ffs0vB2mTZt1rpm7EwxssLOCWESpkcwSLzlIxB8SYX39
Zu1/U5bnOKN9bqI/U7TRs/ijAtGI8/HJ5ye+jkf+bZwIX7byMxfVR7Tcs/h+c1D5WYVib6NCBswC
MaugYo8q72PrlOomPHPTOhlS+c4WyhS2gkBVTIhFDRkjwv+b0Rfg/7YQ7trUJRRwBlPdmV7n5/ZJ
8v+kfOsNYPd+xwm30guZJScoP0koM3ufEw9GIUVsFJ/cpkr72rFLWj7T/eieoE9+OQAfE6W5/0w9
CiIYzxbd83DSE45l1/p0Mm4F7ZPg9lVsN0VW9TJ4wn1k3wkA9HOMzQGSS7+KEq2Shze06sgvySwD
eG8BnJNQ7Vpou1rq+T2D4MUW4k0q1Rq3a3KAsFfRKrZUE4Q6dVu1kAqNCSTSFEqZ6r7ge4c6yUQV
8/pdg2btIFB4fZf9CAS/QRxbOXomsYcuHUeyW0bgEnaMPLCQUxLHPDoYElK2szDqV2SHZUn2CcvS
mAHfyo8Ji/AnkAmmOyYTZ9ERwwQW0vDcJaSYzL/A4yStEFJBNKE4+eN4xAyKIBAtbTJgNCKmh48H
QneJuky9C2mJb5coynkN0z0hxSzmdYK3mriwJgcEXBUAUXiRR7cVa+GA7luR0CsB5O32MmEA5jrQ
7e3NDVR4wdDaPSZk7dIVVRZbQ40M5p3svgNtv2iZmRQRAl4IKqkYxEV9cHZzk8l6q7lwRwkVhSXm
GDPBFV2rXsKHJ5Aeg3BXo6xFBtjoyeMSijH2B0sE0b2gQer2qsFGtOQXyHjLVgUCc4OqzxX4PHBP
qTF2jOAXeuO66m3wwnqLkcYmxls3rtg94CYIVgwq19n752i+SxkdcbU9MTTnFxwHUQdftnQqV6ve
co9QCl0enwZgUrh9a4IGKZHhLSDb9NDzT3wYUnO/W4IPdEeFCGZe/aSteHtHT8YdJlDzSwu3+KEh
Z8g9KTaFXfe1Sod+5xCmkj7K813qjHXSY8sxtm6UGHuugJKXC9ZRaZdk0CIP/5emd2BszIjVZ+qR
yPvLEkTXpVwYy4C40EK0H3vZHJ4Ct2EGSckrvfjasHRyS1dZjKIniOnyLJDZ/VYL0kOarZckRdXt
o2YalN0uyh79ZFvmL+oyPweBEGJgX+sOZXvBnL/6b8vOrlghq5Gh4itqvGVmbB8iQc2uUWrDqbsw
O7uNyxnhNFU5UBbgmZIZYM3ZDgbgqN/qmvffVhGG947SzIpLT3bq2htxEW3c9Iv2Iy5VAfx0sSux
J8TJX7b5fXJoXt5jTYzjh6VyzBtrOn23zlDQbB387PA+8dv5V/tbiq81JCXYc06jllxvbqGTclQc
+dst3gVqJE36nJ3CyVUBcc73PbZy4KoAeKRAFJq0x+Moh4XSsq9cTT2LQ4e/02p+Jxf52PM9OZE3
SWzkjwzIA2jyRiOUDRYrCPA7pi6eR+FPbjNcAi/CX/Oqlld9vDq6E9TSNIzLbNLiduwaJ2dlvRmE
BS2RN+QWUdOASq+6/2m7wN79HGydAEU1nkk980n8gmzoNygxOxgb6HuW97VVLbqU2+ptFV88b/0a
9aS1zZsZ8vxl9uS5b3ZG3+j3WZaJXFJWY1MXcbRj2HIDi6urYzymnRMETZRALEnfhGHL6SYmiYty
D+uHUqkPPd6+Z4maMLbbMzZGqdiKwSxGwWmJzyC56HwXDMB3fIaFsUd4+vgfgSFOif6MeHVOYL0g
nK1xYCK3qHK1L4KF24RBf1JVbJEaQCj5yLfd1aLW1NAjRZx9jJbKSsZRUvFhDGg+qpmXMJG/vGrO
cpEsafEOFxXg7pbu1NTAiEP1bEyK1S2YjZJq3JHp3WWUInM3piXDPN2nEdtKFa5GJZZg4gwSmIKu
Kb/+wVkSBUA065UQIsCSzQDZnmy+RF28XCqOhFFJByj69laW/tpC4wIZXGIIjK2zOMNFgTFtN9ts
lk+uu6OUS3NdmuN9WClk4ASo0mmNvMslMev5qOJVETT1ZqnrVcA5bsUTFCr3MxxZGVZl1+yj1+u+
WwYvfU5ukRZ2aEflLzd5afRYesklU7DoXXM+/x2vCrB3ZD1jMhA7fwSsrZVBdn6AjwYGMXZ3TSVI
HQC7hKBzwsIRvT+1bn30CW6WOfzn0mjbEpu1XICpDp3042n7wVl+7WwERvuHsvVl40mPTof88l87
lHYrwFNp7IPieQlti5tjVrnTTvTldNxF0+pR1erg8tMMGImUXUdF6hCGK+ihvUXCbhdoonKS36CF
QVpMMnseNHQ49qeXloJOV+YjVKvtsN/hl1xA2VugkzBsoPRnWlkn67BYKBtCP8DVnAeItJ2hGa1G
mWqEj2Yb2KPpamSJ1EX7vxFn81EYEKp6U1svsjSVFSDaTb+6Eu5PPfkiVtLvniQ6D1Wvd2LgRyKX
AZ/FKjvZKf4LDunGQOa/5MC0rjB7LxLQ8Kn4f1KXkum8yZA36SUIzt2pUlelVdJguevLEPrCN9dH
h2BrUz4WVa1HMewt/HoMTO9UjqVmctQV1a6ZbJn5Lx6btNMAPv1OosG1Km1kU8e+ORwcIiLv7wZW
+cylCGJHtSnvy+hqfvYMxNk3V/WlRrkSj/xO1PPSRSeAFZaIu5/l6xjLxwWph5Y+uN5XYafPfgca
X3o3LPk5bG5fk0KZGs/fMD957JJa52Hu79eN83RpfSi8thgliTFMann6DYe8LUuITjyPgN4U2JsV
qAYDRtClDSESDqjnJNMkTZiQBtMkI5spO2O5vf7y3tqBf3ogNKI2Uj82YK9pSbx1pdM0MeVucPMQ
CaKlNTLrBNE+ehKJOveGZsZLwVNePAXclbkZNUnmqUhl2GgUWi2skZDK/CRmR4OwbZKIesHFSbYS
3KE9DxDB4euSldXejpIsFza7dO2p1sjKteHqtsaTk1RC+KzFoYcxBLn8tA1pxTZorjbpWvXM7Ctf
k40aUSJtaaEMgI36qsosdYX2/NkmpWD3OkH9A0Wd0DFZbJ1lqzBO/jk5+Uez7dRV6yYnjX0yCW3s
Vb014W2RBiMzZtxcpKGhCDo5DY1Ck14y+qi0sqCIdDhTLMecvS58VzQ7eBbHx7LhiIszQgZywAcZ
oK0xvK0zkmGHYy8KHNKg6VB6bTNCiTvEGrosqPu8CkypIBpW8t0CEcrCw3xU2OCBDXnhjJv4AOfS
vJW64+IemrTc0WHCX6QEChNwVfyf9KSo2jrJ4lR7srRM8V5ghpz2jmXd0uRR7r86ksInVbatl8/A
f+aIqUbIddZ4fe7QxKKdM3mHTNcnlzLFLYpXiVPEvwkmtQdU5liLZzbwFiRrsKQiisrZ+f3xWgVG
3GcOqc2kBErQwknHzBYTLXJsAwSzYwoG+oszvXPrrxP6KpUC2LQp1T221dzV/R6zyyqj1VLdbMKo
D9LcdGBBw6lRwCpsbtgo3b8IS3tKYiZZN/iUiUoZg1EkO548IJymHAJWDPQInx6pVVNpqiqdGA/2
Ood7N1S9lnBAOJEz36vA0QCUhBWZZnTtQldbgnm++NC0GkK3J0q7lhsrRO1JbagIxpLw7i2QjGnw
NEZWNZHcchoqq+U4YzheiCo3EroJ8dQ0cPAseqYTVVf4ODcmygZE2dG/j/e34/chzSh7EQLCD6B4
6S2gvh/KWPHtkT1xk3PyOlURF/fT9CeHWgGJYS7yKXrtTGnfxcC0egzcWH/2LSFamIqZdXyfLCSp
GqF1X8LfFuZOuRmuWr4i5r3LFDHuKsraRgIDLx03Y7QFOhRFWI3bhiSWlHvtr4n/3esLi3OQoYxA
6UAvVW+nVldeRRJ2syQQL96Ne5ho08MpiTQRLgw46ZTpox1hBJifhkl9cr2ReYdxJzBSJlPQ/ZEo
r8+in8guQwSlfBfja/a6UI8w4T6iTl2bqYYewpENVohkmCheg6d4+ne9RabvqHjII6viV/6+dmyc
ig0uMmZZ+mMJt30z0xbvQwTomAtrw55DFNIOE6SKoBR723U3CWyheo68cVJ3n2h+84hv3XaiLvuX
LImtsVBwsCWK6EYmJREYgIY3xIEd+cFwukdWYWYSFBSiQaPZKtUwMMGQFoMM/0IwXOxGElh9BU4L
MkwR0EtSCSifVZgTd1acgoejlHf2FizDmqPArj2YYP261d9BzL185TCf3aussgqQcdw07MYvELPp
cBTBuwmJp6CH5IdgIBb3b8PHbPSdML3/LQDHVzn+4X/+eDDqjrViNiEDAJoavhXb86hSMp7375Z7
17VLxJ+ij6vFkHcrkVJ5lyCPDDHAGCPfq113fVW3UiqTqypPp/zEtD61poOoNDJzYtXuHQqaHPAL
NzL20SEN+viOFauCki8oiYvZWsOsOvxPoIcoKCFFyMTD6kZfQNiOlAVyYpgx6tBqveZK0aTK4YI+
EwnEHXyNOjhS33flszWoQ7sooIe9nP4RqcQPhKYLVqOlccYXyyHypMrkGQCJM8onh6PElp2Y8MFh
fwgMNvxcGA6ZJz1Klrl1B7qhmhryFI3D095sZui9YF19idJ2L0w67i/h9lsN/1t6OD/tv2LmSWrR
aK4BqLEC8BBm9lS0wuObIkrxhCZHOBAGByJUWJl8hVr8MJdfFz2AfsY0tTL3VwV0TGQmk4LAAF0Q
oBALqC38Mc7GFQ6D/cBM/7NSx+B0Zy/nww+w/beHEoZC7ouWj7YWbTBVCPoT/cIaq4hXooLAb4EV
T6OsTShOSxH9H7C0wmu0gbVtEVvLdwsyvb0gVMX9Ch/htNmr4JBn5ku2i/dHBlINDCjgN2kDQMh2
tlG7IyHe5EPTEc4i/SU+oYIM0hMDfMzMfbVDrat9L0Kldsk+yzpJTRGK+jOrB/NXTBr2qW/oZLID
JqcSgpOm0L5BR92Rm5VF7T+Ihqhz9OGd07b8dkGCnUoQRfKI4OIQHYcX5bnQSTCHIgEL+nrK1DuP
qhkzP8Qq0j+b+RsNu2u9jAi1EkFCYFRtLksLV8GUNv1Wgm/DBYQGpHQ3UsGwk0Hia5fKeIzPy1Fj
gslXPYv/rlaHLUQYFKjJUIz0SWlfgzlfEctRiRvwzc90zrcbOiW7txpMuNO3KDuoKnxMgy4METB2
+6Xpp1qZ+mAzNC0pTc/x17Kq0MJXd1JAbOyHs6HRRSywzS7B5sQKTnRbiuxO5y0KtSTIFSm2ve6E
54cLxeMBrtlFTRr06V/AL/zIaCdwltO3Bx1IxKO2ArbXTRqR9XbifWYG4BwYNp6AwWuU7GoBt/nw
gD0RIFMDbKVRfVPWVgM7lgdzZWAYabXcQBqhGzHte36APb5+ptW6Ga+NMEQmb5tJbhDipRoGkjCd
CF3ew8bSJCVDjre/IXyY2DUqL+U8SpxaMgJSPTdRl4Xa56Hd77pbOl3oGtrq0DcZc153DbgQTKLP
YMR3qAB/T3F/90xaEDNeYDNF60IraBd3akBk6l90KnBlygufKCfOAYOgd2Vv0cOWUVHtEmJbMNb0
Z3/B3qHuyUe7QbIKJZ5+yK/R9kPSdJqhqB//ShwAfOG49g8/sXFslZl7lt6ZMJk3EjZXZx817P7D
dTsX8hwBgxDUtC/g2hYw2cezfDNwUvX3BpInB+W6y9GCL0vZPa1dfHFLZ2PmMG7vgBZH2SI77eUQ
VhbhkeoHipr2JpVau7QlmG7VT9zOcRewC2Myj+03DkvdDRC3/4O27Y28RwCLFAYyxdRIW1v1FHc5
GzKALlP+TlBSM+zhzqUvK3SuVy91r7bL8oEXJi6NCTntU4NryMC+K3mJGvaOwtYJsI5bje+fORV/
WQHWWeRON5IQ1dZn1schsh9/4N+nz8tR8xsztEpAJuwg0qTzg5fHPtaNa/KEJZCmvCrOskIfr8N3
F4Ghak9V5CGiy142UMgea2pQRa88NRRJY+CDaNWdpyImWZ/OHgQambOdsewxSPfuWAFdDj66IGSX
jN09ir7gGgLnCCSqKn0VbqPEprf0qx5/jeujYeydrouc5PP7RZ2iBG5VtbeAzMbVx8KkXGyWTV/A
Eg8cq7W73pt9wEpoz1wGA8fYLL0O+GEaG6lJB11jR3eaSS5ZZ/eX9xtGkm5y5rW8ehSlH2fxoa4Z
JVWfGW46lkq/9YSoY6EpmUjhrBt4A67WQzOl55JEWBY7Pee2GceyMzGoVNP9KMWmOL8d/9EF02ev
/oxLR0gnAg2sOhGH+wJ2LemBqnVkLPy6uOpsE8TKljhIS1SeSy6NhTz2ni/uvjUoCWzAljoT6Bcs
8pmLkj4hT0QS2nr2xTYUTyR6wWsrmVgbGywVEs8IlahGXyMMYUy9gcck4mfyO31tpU1Ry8/Fvqk9
vi09G+rM0duBxdWlneIMBLFe07LF962jMFLM8fEw1T3aqtCSBtEa/JRHSkJXaIToLOeIcB5g4pep
MO7piJxuUlb8RnQiVW5QoaSwU5q+FW2GGdQgsa+dFcZmRpRjqZfaNAJQP+I2o7ln6brEzs2YjBYq
zeuZU9RPADJEAgZrI8VcGjZkyjVPqb0MkFziKll52KT59msJyoTuOc567AepXQADq8gi/odw3wys
7pxr4jmjCmB1rb8F4H2mdgrYSe7Nv1Tbtyhxxoh9yi/yXqfDyTWO32s+kug4o/DwUYXltPxtbjhL
7b3vhVEQxkd0SjYXVeaxIbU4hRenO4W0AEPgh/S0HIs2RKw08n3IR0wempjIpaP4cBR4bEXGSIdi
df356L7tVDpOxiKt1FoYPZ/Jf4/Gigiy3BGdHN2GVqEk/a9ujQO2lMbPfNy0WaTlTedmuVJ/Egp8
F9R4NSgqIV6ySNVimH6vhZuPfk/A+HxeunITz7rS9je4EY/Ru1KArKcTCR8t0i7VhFx//NGftsIh
7xK/RBTkFbo99UyHdxUmTMg5aaJJJP3qNoIlxtrrFzT7MHLgyQGfeBKS/rF9bzDOT69yFbaBJKQ9
KSk31v3aZ7kc/898nsYdD6r0LEH1Y1qmy1XvnGrs7dnVO4RrAuOcy7XEfyCtIh/3+PeY5nF8vYN5
afulTArgO3Pr1zzbh09ScOqCGFXyHODBlFdxcmgQpGp8H6grjLj+I046xlx9BpKvrufNgJzBVtwj
dL+vXhOa18K+Hh2iN0oYVB8EvgAJMZH62FsHVWjWXswFMLR/Po5XmxyRAHsY9x2rDvuUJW/Umkmq
xwvnv0FSzddS7brM6I9Oba+I+BmLmQTEBaul2XPPwfCSvf9V2j410SdDI81hOSKa+OmSrE8HDdke
QIan7/vr/apOo/uP4dXRMWL1UZ3mTufE1GGTqTiD7IwjaV9KLcLfQ07D1zAE3UXTgUcUAbliMEe9
nt4SJNyvanasJNfQQJRu3h4E0u4xoUQoHkil15Udau9FzBMUqzvmb2JJKQuca1C5gJy9TLGPm4X9
G/kYKF0l6Vqq9t529Wq4ny6eViA0vuZxSr7v455daGzM09Z2oEiwjgG7yBlInU/eJLV2eextSntG
0oRIbQ9N3I+eAN5DT7P8BIQKou7ZMHxmsISGGCIeFxX+5o1nS38NpDUXZXRWmtkoIaEuAVIIdjFY
aoecnAnVJOdO+YgGqpYpJiwelaDcwy1DcfVnDmwQI8T01V9E8u12ury3FuctUaktr1zlPUcnQObk
TMicCBKqqdfdk12F4MiaXm8d2Gg8DQAkX+MNVRbbxRKVu7CXf/DTzopRLEf0bbOr1z0uCv491G8K
yHlx/XXYFMwRhDZfHZnBNCtyxGP1zHUcuzBkg5VmkvMLmoQmcBUgK3hYfKGLUPE1MB4U9gu8Fk85
CCmT8PYAr/DKySN0uWfemlUFzDsHY5Ome7v2TSpVnH34wJjEFQWPYOBzjbZ/v/7SbR4HkRDV6zJt
WAluyaSKR6CdJYbhjUNe+FBaEeh8yRLdFC6hMAk/k7De+eQyHLxiCl+O70mHyLOl7lutY46ZZZQH
1xhQddZTf81bv2fOF5wO54YlmKMkV5Qdw4OuO7tbLq0xt7AFaiJeDz1e3yA8NHYS0rOVDfZ1P9EQ
5Jzi0fIiXflH/w5z1dIS4SVhfapWBhn+OsTzjK6GmuM4zk9M4f6e3FFRe+3dhdTSfBO5l8SB3Kvb
gyCuYbBnSYjuXK5AJVyFCULLWQ99q1oZkreHXTIuyZNiUC6TfdqZP1/jdO88pDC58pciccf6smLO
ICaiYsBJlikGtlQYaN/9Hchsddb2lJiR5bsbHeqN60g/128BVPchVR2j/UTcd5yFLB+Y+4Gvl4/i
Nhucl+hBK49bvxVmJ62yRd9u+8sq4f6pvOLh07Cql6yFoLQ9y4zbI0L94vpK74dJCxTR4rHTGS3S
NlIbY5fVXW3fRhcO7v+1ow7LHn4csPrca8N5KRdBc9zuC9od4+VX+qqOJXxAHADKj6IgfJds7gjb
WxRm854RtdHukfrJuTzn3pWoK9z6WgwXY7HlQjCv90cmat/jytshO7FrunTvw/LUoBKl5MWTo+fv
of4XiFwmjiKaZyA6eC+xm6+7dnpxL3Hte7buj0Y43/TVxNuHyRIO5PknqXLYL0l/ngA4dxVglbvo
KBsAUw4QbqAFtpZSHsnJNkOBfxS9kQeaq8UcMY7xk0wiUTCl7XSLHrNG4+WHCJ/XtE0S57Oij1RX
udLb8tVn4eznq+iPxlVJnduRIAJgxfJCphbZoAcF4NFYsVfP3rwI5TSAPmSAK88kltrVfXrHB9Qx
r4NhZOcloy/gRKeWm//jgmb4cDPlYbb1Gk7yNURDseW5OD4BZZHy63JDdhHY6NxDZRUtRHXw38qd
5coFb+NjLFM9tayGJdRClhw7QgdiuuatbFx7AmJjTcZr3b6EOkrnEecu2ndJzfTMC8wszHLQhfRe
1eQYYWzIG+vwFWdsdEqlTxpqnafy5blcBTeohOvEnRVfcoMaW0fAxnmtwJ0SOFVMqktzyEGVGcrE
YEPi1FIOx1UrPotij7y/lGj/Pn4dPbkXKm09dfCRiqUAVIo6jXAeMVPCgrATepiRVElQWB5Avqm0
KbQgGvE824PVVfdQ40v3yqsPY2WegP9BFVD+dQ1sKjdQ8wc/8HdP0xvykBm1gUI/wyqbQMqUg68Z
6eEyu5GcAH8Ui/k6u/fnFIV5aZeg9htezw+o5/PAXhStb0VBLqJfhNI/v9Llqw9Sc1z0hXX8cNnS
dmDYBhBVX9P24IMP0hbRkwURLuNzB7FszRXBUAc9doMOOvXOvtHkxm4Ml+vL1MJ4lLVwXazyIN2d
D2BHHLZ9kjEPbNzIIkc4wWOQsTu6gDEV4LSRDEmlIoN/Bj5e1fOZK1lApDdrEkyMn/62hrxZyCDN
4rN+Jo3czuyqo77viQA5eJtAXPfLTb9nDcJzatAJ3svK0H1dKHy7oMjOaPhoc7bZcHjnN0wRblKG
fbUtVlDkQI4zegd3XDHWkzGKziI9KzTj1RJIPvjNEvIKhixptQaO0FQltQntHWQkQwBBb64Cmh+4
WsQqKO7SwbNFbNoRDt2xlhl1HPa/CJLVJDEzwpe+OnGd+UfoqcJSfn0KmBTYcirVFHs5Qons8xpE
nk1aSdn+btoQ/Q5feNyqn9UJsMnD40HonwolxXUYL9IwQ+zBliOSNWknE/eYXeTkHkAUF7iVpqm+
2koeAcLPUQunbGkLpNZoySjK7iCSM+K8angGhTa6MhyuPXwqKeHkoaMWI/+L8IORzfU++DTQCwzK
Rnblfbf0nB2aINFAACQIVHmQf9F7skbybzJBxmnONJmw2Z9hPxPlbSd58TBwdCXCC2xqe88GSqTM
fckXMzrMQAup0SlrPj9IbifSKH+nWRHzCmZ9agRMGDGgmJm2JM9GQT+AVZMJ0p84kBUZDIBIxsPq
1icbspJ+SP7TpY8Pk+6Hv/Fi+ZvVfJlCIl6d2ZenBc2HJNL3hEO3T49GyFIHSFfoxMKbnvg+rOp4
lb9qU/BMxv4m72PsstC8Z5Jds+m+v0vWzfDD5kzOyTGip9UKbMR2dKpepjALv2MQz6K3R6eFn+cZ
0KccL+RhDn9GJTUlItttdTHdXIcCKvo/LTlzgNO37lP0KwsU2/igbVidWKd4m09Ooh0CvarHmdSV
HUDfvSGr8EpC7ezhqTlSUxSkpfJ9kHohZVpa0RodG1/khyB7VRMyCyf/5fojStrcVRwrUW4RUg/6
oRSdvVTu6h2F/jiO+TvzaMiS4Rx5PFHt9um2z4eW+DTCypAK4bJSZzaiqf3cgkr/AOP+X1iSqx06
pATHdXD1l0H3x9qUYXKongz5OLcRJhJuwfD6PbT1pkR3ERb6sfnOduH1O/5wLlchqAKo7R3657tI
tpnGViqbkHcjQnrItXQ3DU/sH+cYnylaV/ctTFOTtbcXKXWI/89VV2cWOKM/Z0FMTzmABlnrLajq
s5MwSH/aJ6WXP0jTergWg3Gh7dUgly0mGS7ml5jD5LJqf/nx4SgdHqbZ3vWXjpUtn9ywkYK/tP1G
IgJ9/FpUcAnrOiUpNQIGfn6gzWUIh3NZkcNSk1BoWSNv8IDxAZew7hAOElNS1jt4qUR9oBT0cB+B
OnmWa7Ahk7PMm9/JKgcjIRcMbFik3pA6Zb0bljyo/pKz/ku0wEUEAgP2UQJ9dpMSh2i4bYGjdYUC
0d1vqqf+/jzjUAm81ZpP0fpQOXLGe9HIDHScToW+EQH37BN9APotn4To/zPprxufGZd0MHeQz2h8
OYRnWd8TSMxVfDsmwwzDzk9NhRHgSz36VO5NFuHAf9ifYybJxiKRnYfYVH04/7Fl9v82KY94vnqP
hwe16K9YeHFrV4DATXBRUXPDWqrHEYV1OumzPUtFYzk7AyxVyh3C+k13YyVEns+cX5i725QvieTL
QiKlkmw5BUhPUQFrTwoJJyp9hD2Md4RtoDvaHdOuzFTjGAC3MrErZrs3BdPQmPDlISzuTrjvojBz
bLZePQ8qZcK9+2nUcnNiYcmgMFzCflwq2mOP9d0/BmUKs09UoXng/FkBnzP12JTKMmAes5VpjsYp
EDFgFURloXQYQa7JmSrFR8n/XLU9UIv1Caa5gYqfaOAIxttdnMtpHN7g8+SrOmPOy+2mvcFFE8VM
jAMREhiIR59R0AARSwqcK/dswZR5D821O1KxsRV2Z+6klYfYh7JYSWPHvYE17h0zPturGYqciljz
oQU4MM8YK9WDdWxFypqKNVE7S42g7tPSbS4Ppci9MTLn+9xzd4Tp+XqQpn4qvt0yaCOBRxY1EG9z
iXyDODTCQuAOeZNXh7cntGuOeNNqDSuxF/vH7ZtrpeoCR77FJoMoevuxnaZ2mB1XqB7VOly6pe7m
rFqBYaE95mXvHsGF+cCeZxEjxABtco7iDyEmt+IhOdZnA4H2aYyFJ4pFGI32RD31/iqaWOViJdvY
L7Nzr6dX3x3N+DBXLlSTCBAC+ExJRyQLh0yiHatQDDLSuB+2DXVYsEjm0/0piUDqWLqzQIvbA/0i
IXExFaanVAWc5BdPh+0TAVICJSJp+ATAyO0HbjZqQZ7B4OVVSnD6QiUVD9NnHWDrX/HA5OohxuOU
fc99CBH6RK1zIMlAw2Uho/P/njlA+BtU1utHpfTUfqhYZL7rj+FtB5iewebsRUZ04GFaY0onH/jQ
unBmLSUJc6+IO71M8tXyqykhliO1+dhHmjCUT2W5gj6o+KHq3GUmwGtlR27shRD8MZzeVktIXNPa
9uVr3aT54VrZrXlYHm6+rn2j3j6/8NxBunUa/4QdvO4hkyOVP+iiQwL2fdOBScb3xY3x9b/j5sd6
4TLMquMTaq1kBlCBbYau7Zo4Sp96mEy8+PsNYMlCJ1IE04zjUwgncqRFZ/m8QVBmpE2jrlYdE5qa
hAoFymUnmnEb8CMIR6x1IoKRQwFNDVTAJicJi5OjMm1sV4q+m4IouQvXMDG0XK1r0n5VlS9/RnW1
UwdOQMsgz9i4iBg00infXtl8IVeglKhh3tggjY1x9gphd+keUyRgAi4PDTzV/zOvF3WBZK+3FEAz
bWUtT+mX70ujfPXHHdDwmMWs+eVLByiqBSpzhkjSEk+zlRmejtJmJqBRorC0xBBNIrX7ncHQKv4o
MV0VZfuXnvhbmbhlqJUlRTDzldj5M7fgCR/DWYkw5e9+kWgJjkvc4E07kfjyTVtY7Ymy8P9hZdtb
PdLVlTGC4nd6HDKq9s/xNtazuBwKUXOujy5/g4Nb+cdlr+803DaoByGIyR4S4dGyb6Oobmh8dB+V
ccT8xnfyAlIKJ8xQPqWT5DrGw0UZbdHSGLDuV7Xn4CgVxRvzCktiiiVvvTOyXsvnR9wnjoKwQAgQ
6vwIWKR7MuntNnF+A7Ejffs4Z6aJuaQXL0prKoTj/FkSh4LuQM2FIji/Nh0970mXJ6HLDfkKS1f1
WiICfcEwdQMQ/ogK0ft48GZrOIg+7aU1B31Dvp1XE5vo1viUjfoD7NuikAsDU+T7SwcOjkEpPGUU
5wOKs+wJQQmI5DARJKV3zv88cnaMfchsyArocknxnxaHbi0Hs2xhe3uMkhKc4TsM3JxazyDn6GPB
2QZBpHJ0lD3LN3Tb71LaTX5AlFxAPvHiMXIGWHu0dLLm3zY2zpDuMYL2U3Qb+cB21xbN4ZpT4mus
56fZ9HdKl7nEdV0wi9lPwOBbDMZAvOoR8qLqALmUxlQB83JbR4qTy1VYknckvji1uksbSl3slJnZ
z3Uaw8Dg1VNuIR5d44lqaLn9rUer0aJmJsUeNH3Zzx01aRDiwRwU08n0/6QiLveQs+UvMqyqv5T3
TXErngzQGFjZhM225VwCc6Hn8Th6g7iDp+JxgejmYb4Hkcx5sqhDJCEirDsQpK+R45lF6GRG6BSs
EaeoD1Z2GrB9fqoWcePSVtes0hNYYFOmLiACenIdZ8wf5vxEz1zR3OKAUmXcjbHwPoDOgdxojTFi
6Eu7mts0ZAMqF5UTc/tFZdnhrqvsuOC6kuxlqdkDkOqs1puD0r9K96967ZEVpg4qJRSbnIuhOhSM
qTPnBlmFH6eb1cy2p9kNjGqL/jTjrXzgPbGMKu++URP+4lmEnS/rLxfTUUF3fEBu+CGoyegGNLOI
IfuQJE+f+E1bxq6gGEe4aLuOjeDDRTaGKWPMR9ReVjt7Om9Xm0+sT7tJhGJtB/BuVFzzplm6x5yL
Wzc6Kb7UiNC+uEHJUq1Xs3FGDV3cA7bIjw+P8lKe2327uRL5OODADZeyGwN58KzqLX3AxeiUb4Pa
7LfTRn9W8SMWCZcv/bn5wm0Ufd7XRc6C6sFCwwaE/4am9+mezYdZFJKt0emGdbGERGig2yxW12MQ
fL6w7E8KBpbqLRr4gTS6Ggx4kpXHp6mPMNrS9ePCwRkK3nfwZxCE+kkvAYEhi8OeVc4DLKG5YmQ2
aDRNo3FVlgja0sBYL6Z7htxNU/LomY4OByH2gwAkNIw4cA0NgFHAm8sQsFBkQb4b6GfikJrlspdJ
+RtyLGtL7ldMjePZNgBRgkyiHGNrIXsS/e0TZEOaUpbO/KWYcGYwBKUK4YtC+Jm2fsxAVhib8QZA
R5bxgDeBQ4jJKtMdnnswgTkydKRzuvrq5kNkpz+NDOePmiYW6O63CEeem27blt16IY8Uv553BHGb
LXPOk6MFR8W73oTRILkgAaRjnhnsk20tB1GN4NPpIDmvtPXJK7aCwtXU7UNxj9Vbeu52cdqBVdfG
YFf3JaT/dywsIhjqqfoK41MgOZjo/gSCZ9KTqykNPBXpRfu77c79L2dSXdzAtFcUdjZYqnTSQtD1
kCUBWamBnkicGWJCFpD2Qe26nq4NXCKsDpSqOBHaSxt8/Hg1RcZyGl7eGTthruPeJH0rld+YFFGt
1OBkiRaHTWbSCWFzypK5oBWaUWpNKIg3Q2WuX/ARDrx22unk1dC2cKonZPazWSuhnHUu9qE0U7wA
L9UKKmTVF1y9AGZQ1xEE0mLyahSSIFkru5sUYjVGoQN3zKxThEHY+uVsgPB4ONAaNPRgppmIUYpC
aCOY0iGgkduogluPYRHGc0ruahbp+B9Z6e4ibyqZaqSJhnqWUdyNxiIwF0gAsMk2zDHMjh63yGMT
IHyFxD4kKK0Cxxr4JzvlwglStu3hWSZnjc8qHDGnczJ5G8zfhq4pLVgppeZPfqxBf/6tzfRGPQJ3
xIB9nffClC/uU4sGRJAbOxjWV7NZXvD6LXm5GpyFy0CURHWCpNZLoxgViXxLZDptsJhfd/90DT2k
citljD3A+o/MlEysGLv+UazTkMmMV8XamRYz0A0xoISa/YMe2YjJRFRdJkJji6Gwasbr+Ilzo9np
BijpA0a8Y6GSErd683lbzc4cPj8pokt6cqtGo7bUs6J6U89+o8bRHKVCGicABQ/s8/yamhOTi59D
LsA0AOaXQNaobc698FvS0FSxH8wy7idR8+ifuNwUrKiLz/qKtF45GUK4dKn12Da0TDw9YZKkZjSN
0JGulmFgozVhtYWYhZV9azfgNHRJ5dku2fX6SguPhzB8a8GlU9vufVMSRnc8JRF/S9jo3iEvjxLJ
mUC81OhTplR3MQSm+ZROGvi/AazAEefPyF7wLdS9X8gfDgCdX8hvqD0WxgRM6mGlPf6mtEYoCSuX
G0hDera5DwBICPg2K1264RuBY7Mgw/XW/9urf6ZUatLw8NAQ4JFhHM/3IkZDWL+/8HqieQnHsNyc
1Ue8wsDFh5cGGMI3n4pdBSHpIjj6DFwhUB2SHXY0JlSeX7LD8Gk2X4PlTlZQUHDl0Y4zyimsF9pa
LzNQui07VwG7uw5flotzjHWeHu3A0FRfKo5NMQiH1E6qJkkGOtyFXsXpwr3ilbL41gOsm0zmHNYl
shXXMKgbGjX9GLxt0bk0z8Ef4psQM3+5tcFTkfZuhzahFqxMCAVfdGyl9hcQhUVMaB+oVzAfOBeV
pkmN9f9c3J8SNKQHkg4Q/ptYWggNlESF7/JIH/0rhYBaS1116Epi8h3VKi0p7ylfIdZzkwfdXXNJ
Wo+bwdjwl8CuuM5jq2ICGa3y8MM32cM8hyNk33d4evWs0HtmMUAE6qMS0SUdqcbBP2mI1eJQL1XY
vYtvd1TPwq4I6XYn1VR7A9+kwPt65Qp8XXAvn1sHkfQKRiCCzu7RSDDkT6JIKLe2gEx2+DUfJ7Ms
JrqL/cq6vbPImCm5ONQBvFQq+nDajVwSnJ0DtqJwjaPWEYQet/lHM38J5HIgkKmP3Y+mB+JcVt0n
X1B07kpLeEpxg+Ba5PzZOnaYuAtQ+4EihUaEmIfWGSALea9qT7dY2axPnbBMH2Pn5B6iglrZUsLL
yczH66MQ3e14VyNzRwuGOslsQbJpITGrY0+y5p6K+LNrfRwMyOHmMcew+M4RDl4TS2M1cJCyOHMx
DXkzy9WHu4fVQtuIwjZm3HyqwS0kxg29sDkYh9z9+dP1W7EZ4Tom1wpI6RVimAXf1mP71c1TTooa
rXGFJjaufM2Xy9+eQqMnijqvWmy7A3AsOEL6owXv1PT+liGphycV51YyF25fkbGy56U46ct8yrqk
ywq8dsEsdLy+kPZNe2HIOtfFvnmyUu5x4SSWnm1vvy9HuC2GDvPevqQgiB3YOzIDiGrZn4FS2Q77
HtlmToWk+qlufUVwCdKJC3K3CKpOrRGi1FNHq8qloJ4ChXue9RCmtHVi9WNpEj4yueslxumCLvHW
oL+v8pBbWWARAz0yu2YpD0UeG6VSkHUUITzA5bDUoq59yo/+ErhS3+GWs4QH7usQdF+isPeRnuDz
lWPrl7slIjwIJfGE4KTOtL+MrrzgUoEBp4ZpGFAMkC+o3APQDLGDB7ZpOE0t0onvI2lZ2FIbsjnx
1XrlDXI0F88GmlPQGPzkPdNQ4O7riqeInzFLKA/POULMFvNyNX+uinq/wabptUAGtutgEOd3ny9O
DBJyN+FgMbrIga+k78lfZtJiA72K1shesIVcNyF/XN1Xx+HxnF9pckEiBsbWLq7JjBR+8GVzs1d/
xPV+S7p9nh7YmrFXNTXYCkr/8v4TcXnWE0OHzgj3yDT6HPioobHgg6Vgg4LhWwKPR/EJwL/0ljDO
67vmwt1Om3hQOC4aEOQenKrCn0kgrOjaPDw4pjJPLf1u/CZTlvfnM6t+80oD4/GovzngtVzE9X/a
ANfuf786gI5TFBZ1p+X5cFs7HCeWH/SAmb9KoZdrhJ972ehj17esgIjqZ8vW8li9AwuwcS9YM3yk
01J6Y3upo01EOxP18Ea+Lp+wQwE/FD4D0g8MdL2PbvBht5FArVkGWHhJoZopwCJB9crOY4GdvKdo
ENhuX2HTePGEk2x+5ESuC804qeqXKHHL+yW807FPt7P9BNFLcLChShoGB80wak4sEeBjBPAwSZyt
OEZL6xkp82hVWO4RwngMPAbt1S0egXlG7NtR3yOoXXRIMpYBjNQnPbU+7wBwabtzR14tf+QTRrSQ
AbV0k9ip2jOt52yDShp/EzAnfAzF6t7/MnUtZbByk665VtG3F8gHHn4xAUcZOfSpv4SO6ehdZcKb
c5OXDpKFoJdNcM45K7+38BY2Jk8m3NXnL4TLd4Xs9hLWe8rnSgVoeAsPaSmIizgMIDMorqjUB/8U
CLDJthePOp4Cq4M7ituoUEYj7+ef3QHJwYi6GtQqu0kHStpfddG77c4KOgjwcZPoWpTJknPb9JhR
WDm8UoD8EAOiFPPP26OrfGpUYFI57EAj9ZVKaCsmDETXYFb8krMUQG8Fa7GG4OuGDrFlkFMy05It
5WPpGTt7/qG5taV6WuouwaShMa4DSXI1pjJe0h6bN8luGnRPQ4iGyRsYQ5FMQsCpbhSf7vLzd5h2
gzJX039j1B8gwRl7i+A3L9M1Jqks3ipbCoxuaUntlW3IjQuqLtLc7FqAVS34qUC7WMU+DmQdZuLy
9yjEs5uPJeaFHLzo/9CMNH80izIyYTpm0hwUv4cQIQKlmKJdTeYeGS01yFN2+cRCKCtPlBJxbqey
1cYa43r37+svD2JTOOwsQYOLJSkpERoq7RrrCRDqT4JknDReN/75e5mYsNzwZVoG7JxespdhOpHt
Ek8jz7aq7sDdUDJEnlAYe8rV2C/oW85TEzftDe+yoSqct971C7wwn1Sghzoy2GlUoUdRVNq5ChA/
6LczaqNMRXqwhG3dmKDwS+Il7M9SxxvCrNQw8vJwrjGIcg7lu/teiH7x2PsntYH3Ju09pv3KDMA/
1QkISatmK9uVDF4g3bp/du3SvsgV93q+luJhz99vA8O2kk2zaeM9ibGEL4U7TjeSMFDtgrzBp+Wz
x3s7uSBm1X5/aZvs2Ivow98sMpHJFoyhCo1yaBtHGkqmy2p6dpuwITpCxd3jpp0rDngf2ii6v/D+
nG/eZJrSjSS1COT+E/ijqXh5dcwWi71oukb2wG1K6Qi20UcIt4BrccgELGx1ETSPAYhF3kM8X7i9
SrAeicui4OHqvUfRLnDlQfNQSv6R6Rm+ru7YP3IQIt1u4esL2ySP6eXNs4lZR31v1AYeExUfOPA2
YzzSWO/VvgDAVr+57+Trbam9n8KhLd39wu5nDkF73CZd4MD6GmJ08jfz6SoqwfcIiP0jZ28Dpm11
ZljB9YmnU5RFVRtOiR0mYImq711TqyYQkc2gqtMNROEsBSmI4XXtgrQre7siy1dMD3mAZ8qU9gcr
bdjFvGT+Dz8FGKmrQTivW/0/jt1jgKg5wQK+2hpkMIe5Je/MJ0cUuYFepInMJHeH7+6Gk3zMAj4F
LPk+VBJzwhh7LKKz20Tb9gcRuSpUZfIRAkp67enf/biRLcALeTTREq9xyQ4i9TYzoU+74noP6Jxf
oEiUcJNaDVF+Hv7XKVPMF8IRppUXmECMbYPDHjz7CW4uOjqVwYVsQVf6RsVB3L7Dh7FvTPS/zzS1
oQKxperOMfPiSP/t71PNKBfyEDlO5ohwteao2TDkg7OWlbNT4kWhBUgXcgAqZk6B1s9Cgj1xp6vB
p2biVzthe+Gu7p/MmL/VpaDn+5KnFCH0SR8NN8qdMyJy+pJdoVGcGvzgArbwLhmwQSDJzT85xyTL
js2RiNhqLGjU6vGYnP901Ud23margjfSNwi5lXJiyTDrIF0Q2JFRdnWsWtsXAq/o02zUxus8rZ0N
zl3TmWxs71JQbm6KCj0HiS3kLvGVJQY3d0jMurLj1XIcd2zY30NDHKg5RfVZVX+KSTuatls1ElZC
BlvjV+eNY3xESNonesRKVXCYgE0auW3p6qVmwuVnehfGk2b4wUiNUSaUdYqZ47X96LMHVGLogBQJ
wTDF61B80vtBBfDCAXyacMe2FC5cRMa6lH6jMVhUEE4kcBlC5tlLogUdVCsjidfpLfcwNnbmxxow
lBneipB1gOzfa7dFuwKH0nMR1QYqeX4uxm9Hg3AolGlZ+XDfUEWr1CfjeAbzoh6/sMTdo+Y7mQiD
0saUuaGf2ZygN8VaHN9HE88V2mZsGX+S7MwJFutvZj4A5+skGqZ3LZNGc8pe/amgH8nbjREzwtbh
YlS2ZGF6kXYqB4sQV95AynRUhCg/TC2+MNwMVdm5C1tQDjfrCVPn1OfokxNIUg1za66OF+al2uNu
GKrqIT0kye7kxUrCspRlXeYF5DImb1sVkFzR+MNvW9hn+UpLUxzQEow9m64YrMVG7LxtuG3zejsU
I0HRf+VShsu/AojRKGngo7LtBz9M0lu/t0M6ZlSqmz++MuT4Y2qEkBCoRGB86wX+nkRbVSdRPI8Z
57Deuj+HXQlqSb9tUBcGsPJ1u6paeTS/+6wtR7SnQhHtvziOj5g3rSR/05IYeiFLyxb4UkK9ADNc
+/uB/g0K5ftWUZ9ui1KOZkBwTU+kA9obUdEumgbQZS7e57kNCwnb67y97DwLwcEkZMj7VwjPGjTb
nbHIsJdi1ZLHsGK3AN009DVZtCj4QdnWCvAmB51zy6J93ZhATGCfohdKu8WDLNJGm5AYdnTUU+lY
7gg2gKp0HftHSohHaPZMMX4vkEx22HV+MYD83A7F9mnc3ajAkE82mUrVbp4PU69YvJVZa94DV7Eg
G4cFhLbRX7DYYh8e+h4O4idwIPNcPELsoF3CpdbB764GYOVRAEBI/dPSfGwLafktEXgIpJV9ZkRe
Rcwt9GQjTAzySZecQn54JfBQj0n7b6MxloeFB8+6jNnGk/323n98YF5XUio6rB8ioAiW9oQJ105x
niW+mrcRBnVavYVv4W8dvzhQr9i4lUG1teqGNn+h7eJBEd0/fYCzzfnho3vYGp/4NttV/aJAneOF
VjFy+EwSui8x290euFWI+5TEAvZbr5WVfAtx2H+2ri8j02oqmrK1BCAo8b+gIhPuDxUx+fi+bbC+
+yjJcbh6Z/6UbVZ1Rwi47aX674+eAlzljy4LBohcaDBlejLO+PhQUF2P16r6il5BYTP6UigssSaz
Qr5AyUImNF+SnR4NCVCo2VChnOcB5WFEJ3U1xXaZYT7KbzxrUy9vgUO9MMGZG/7SOesBvSSSZT9t
EUU3WgWOs0ijRgourn1SoSlQ3p5u4SqCHH/rJzPULGrG6ko8AAsLEFf9SIkHK75Ggtr9GqU6096z
c85FJvMBH0RMvEDuzes8glAMpZJhykYCOTTZ4EuUUg6aYDd0i0PQWObOOAlj4dYNjnI9Bmzk3bxo
JtDkt1FMFgFVLKSsiQZeEZDTWI0EEkr+3DxB8Gu9RYpRD1fIP6oeVMmzjfmaizJlxPeiU71owSei
L4E25JUk99cuGznt3KexsyqXBnnGetd+VyFrgf4ccE5MsSU9QJNH/+66uZ2LhiDlxRbSZJtrGFgg
wKG6c0AJyy3Iyj6v8j7SjrNiVeKmGFRgkuJlejAKjFhJbko6goA/0I+Dxyqj7fnuMwcxSIlgPlRg
XKpfNu9kUeEa/vTclUim8yhDGT6syiyMIQCt4x6fJdC3ppIpeJWpFntfEQSoIaakg9MLCfzVA3s/
dPmPXso7mneEeVZaqKAYxoEz6a2h3FmjX2dt+lDv5V5XHEFlSgo/j86VtPgxUyc493v0oNFlYynh
UOH0QBRMdC+Y2dvYHALYI3PEQRnsowYAeJUf22SDBQq4k02OF6znZblMBMW+fjYJ6lkbjV/tT1XE
0HrIg6xSrKKGOUMUbpyp1s5+LQSuh5msZlkboJhiFKFjvYfhN6ct+MQdiiHXwn6/nen+dYwuzN9x
BJV9YT0IQVLp2eZgrewqzIFQIVKsa2TM4Y7XKCylvq3sjUTp90Bq8Dh+IPqQKueYIVmnSY9Q0S+o
J6gbjyNoJWrCxI5sOlLTBIrlFrviJF/5/mnFMbRc/psTkkspPL+UcYtCXPk8jyMht5aUVSSGNxmm
jw399CJg9LSJWB1yEwbCNn3pOmW2pavn0s3nqUJBsMPKrDuRpLfDKbbhWHWCqmk+RMPgBp5kKaYI
WWXY42tiOEkb+AAXgJQb4N5ts/Y5iGLLTW1gpdQHkaj+6BHjO4cKrMTgwaQPAreb0QGEW8HwbNNB
jMqY8kmEAeHUEvBRTyuAmKAlpX+RDNv1d5eFVH5Kk25iMo1oUxy/AI/Yt0Xpi1lMCdFZgmiyRPsq
1DnGi1gws5YBAxpya4pUKsudKBhQOCQ5OoiTo24o0btWUXWQwbN6SZVNBdkMT8QvEkTEQ73SYFXX
JuKIZFZ5S72dr0taRaPgKS4y192xPpY1jMipZFRoPMfN1faKnuslQq4g7c7gDY7dcDJ1yEeLR/eZ
H2mON5BtV7NlMkreQn1Ke0UVNglHjkP9xad7CLmdTZ0ooSbeip/vrbS+7FE6WwdBlEblf8vt45+1
niRibVALnKyO81mPDeoJfiZcGPvE2yq1RxQ24BZxHOyC79ulUbwTfFMizp2rDHOBAse9fkV8n/T8
rSSCVhin67tzUIkWCqnmu/wuBzIyVOV2u2HZy1ucs1vbE1i38P5QM6lVsuAUmwR+sgbXB0E2UvCO
SNtql/XyE1UEE/g1spnIZ51t+cozB1L/9DROYvT3gnbohIqAjvvDnG5BQi/hTAcHZY+DMSKwZdLu
o4ZF5IpwRM4bXErG6LY6Q9yNKJY6Vz9oAdkArJlgF6hRZDwImKiddGsXVVXUiQ8OQVVt/gBWkemy
gVI0SxXG4rNZNGwHlFalW6iD8LUQlT83qrAZThvL1jNVIjtbpc91Ay9QMJIAqbXsq8FtElr2SSUO
/P8uLwkqIvXbEQ7+WPku51geKY0Q9jD00h01AtizR8TrDC+33ify27niBGYTvx9o4KNM6pwaS3FU
ANOGdzuzMXWvq/uuY93XQv70yJvXAU7nwjj4SYRZJBbSy1ZfPsi+aK+fFLYUN9FsKyhQ0lBbfkH2
SpfayQmw6IUmboTFmDmS0siCyGUS5BaydBCeEBwAhIWcKsHipIFwDSy5xAXKf+HdiQGYdzkcstpz
iYYQ3uYUcn/LFLuxVEEYCyvLk7wF3jIiY97PCq+heUVTxZ2Fz+AzJIlKeDYNDdfbBea2NTe0wLaN
kzFSB4RJda4pGxqJgungewbNEp1RTaL40fDYRKUbcu+VX8z3YAu6HtHliMK9vulEBpwuofY+uZKp
U/T/yYJcDKy2qBaZpPBFAXMGLoZC+f5ksoIomB6oAb2GI0dhnJphxO2Frwpa/taoTIYy8jGqrnEn
m5FWDAhDbdfmTRPtzjGmhJ0g41syqWnUogDdXpAgcKQJRZ6IfiYZHk6L58nqGpJ+07W00zE9pZv9
39MLG3BrgifgaGT/MJh9QW9ua6FpsELjEVBKopJ2A/nlIOkKmKlwrJpvJAs7RAP1YqMWZmaDWgsd
v+ED6UMJbrWZOD+M4eA08hOp0NGxC4jdBDuA1AxumLtcx46F2aQP4i4DUtVOp7VQHwzGKjd75umf
yXRqxXEBODz+97C1b39J5pyD7S4gAr3jt49+PZ2sqC7EZv+W0GpbUD+jPpj1WhD7JqMaRBYy+l3k
EkH9Omd9th8P2KajCVsSlEIs3hlzUZ68MG7553ifkM0VS8XD2oY8DAoc6ZD1CQT3tBsG69EVZfom
IXWmEGzamXkc3D6ThH1IJougKOuww8v9bepJFUmmz6oRPVq/7XXSPnGB2mwri1+B5zokT/ZQM6sd
WxrXnO9AZsdrmkn0rvPQQdixog6QqUTtE5Rq5AF2Li4ZTk+M+3PLQbbE58gglzDln3U5InMzY6LQ
m0wU+vHRecC6WN9osgyDCKAS5qcrKJJnwXxRtEiXII2wTyhR8eejBUN5vaA/Za2d8cLFQ4pRD7CH
GpwgKyH3HE5SxU+nWaPN7jAPxYdmz6JMBfIfE1OgFopDEdDZkEE4VjlPuit9FbCUSatboEcrBbeD
G+uvx7CqDDcb85AQCHiJ9n790wENHyoeOUE6Md1z7xZpQDAgoHbhPVEHt8lHyjDcw9TFMo26iZbP
4MxFVoLbNGgVaxn0akMvZjemZEUPGSTtm1hKEd5u6XYTJz6N9bKPIJeUBNN2vJrjBskYA/U32n1v
qgq1kv+foz6GqLRG1GojswWIOX5wioT8aQzqb8kYp1dvey1BvwfsQArse6IDpjYt0ejVpRw1BVrN
5RsMGnZOKdhHQco+OjYn1wNx2TJcAg6QqN0uQguWDtjsFawI41G+yOj9DKtC1EH/cHWQ7gv3T13S
KenKJqwLwTSQIxy6tKnJ2XD1m/RFKD0fx4afpxsgXucmJznpBlAOYQymGWfZQqOpghh6VFCGmOjq
3JfkBlbwm7kzdF4r/tle6XR42gogbwx+1uQrq9lXdiJxb8M3e16s21jPmGB1++Ny69Pz7JXUQEkX
nFyD8bFba11eZMppUw3Wc3w6OJS3jdmJHK0cEQF0eSpL9v5QWzKXyDYqR3aWvCdVpea0r8oRpmjX
01Wp7BvobQCbGYbhAA+g5qwpgdiwC0HOx9+sB+na0yfBIiAu8eJNzwryRFWkIDGkk4xzwy5zsowZ
6Vwvp+DYA1GzIb9rXwUOFiHgmj+N9F7WYsXNGlS5FCP/6Ol9kifXXLjhi0ksG07fbPz2D2ooXFW5
EeEWb0sdls68HCTTcLLKv5qEvjwpeR1q4sYJMtcmNXxkkkmA7kw0Ds6xCar/g+uJTQ3EuGlPgMjK
tM3uLLuBsDaf4t3SZIJmXd6DXQKPrTYbcfIm3RHA2u9jPFMXDrX/lUj7rJc5J6SR+Cn2CH3f+KBZ
jghAjtxY49OW29pw3DWCi6sebvvXzNqLqx7rCX7LetsEc3QMw9ft+vdVr6VSdklGJ2FQbG4RTurA
Tm3iyU5498bDE+HXhREVJxUVOv0JZ2VoG4Y6svg8HPGNmpctWUu7XrX2SbTv3me2fk8AVVBWwGGd
1xm/lgLu1iIsGnzpC5T0g5qcSkZUM86qM91DE8y9F6dpHZOxzyM5Zc0eXtO1izWJP39dYua36qFt
2DOLZNbXRQfnyIxo/gqzMoE/Ww81B7Kfo3goeDe+KkUZN6y0AZXwKn911rO/alBfsd1JheklI5iy
NRliswrmkg3YP7ZwF/s8gHj+muoZpKoYwLciIdPFu/R0FB1SHWYWfgg3ihB0od6P/UWN16m7lkUC
z3aPTc70qs2jbUg1h5hH5Cw3R5rj7z3RYGxPVX7iRlrC2cB13XZiHXvL163hawGrfsG7XLeWevtn
AhxbrWs4scywk7UeCfJIzLwVUuYScpvY4k5r8sYHm9XM+rTbNpbqigjP+b4QTOGqLs5bqtWQ1yh6
mAOZ5xp0UfMj24wNg5hRv+4vgRQbS+3xvTALo8aF/ii4rVMm5MuY7r+1LwCzP/abJGNUST5CYM4m
zdSU42jfSlgwPHLCW1YMz0GUx0ZMOVJVU2wxWhuqzYjton5bPCrK3CxE27/L0qoWHJOIycMuPfZj
J+AyUWFEvQG+qUqLpAsBLsQ6suNDU21MEHlYb9+HLQVpXZjuDu+zk+WospnBCCm9k5bU+A6UONwG
L8Zg/+hC/hWSD/khoBHOlZTO31Bwvjjl7a+gkV0D6d1a3BP4kQ5M613nZrDuvCwRJJalFYJJX098
2it0H5eKD1fXz54TfT7+uMq2tlOQlvAuUVeXrN2sEoPiXRL92EqGWeCQSle34GPO70umhfxzlzIL
+ph4AYQJF3yT2Y9sb31zZywm/HPUqWa3f3Xdm0KaIrMC1Zdy0CsX3PuiFEiCW1cRV76indDlYT8M
NqRI4QXozUOW8Gql5hfqb77yvnk0+Imr/LxzTDcES9N6yNxsuMstOlCM5Gbe2plg6vGP0quClAx3
asNXdf+YFfv/eS1YEaRwbuKtp0B7oaKMurfX71y3R6r9losa4mGt4VWfraZ/jd6T6heqjx23IZSn
npDc3MmuX02GDm9LAupbVAjz4WrwP+CXOVf3HF+l1gCbLlfHmb/r+hhxI8pyuLN+P2sYq6QKUdgn
RHM9tTDTa+x+ho+NOzMn+reVWb9ZFYUrrvdNxM8M6TzClb8EgdDbm1wpIcU1fvwbko0T3Q0cAcSF
oeWZil9X8WtpehP/n4nzIKssrajvjnoKyXnXR0iYou9QWfQ2B1VJNA8DivjyxYeSFZBpK/UraQkY
vFU/M575c2wYFI+tmvyJwmMhMvghtsz3/u8UF20tKjrOxlfvRYjUvsQtG6GSbUDI2a/QUyX1kKIM
xdI4dWiKKXrLTEV0KJIxgeUKnBiWpZKqJLWOPnke0DyWiK3/Zm03nd1bThs6jw4IqeUoM2RKVhfm
4I+/yW8+bKgYs79N+AXSwqoR4Wp3ObGjdQTBjxFJiFyemhBBPcqVc4T67/C/9jkfd+LnqaOPeGCR
ltBc/FxK0Ts5hWarUUoKS32sOxJxC5noJWvt4vmv+/E1uJF9TUVf63JZvpDx2iPbX0kOmNxtB0RJ
W3oEqlki0RypirfUST0lQAWMnULKHkdnBCwTKGn3FgjGnaX8PxBGB65pj/85+SWvoQn1nzD881rW
caFK8s4c4HZ/cuzpgqFcyTk+J0brgobUK5Mi7SSqNxUpKpLat6vHQ11U3bW7MP0PJxslBt5xd+gu
iJSZmEGvT7DJKufsl25sL3Fy47cBnu5zw7njfLoKddKNLlWl/wcaja4Qy8NscV+BU12aFo3gztMB
UqmFbVUZIRn7+2noi1fHMJXJs0vS9NGZ6hMT7MjD7RfKz/C9scQvDPaQDw9siwIEr+8oJzFZxIIU
UeNGdZV8bnZHu8d8LVAYvyv41aC4w18WaHFPgZC5sQnsbzBS9i9rh0q4JdmdSyRQLFkr8+Dqmu1i
//j/DknAxPEjTDAok8YtTNeTkHZ+hYnK7VYKCOtLXdAODbfVXyya3AVGk2z7I51z+JsQog2Xy0Lt
9S1NZ9T2eD27fXsQ92LkPgOj4Rd09WbLjRmel6NAtRBO8PwVSJa0KGjj82oSSJcu6RJy6QofOF9j
gp0b/wD+/dWrQsTzER9IPknf0qR7F6dLJie8JPvVd7ZQRvcvHYFsZ1Hyal6GEkzxM7TIJia/bA2h
8m6Oa7LDrguaRA8/wk1T7GPvRmoHFWy3R2N+uhoD6M8Qdp4CTOnnVBTHtO+xk5jKvl/iA2o/Hk5J
335L0Nu6ruREW0pgiZvGmu7atpdl0X464bONNRhfRk7PGOVa6UJEmWMRPEOF8vBgtzHkMFwUUZ9A
l/Wvdp/6uncbPJ3N6a+00CuVzojY7ZC1ydfmQK/2LjClseX7D+yeGS3G0rofcVmMNL0zwflrR0VT
oSuh6zMr1BWYNZkeEJ6YGSQsXngYJkCmD3RzsWk65kyk5N6G88B9dovNcBkVenqHYsKFBHf7fthq
CBb3NJ1cg6nBFAgauLu0ZTAS8wVvy4EMXwHWBMR+0gTTHkGDoAuE/NPTm0a6KzWov79mXLD2G03l
xyw14bUvLZBx7SGePMxUB9y6S3T4AyWezujXVgBTlSneLKRWKdpcsWaLwPywqmb2kA2P3NIaYRdn
0r0865MpXtSpK2ffxlQT262baUt0Dc+i7tNRSOWXi6JpbihRoodnWRxzCp1hgnCzm0LO02+f1MoN
9GYyBuQ5enhFAoS1s8flnC5HFU+RPh7jNsaGPQGK8Hl6r1CiksdaKrLPpZZ/5qkr4QUhCQBIah72
Yr40rFYi+gJmtvwuutx2XWQUoK4fR986pKpAKIIh9CfV7pokUrtY0I7bmNrfH9RbvWY3QLnwzTGm
/4m2zrhFsshwP6eVsJqdBdUD27TekgEb2Sqb9HiG9qEVvb3aMsvY5hZBjWKOBwOOH8yDqj3TaS6/
kwC70NlT0HATNlNRxU2SrMRFYth5NbLmkwPvnnhhJozsLJVJfwxl3MPBCTyTkxYn3rb4OrzzG7JP
IJzhx+/3B+W//NSokiz2PCLoj/JCcEJrgPNt0OVSCYSXrCWAMJJq1BFTf71Te9agJfk8MAMQHc6D
wgL+Q8PmbFXGdCE+Wa8d2yTwn89G91kbiR1XT6nxdWvrODKEjsasPPQf2usy86a/ZH88iWLJWQAc
yKLNBg/oFlzOi4dPAqD+V88fJ7xtTOml59N9BW6TKK16VNN7QllhZNQWDfE6KlZJzBd/jmONUPrb
Vnn4RqbN8A6/xqP8rrRw4RfVW/UwRN/Yh8TY3iVUQyH8Hze4TbCkqLtcFXRzJjxxmFiQxRks2g43
v+DuVjoKx6C+qbFKVZwY/vfe4cikssLN+ngfx7XTN9HO6krSqTxgG/JD0NEftKUJyANg7vSAqa9X
B5qlJDSjhkHLYjx8Jb4DGfos+1CH+lZqS+MVznuli1DEbEqKicYP3vmGX3ZL1xV2RyvgPeYgxXmk
FNEwuVUYj68OkZ/ZqdIe3Mnr+/PehvkZAGSK1RSJ2Dsx2e7vveJK71Jt235XzmabDWDNNlrTi5+n
KNYCAr9tubb/3H+ZrKVWJ+9ic3Oiqag5KPJRc/KQYqW8I83b7qc+j6MnXnwUpFzhauDhplvMasU9
DVHcYL2+Os+B7u4vQxPgrNxwy3uQ5BeHizyz8c7cDYkcK4mnry+zAO/9cTosg58u2aqXRYKGgQSn
osEmqPpjFDPoyWTb6chowBe8UPEOy7LsWqY6CH40LFOTlDsJxfWrzOd4cA2YGEqm03TjBBiIBfOv
Y+MmsPE2+IZYqOHGK34m0etvVjaonQpMDPLU06Ln/8D//Y3HEjDhPI3xN/iIiB/vezHTySCvqvfv
kV8gp+PUPowS+Cw6AtOlvcNWQ2A82yaMypk5k1oS4wFGF5xty40y1uoWbW3cg7hWqcSGQPe+wis3
ogUkMX5qdiztQbJAMqSLPfrZm7EYy1xTJ3O0X86uhl7n58Qpf1/nq55HtescT3vQ+0hrVsNvKE8K
GUOZNeaXrEfuUvBklqa0C1I8vTcsrHQGqtSAfO+SDdzT7cr2n+Q23B50IsiR7rYpZNlDx/a021x4
lgBqn4h0QwoCrY/CbzhujdrvAxm/Vw6Mtu6v+AqmclMc9UwmfUiRdEmoYA55qL0X8DJYldtGRPkJ
JWN7rgsOmnvICvQo2JfO8dtlg4TzvYqDvhIHWyjMIJAhkv9RdbZYvl8OUuRFpcanzWuy7LGabTey
IvfBiFDEFpwmEFqzZrOWOJB2SDY5CJKZQffM6Rp2xxSETWPxY9FnjeMBjoB+X+VKQwDVOHN5cFZf
z0R6/cQKQ1t5/oNHJnnOVCIwhPucJHQOy4QkPdQ3yZZdKDaYPuKUTVTdk5PGip9dAT/s0LzwnJ4H
sBW8YznogoqAbMIokyRjeHWSdBM7iUU09mHnAFeO7HHDRygIFB+IzLJWhYk7gfFvHBNu8I20gabg
K3gXMXZ/8QP8s0QABWqTQ+P2VNZpuZo5jTx4Gxh5ul7pxSxn4vLizRU/TsT/aRXh+blpd0N2lY/i
86kbz4H2GVMNpXpx/ZCo6KkHOkbPwZTCaQTj3GmR01AAbmoRP86ifrCUXBp03brD2RqedT3K9/kb
HnCC2FOad8XrXj78Fi7YoFqqZ3Mi8fHHakPL9pBzg0wJO2RDDmOVu8IV57ywC18GqRaZYm1BjUG6
+eF0RzS1O0KTSAkkjO+MkmINM55rJQ0otOHe3hddzW/8w0i1vxCGzJrY+2coQr+PF6hyUHnxQyC5
Ozy6r9EInoqxp0Fxpe7y4ISmAK7Y6e+L35n/h3iYBRPvapUO5GzWEq8WL1geZZx+oBOhnJ0zw8Va
KJ4s3BCe0tahavkFIzDifJAkLY/vlBbNuU4TEvRTRPkP0QGblWhOJtpBk8b2ys3blqJ10hVwH5yy
V9Bx6lM5kedtOI+uQ+AcRKXcibYsApV2TjF/cVkOo42uphn96WnnoKeD5rNlp3031bkcOpZU3W29
GSbfqLf1k0gzoJqKJLhXaAAMYWvdcKEFePtCzkG4s0V3SwsrT2nldt4gPvRYcRbaKS2wsAchoAYd
Q4+F55vZmYBkZGWsPfyTUJtscDyGDrI7ZoSgJ7K0xs5ImU27yDH+GZ+kfcese8dthvIbAPJ20LMz
6hShdjORNcYjnznZ7t1CZJ9jSRPfw/MtNjmp+GLgsTeeRXTte+09uVj4McIfO+dTYb55wuz0i2ky
M3cMcKv1am//gEf+FutPR3bnjTKaj1ftoPuIsOKAODsajMHjg11P0b66rAnF1KefwL5dscrFy2us
709pVHIIZw0cSHARVgNVx+t63WdzbWbCi87wEasta1tSEP+lPQVBcbBDWKuAjweH5c0wpRj0MYsL
Xa7NzgMd56MoI4y8j5lgR+Qb40Pxek43E4SQU/9Pp7uB80V3+IobO+ciJAyaAfmDWckz2r/JMWkC
3Jntv6RpeYNZdHpq3tOdcTEg4mRG0adzNl95C3QVtl6Lddl7J7GWs8WpKiEGELm/ePNa+kwy5JM0
z8ErKCcs1cYDHDfB5ymb8wxqx0Wa62t+MQwsqlIqC0es1cnOivNmYw784DIyC1LB8zbLbghk/yGh
TlQ7PhOMrsa+isVLB7F7OArzput7Ri4zgzTaau0YiuYWCiPgkN6iqd5y9otUje0fVoavNW1e8/st
ylhwZUMex2YR7iHdxFwpVkzNwfR2wJNK+C5UvBBzWoySA1/LDue54vObheiRfA1QnohGZKvUlcrp
R2twRPXK0gJK7NAaT1uu2Sf6+ic05dyIGEpq7nJ/Nsxt4gus2OKm3B7AkBUB3yZ40wG/PGMUbb26
c0roYfpjTZ4E1VDjMJs0qyF8b/jxH6nBvf+3G5Y/YlrAA1dhTtENfWZzw2hrovq0zX3aZPf5RZDo
LtDIScIAbzV4Wr53eXDAewhPoPFjHewfEJBKCvF5Il0Ocf++5H5GYngXHeWX5eQ3PbebVnpHWYVa
nbyuvvroBTzEKOw6mpXP/tJ6Na3+gGAd/DMVd1EmwODeC92XhRsGnK52rvLgd21pEI+yvZFyQuxJ
11XQMRmFClcNp77lrSmqqEaMr2JlQkeJEghI0mcRCSpMgEuBu9nwR6YvU5k2gXrgla1jojVtcZ10
bIhXvlu3IF5QA1sS5lg/zQCizE32PXH/NRhViUCxVm9Zh18yndTwfrkmvcQkSTgRzTQu/ryZ2Pwz
Rk0YPMC2RhPAblS3X8GinBjYhqMbdPAu6aS2R1jcV9WAq+Qn9xB0YpNCkYPzTiBwd+WU7T4/DwAX
DYzSo0AVPcfrKBONXMszPdl9GVQgU5C9q9K1tEV39jWJ1kMRjFOsyBMJSqZOwyWWdzGBTtyX2Hwr
ZzcUmu3UwAVnolycAcSdEhLYYZ3ONhWM2EDVaqQQCQ7NrS5EbcSwFgHZNGDzg8CDcbCUDJgdjK3v
X6TWEEHT7AVmQJb7Dex4VYmNQj4/1Ksyhk+uEpKkpYiaZiXSK8ff3fCp6TbGw9s3S5Nv6pK/O5qN
qxz5t/HBbh6j3QLOSpDJk7JcalyCo8IvigkrR5XddtX/GT7Rs2lqi1vaMbVreTaYjIVcIX52fgpI
KQHUbq4/CJgiC3UNGKWsFDPWBGE71wdUouFP1ACSJnMqLpP3+YXNYueU1MfUj6Rlvb8dT0Yl4DOJ
g590TgbNsIBpHG2Mewddr9s5rcpV0q43zLznSvD9iZ4VSAA6yGUpAB5ugEM0P45ctFKrvKWJ5yiV
Sdem2HQJttqNrE41E2LOgI9ib4F6Kq+WtfsQBoRbToIC+GItCgcjUYURW7C9OO2Aksd8PNKdPaJd
ErIhN0JBPr5ybxMjc4mRNhC9RTqAhRit4c2lO7q6AfU9EU2dcL5c74MUzq6DNpiUlKCdrwA355uZ
BQyXPhmsyQtDUij4bq5FFc7pAGVsMI64Vm7g7sfU5ZXAJ0oWQJp8jneEnU7BfTWWFFXqAjkLRtR2
yT3dyFFF9p9d9roh7fp5R9adu5UPurZwcpSekZTWZxrbNiEpJ4i/6VF9xgJC2b327l4ynQSedeUT
3/Pl/HNxsDKDYOeW62NjsCoO9nhtVXXDg1BiPLWPJ0bT89Zc31D2bjOTprlEQQEiJSVIDGygOwpt
hesErZnGa59UloiGH4nsqlkmYjAODMOiPPlkdqeJMRITl7RV/hVbC2l1b2OLiDF0fIlernMcjfAk
PxZid8ZpFH//mJ32IGYTZs6Si1tBoTEMiy/GE3usTmz9AxeTfufvG2fj+m95mPnIdYdZf1x4T1Bj
whi+FvzHZiqi7onaJ9EB8zqdXAPq7oL5j7kMnEr8uM8n8VGpL01i5zdC9bPyhYvG0hJD+rLWbgVX
y7+t7NZ4ztKSWYoObKU7K3uhR4Wb9gZMTSLv5PAsiXikp33XaEeD85KLN1iDTbPmu2K6n1s3mCDN
EfH5FDwVwl9wtvpJUK6yA8wzRSgPpwGHmeOof617foSzkRa1yyf1DIfHErDak4q28GTZKmHgCsR/
dnilSeWwB9zNsFpYniWZYcrL5c4XbmoSYKtz3vq6LJduHe8XwTuKPs7ScuIDdlQv5keonvHB3aCu
Lq8Mx9kPtXcljLNd9tQE2azeEiKdXcNi1yswSPOl8FRLGMPvqp+jCJ0fHZmc4bqfF5uzVyyOH2YB
eVJIj6Z734FhjGx3mGkJkfs07BLK5fzD+eV9rnNU6uTsZWczNbgb/oND0xcrpaFoGp5WRk4HIuft
X/h0xfaQ1nBvycZtGVDa+KdrxYqjswZk3AHJfWASfqP5zQTbWmYj8jbPb4GBKV7PSgcyBS+IH2St
WIN7PNx2Va3d5NM8pZvB9Fwm6YJGrXGblFTXXpfk59ux4DClg8OSr1ZuoynwIIb+D7Ij04Q7JHzh
Vyvy/vEzoCX176thzLR0rHtSv6Qjz5JSe3XKBO8XYN+wV8h5k7pCTw48c558+fAqz07PGm0DIRGg
ZzP39TfWyk376L1nyssp/A7Vz8c4db8CHyegp1YalrEFQ1YIGTXMgCUe1N41+FRxy/DSfjtb11/H
pDuHJNmPUHuwqZ8yb3/tCc3vgE0rGtjt4PPV1EAilZfuaJqvTdGeMpr0MhRjBApzPjEny/u15zDZ
Iyn+OblC1hfS1h63l5MhbOSWEjsQgoI+pZMZrxcJroF/40km4kbougXy2aup7eYrkgWP3srqlE0t
L41fUJK36SWkFigJwdi46CsfkbXjqIfn2/s34qFSVfW86TVHO5ivQvv5K+9W37IjCslsLnt8A6T8
bseOIUjZ3wV2BC+FLDKFGB+9I4fKMJpLVZBrqYInMUBrrgegNRXx+aFRi7K5qwQL5neqZQggOIzz
uWoq55XJV7dc8VvdUqojDWMw5GpmgbMi/7Z0NeRCjCXV4U6IUbtKj+kuBZ4bpNDj8hq+Rb8yObkX
NJbmWnJ4BB2CvjKa4hgY+u/tUEfOFLtgYY959DWamnhUvqUzImSodIjC04nzcbuQbEgorFk810zF
wF9eDJqsSJLRVPEL/8ojuCUb9Ut0sdIDzBRJRwEA3igxYDw0KIemVLYou+xoDlQq1wZEBXPIGWub
0k43BkU9UmmB28xk2M3vVipqY+IbSmBK2BZLmNNsSqiqCSJjCEXmapIYnryvUkLREZBNUjlnBOdh
QY6ZEGm1zNLketIsLwmrOJZsBjmEvMzUJyrlnb9+lql5KCZj19zwBR66bqISe3p3FTT82D45sQhy
UOOQrF02QV9TRj1BLu9pasttwYmbyDsu7VtHerocTfOBHb+7+kFG8c2ujA4ejrGUrF9f7b4kJC6p
GOQYDfxLGl8ddMcBUdEROxEqLZ5B1QiOQmJSrnxJLdnRukxnT7doTziwHg2PQ0/fdO0cjZ3X9HBa
TcFJXaCV4oMmRjbE2xBKtniKPk0ES82wpCWh1xAcCFSibgiLAx3pwiE1lTo0VAf7OtKsVCwVSbWQ
H79VTk+U5P0fWrQQFv5XsXYLG32ty4JkxTQhGpU5chWj13PSZjT+M4A/1C91xfZYmLiuuWaz3pbE
IKeowetQyuFmukl97VKkk0BA/T7XuFh8SEmJHLuAFIshlgGl4FPfQ4k83QvXwr5NR07uOriTFUoP
0TRT2lSP9d7vB5JtVz2zMvJZ0mPxZv1funfsXJpZjHJbDa3lpwOB4l1Q2zHzP/8FVChJVjSRDCss
s48ESBhZqjvP5Uod3eBmtreV4iWaGN5hzstNh2aIrVFH5ZK3TptA5WP1PdcRasCl8QdC2ob0kTxu
LWshx+/49NehuQz8CU/MyC7yaVX4uj8N621S0I/Ww/tkQBu3yRZDELE6zDAQ4Dj2wG3UbJ7zNT7z
DkQ27AuLdIna6r2fVPNUOHHo/S1rv8A1enhQXlnvHndMOCIGgiz8S+K4jZZsl5/YrmXx9jwaXFHs
2GjF/pKnRQWXL4oZnZbyDzaFsWFeoI/JlGyO9EOc/GWI74CBIJvgHPN9woaezVdjMahnClsdjyJV
t33tRjflpq08Gv/CsgxJtAuYPP7wwzmUy6rG8ivL26OxT6A0lFxBzTQcSChZBHMYGRbVyaS2hcY9
jcGL52JbB/EeIL4HeKsqL3JWp5v5XcUyhm1hqgvm+jhVe1d1UMZOnDY0ALybDfDuljGtUiCOqUjs
Sh8uPlJw0p413hznzKncjh3F2yDufVPTlxLaDjNCOfX1Hh1lCRxLDyO2CzOlEij+QF6JVEXPbdwJ
ts18p5CYZ/ueaVPSiQGwG+nh1OLW0ECPIquKMuDa4gYqQhF662qWlwZA/YA6YWrWYOxC7uCq+VyG
prvuV2Rki9KQoVBYdKfP9w4l0LccWAp7hITSwMoWXafPfmXTUOVn5wQFF0fwUwOwBgJRpLc0ghwe
2HekxZuTFs3YfXUxYfbxw7E8BLyl2IcWTRee3Qsi7SMcLM7S7UTR6AksB/b4NJrKcvXTVrujfC4S
5cG8Uit+s56U7GR6Ak4hqYk9AFm6fROzPCusEk6vXzbQWoJiE77RM8vQXoYkFiVVNZVD9XplcYNk
zcyDZebW8k5ayvPxOvFSAuL2CqiOi0UOvPbow5tzpG6t+E9giTAe4r/1KZJDToE5aJv9nzd6Ehod
QBQ7OeOJCQS578pCd5XH5+GJ+bKNzebPgXoWrKxVH2aSBQt+6Ft1CJqfAfqhrbozawf5XROrxbjv
/jBy6BM/Ky2IZPG6/UC8d90VZU0ipWglRR56Uw909Mc7YfzLvJtZNn/Uzvw30J0r3DmxAK+9f9G2
uqLwP/Y3PQAxJmqpFMdRb5H0GzzavsZ3ECxgy5x0OcHUPaXwzXiwP4U4nVl+DaM9Dz2BslnsgzH7
ZUK2kouRSXA39PrT8EgQXPkMO+O49BuN6G7IzELa4EeoRH0v05uB/byqhNMy/qg9q/5hVhk31Ld1
6HL+Qj6YsERP3ZKWtY4WEqpYXiscaTHZFtN8QVbei23cUdeMC1TU2rUY3ZgDNbcgO1CD3ffrBksw
IRZcnSWqd2koKYYhYrGXudUHt1enO9SLZJQb8MJgAMzPiHFJ6dmFTMrTx45bf0hUmfirMN+6QeIM
St44qRa4JV5AVXBfnflqEX49qRWlSMmx1XAS3IEZvMi24RZACWcnzPMdLbxMfIZUVMyt/nva34sF
ZM4n524GVUKOwR2BXBcUK5ufGigV9whOLz6HVcJ1cHrjyZjhnf7vgzkD1x4MiCuazpdbaCIYZRCY
QIhvZlrprTjh5fJhHijkyUqWXAgDtJblyz1jZ2FDb4NmMgz2p6MeYvkfx8Z18dlN9tI4kd/v/oBx
EJjv/r5M/XIvTTIpnDfPWejzeEuLLokt5fk6h7ISQCpgje/Lb3/XJQrifYT2kyWG9HfhsMchcKtm
/JSdt/bRxsauBoP/ucCLjGnsiDjUbaw5AFY+HDRFpORa1oscxdKQBEX7ny8Pw5As/AcB1taqRuQs
HucEpTSldkgJ8Be2bDZFx5XIsPu12GNFfMZvQIjMo2Eo+vfbmcD/mcP5iKsH9YBYx4oO/WxfcGfI
by6wQuXpCc4jnGT1zy/RXQ5AU2LZLZQfe3wpQ5hv7vb3pei5wgg/CX0dfqtzIhqPMr4qwPCmBoO2
bIJQIUVkXyRGJyj7OsaWfnYuhoffAFCJVaYHMrKQJ7RWD2LTfNe23L5j8IVXfDOqC1+EW6s+IdcG
uQ1tzbfzue0j+kpImsKreFDZOAQXEAWA3nzJVVpO3r9n9g3GToi5uxAP+A7cv6M47H5MGwZnNK7o
6EGi9r9vYbKHqD5sAp2uwVR4Pa0qPJZ75JaJzoRV2GScT09kLFeJznC5Flp6tNTEYhSG+v//QTV5
AMRMmiHcLK6K0ubO9QAyYS7WjwGMqMrkuHsm9hgBquEm0rbri4AqNL0TsOg2cGv53CDNwY+uksIP
JrB179KU3XxGLPVyxnUlG0nPWvhb03mOibxmFQiwCy82fI0QbU7HKfcvOJNT49wkD6JmSl0sFcxy
/yqnFTRxo682ZyHrtqmXY0b1VtZQ1DxqE5NsyxS8wfZaAPrAnobNjznNOrYNXAYCqayIfhp4rqqL
NJiOuljsKYFKmLYN/RcZoE44UzkH4rmetx1WALvk8g9eO5NTa+meuvIC7pcRRfb3u5Uy+oNW9ClI
+94bHthOP+LU1npXXLP13W1/HEGlyWweZS7ZWfI6h/dWcuxER35KWod/+PeqinxSNMM6oLGVqzjh
MBDxZMNWe20b+pKtLnqhR2n/OBfeqMxCBF3WmMIsWmEGkuYXR+4nL8Q2nOn6PQtarlEVS5XMdU7p
k80jYXYodvRmFOzY7nvmjtoUZ10wuqWLhJZtwTJ9gj2ls294+M+8CN9j/2NMQqx1dPdqWBWgys2Z
Ko8jJn7yuC4EmKXJj36nd/1FOGYLkj2bfRaeFBfq0BX6X7msKG0fDFBcaYqqz6sAL8Sp4RL89ndS
mu7PiDN35LmkAHtjPUZF7Brn4F/Rhqnty13og8NTEpFtUWFKw5mzrvGPXhbWVsHfBQbpHNY6mwgy
TDzdhxXLmJ2oPQNNFkejH39IeAPRRiqUyx/VZDLXGHwheJ+f7H3e6O6k8+JxQ4UoPh7pzVQMu6km
Lfw8Dmdmi8AhlOF+BQfnDLJDbNON/VILhjI2pZcnav610qx1B3sBs8eOcI8Jw7quqjpuMSfNHuwe
O3iLOXxNZ4VBBpK50QRR0ObGGcWn6imfA65AvB8PdB2YF0KnzjrdY5KpMgk6UrvZtoWd0MH+YPaT
4rEaB8OCzhLqVGewP65y762xoW2TuSGr0e8zfsviVbv9TKEOyiHMxQmQPWBH9ARBQmRWTzbw03sJ
wACexFIFUSa1p1Vl4KvF6cPqNRUcUUDD+cZwgHsnjdNIfnkoef4D15r0H1S2f7xrhHUGxPMAgsnz
c7cveaZTlL3pE59vIBbFX1TPyNqfM7CJt4N5zm/xFe9pKYJrnglbvise6d3zVNmDC3HMhKLDeoJt
ew1BUp+JSrlqMUup4xoN6GNa6b++nZrRp1MXnjD9yKt237AMP1aBCRbgTf3RyAa4NEIVOJf9xmjf
hfjjpiwdc7NjFigMcUUuU+H4W4o2m+ZHDOWHu8KWo88Oyl39bI5ZxRHPidAZiMlyjgICRf4O7YDx
40bI7JySdhC0af1RPBJeqa3S/Ebzjw1esI4MNfxCtArkie4URpzN7R4IXtckJCwVmBcHXfrmrsVa
X8DZXaUgf3xbXNJ6baq9wFDEvikLXUWg80jDFdbO/vK7Qw/q84M6GJMB3HhKcBMohk6NIQ6DbFyk
JzUD1YuOpRifHIlzNTxidDW5FlyS8d1AX3bcKV+csoV7ndOmXXjdF1mrbBJypdYTRe+sAiDqNL/Z
ihFndt/fBiw5rdAzp5HmlQRF7wqGf8hCUxVcLkQJh8XnjujmxokpUfulGNpwyxn+a38YkpJTo+P3
ebuU6h/wKwJWq3/tfI3Er57c4Prcij190R8poeOfOvyJJInJyaMrtELfcKT91ekh7R/CGfVv+GzX
tUmw67qt9WHfn4aECzTp8sXaNIqp7tgxxV5KUZ9qxgTaiRqYqwBqsdYbLcGg823dnQ6CRqnXOugW
HNbALVinhFS314sAtyaqzh2JJUYz0HduI0EL/1SrJ06uRO1cEUJq8hIBGYZcoO9LyNVF8h+u18Bt
71OL8avd5kHIlMg16fTo46YxHS0nsGwakboL6I74x8ZEdEtkDhuQMmhBvyQOs2ADafbDdb5qwZlK
dokvAQap56zoaeLYJbyLyCTxmF8RhCsp3OtIWiRyLnLwafMfAzGAG0/tgfzHt/ogZMgmMQtb1GWL
vWa0v8GWtYbYYKZF4sHmjlPOmK8+N65K+g/Wc4WVh2/7V2PlL5G9UFJ57lzStOGABZtjQSzw3o1X
Mp/UDoYyA4dTt8HFvRuHQ9+aWEhdmluEN0GCTNUDLWNBu0njO/KmZNsN2qlMlAkNHrzCr7h9fkLY
GAbaSWXqliOMo3RjE0UtHHKLLqGmzPi/qXfDrioHNk0RZId+/nCQLG1hkrX2CO2vyWo+f6GqWadP
45/IKdzDt1mktnkGOOX9sxGfg2qf/SjQFzKQ22MOZF+HXjPhCNnt/TmQeULAqg5SAPm1hZ1jcC38
A87Ywjrab5v1YLchEmuRMWq/kqj9/KLfEUOS7PxJivncHRpkBXDgGb+doCllYlB2kOcZRTyJOdlc
Beexo7q7HNsE79998XbDk/eYOA9CNtdQnLFNwlttlgEg7j4EL3ShlFUSsepRGTaKjymswwCW6f79
fBE+sQQYhHZMzz9BOxZG+Z+/dOho3p3rpjgkgZE5M/+iu6L6iKe6mzaQXb3UjCkG20rGbCmIEWa9
0u6fkVBSMM/ytL6lXW7HPcfg0hMEz11iTImz6bVp1/HJ9wDqT5mhyxhZ8A7MaN8Qyh1eAM9/gjjA
W4O5p3FygPzQLKoPJ6AAEL5/4548b19xSOdUBo6Xx9rBe07IDYngQNYlU+bj3A3jhLv5xB3ZEZQE
UI2EfGofZP/ibS03rBmslsFC4g16Z5dkTT+CBDaIZONL978zuyhQui2AuGOMbK6Txq3N+yiXyjR3
fWPlgUqxD8FmhCQRnGWSKqAsKYTcXtE9bjeD7o0mfWj2gNHCRako9ID6iYvBw1jbd7vFqM/Xe884
Rq5kp8TA4YC2CvHzstHnqE8WzBQOzysiP2wu90RImbBiReDF5+9SEoefGk8HVCITpRHOhIHAWqME
vs+06Z2ajEFZvbQPO9IflNAKahXt11it4ixpMP0ExuXPlbhvPbNhpdv1u93Td0AFrFtozoZSxBq3
hPkwgVZ7i2TeWVDdOgQKUuEYCn6ziNdtT7MRlmVpITN6VXB2VY30dnWjp0gs030ox/EDGnN7Fi+H
GA0nzziChGh2P/idKXWYYNm/LF6HRv3AEfQHCIwr3L+V6bkviozNyZfEQrCNKa1v5ixvYRCSPXr8
ECRXF8A2UibqAevBDEgrcd1Uc9Bog882N5s3i1T+gU7Epdwhy6cqd4X8bj7IwRLcYbNEVJEeW7Vt
aRIfYZm9LsCoe9VkKDyFT7pnjdnySvksZIvQJsexd8Pk5iRNtutIoilvwRRjHotlRsEuyP0KI2/i
OOL3Jz9iW6iiytvWlNp3fgyeLaWdlYjFe2osEAK0ocJFz8Yxje8Y0Q/6Wn64ZeIqrfKCXTEzJaxH
3zPGz4W6f5BwblPALQzo7+Z5owpznlqdr/59FRdjTAWgjUjR4140tSDTkMwTth/Jgw1pRypSi58a
AQJw0nkgtySzWh7Kk15OaS5H0fcYtTMJyl0zcb9nFK3v4Y4yGAwLu6MrzFFEY9QZygJ2VMigL4iu
jegQn5Pm4a2dN5DF4xJinC5hiNrByrI5AcCg/H5Tjn2WwHFR/fLH/eXm1NdYlffL5li3je2KgA+y
Zutv5OSWkd6zlsYENn6jSbe3lsw7gpwkwSEB3iLQ6+DTDi4ztrsANRkEUBagxalTXgqCfIRa4iSt
4O56MermFkVQrHMdVsGD71/RECNluBTYS3x1dftxltjEVE0iYPJjFG+Ks9D731k6qvREugG0cYPB
YLAJOfbdUFZPEhKnvyKogYOTUXAVRsNYTv/za6Wz/T+Tb4oevRwO+YZD/qMfJtz7AehTqxeV+9fv
89aFipLAeeyztpY4As8msqDlsi0xTRAL+7Xo3nXQENCcgWY5I5BXWjnW1bBKtMh5zi3XGc7EEeXO
6DH5TT0wCPOKGrspLms4hOtAasQHGukokcGKLvbPmM6GQzUn97+IqeeScIpgjskoRyPgAfGPhm6j
vr5pLqfBpH9PQE1Pwu0iNpO86XB/wlWQhJUDawM7YtQRqm3QmEEt2G+GraIDIlPWYdlaS5SUYcqg
uGFiVDHjBS/kW1QoM+i5akYunaK1yB8gh3fwWDFhP+wpg9iQ9/mtVCyA7A5HA0teVwrnhubXuhE1
+ssbg3HCoobCciySYzO21JeYzzH51hH/un4YJcRS1/IqrGswlSfhxqU6UaObWgx/ZRsVzulhlMvA
YUL9oYwhsXr0egWjZIq1kn7D6psWhwlPORk9WqIHgcSkfJU7Mn9QeM9BEdsV3DDJA9TasFeRCgfH
e9aUYuYAoG6gYEHx66Y+4XBuZjPMquQAkDWtkPkCXDfAO3f15nvx/s8DLTlEiTGo8BuzF6BOFJ6h
69QWUpOlhBNhvzdXj/uiAfyL/jRw0b2CeJYO/r0+APzFl2qBOoi+idZbPQWBK2XbmNUfLTqL6F10
KP7uMUNcUNqboIhWuNvWQHA94R3eApWu8vof4JPtT6epTSW8oI6KXanFAJKOZkQ+XQ9GOH1qs7pZ
CrUXQvfJoYRmKK1JsGJHZVCN8d2Z12qrrmsn32Mgn4qOnJyP/WwAdtPt/YVxCh4fI2kUJ6OxpbeN
L20b6/1An7qvfGKuoLOhg5mfNzglgUegcNknxCLPkX8X3efTtbnU9gtSg6ds8+NaIW43iMeTGwIH
0OijW2HQ82lJ/YQTIykl5FXzxStW4q68jsc8d6TQuuxzMogNOmUHpaD9y2Onk3MVd1qS+a8CzJUt
RWMubLDzdUgvgArYapzErkwGFhDUw/f4cmc50zyCqKz5broKMw/C+BrN67O5/AhEk18JJZqOd6RJ
V/c3wC7U1HS8lHPnBOBTPQrbUdP9rUOCAeO3c/ZFs6iktjJWczN6cO7ekEQvDPETYbxgGJ5g08Qr
r496C6b2hBK/YWUcnJL3C4Qnb1LI9sYQ4a+XiwhBZwLyDBYT7XW4CyIJXGtM5mJ35W9moOSt7tX9
1CnZkpThASdNTX1UqTNOyzZiQQmMtjyzMNW09XzckJuxiW84qk4bmB0WtgB4vD/XhMRqZE1F9y9H
QwywmNHvN6PAWuPD7yTBNXi6dJZ6B5hKdvrBHE7gHT051KVUb6OhjeQmCSoIUt42bMcYjZDx8e0c
5q9FavzWpiQBpBlYfG95q2LNGfruvyA240yPWBC3it99x81ZeQ1yQ16Osub9mvwEd1HBDhj7bW6h
Ydg3rj2Wb8OtdK8r33Dn/fW/i9D3Ex70YbhZMUIw3+ZnDBKeA2W3nVS8ADNlBQ3zgGZPaspvMi8y
SK78AVIQvlLJqexRXLVg+Zm4XNdqnXKS4BO0SiDPDWQML+U6o/j6XsMZGV9WPYS4TvWQg6WnFnkO
VJcUlx1OMzCWrUdMq5Sb9khe8uUsWoa3939I7nfjvHF2vTCL89cLpsV6JKJRY7IUr8og5/xsk4Ra
qqFUXB8gOHX3ctXHhnACobHZ5B8xJX6wFv1Y/NakHji7aWq2BwR9I1Q7AWlw4MUr0w/5rtU0wTXp
dkETAFjJtyUf3ha5ItB36VnieMwko0IxgiWJdux7z98HkmcU8jGxb90Sf05Qd2dfNcYNXw+saiT9
oE8zQGvBlRBBQCL7n2Jc+02Cmt4m2cz/8qChOvHz4ePDHh7AqUlRNviGtYKzcR+1saKeDNoJzleh
wnMH7t8LXdkYJtHzLbe1d0WuAEzLPH3ahS3/Axob2Ty9LENpHKljXPt/XSRQPZWqXgq8G4POoq4Q
V5LyeQYgnetG5zJ2TcyionLtTJwJJSBb0VW/tNXDFvU2v+QuRuX+1hSZcpV3BN1lG85GsETDHZCQ
/qHrrxq9KfHuvOLIlquTZUP2A5SJanwl53DjW/hlwNfaZTrTbKjnqOFZcZ58UiXn8jiH1D4wco+6
TcKdR23psDY7HXndwS1RQc+DfmpAE7pRRTiReEjbpQ54xourkf+edLY37O5FTJi/Ze4f5BYk2+yu
bJw7+2ooj4UUZonFw3nVnqPWoYL6EoZPAErCsMbEMYjLP7j16MJCeK4cHJ5VZLJJEleFkZedC2RB
K24iNONcc8x4ozuSbQ7kq82x/Mgip4YYFjkBzyNFyrCxwiip2O0G8i/MTrC94lUXp3UgS/7kaR6s
OAPRYYZvnYFYN41IQnROM2hCKZmuT7vLZ4nCvyMjrSJIqq1jJvMuQyvuNkOXdG/kNA0Kw/XVMRwn
eKn9UI1/GdJSsPq7FfOH5hU5H38/LKVe4l+Yn/ShmsfwrEcCR7nsl2EnY1ap51CADvkwZ/gYLsjF
c9j4qc9MaiA2ghjUEoiR1G1bThR9HYGXAgsYZvQjeUPCim0WHsdfgut5WR5dlywef/VdgHeHPcAW
X/JUr8kjrrA+N5Bi5ADscy8CS701donclNDOGJtswxAz3TiSDSDvcAj3WtxV2qwDOjrEqXAtdZCt
0mN6iWvApOrgXzhOp70DMUlcMNicIPPC8Obz718EQrsaL9TJbjShtvkzegwqUTfnSqafFexknQgc
WZzEXNs0He2meJbyFRCVGWUz2894mmWifJM3dwU+YPdfW4LoM73xpa2yF8jye3uc+Nxz6W/jgc7u
IpwUqn0OTvmqDojN/2aYuPFT3Y8g/OPQOOVu9+Ijxik3/H65+btSNfh611FmbFLSGKP8l/7QMsmS
Bf7YsTg8obzyl3bfyvz5gpngMfWN/NHs9wlVIiCFpyK2QwRdk0hSh5nSEl1zwK962ld0zCXjjDxJ
FnDPh04i1l4Nab7jpYn3UIf2E0ICr1mJGmiUknOONMBfdi3Ki10Qj/W5JDCE6t7UzHVLPWE6Nwcn
ctN0n+j7x+z8pYVSbCZRZFujIdas+q2sUGOSjnEvTRmO/Wg4LYC2im6RaO3hMpfxyTtWQvnjGNtC
fe+wtw3IDJvuytFpPQ5Rq/s3JR2RFUCerXXidPaheIO/W4dLIqJzxYTGuXVHhVOFXYxFIP/z09WJ
z38buEAkLJCiT0HDNmebOTF/6FxDZrB46frXIgZ/CpMYxI84qTSGMzfZjKDo92HvFOwEYDnr28AO
6fWvbsixo2xkQiOSV2nl7w/lvo0lg4vP8LyoK1w1T7he5Y6jH052Xd+qf3+uEwKuYXtmP1wQyyoa
7pxKNO7WaueNiXXkNsP+5le5u2PYdz/S0ebsXKy7TzawyjzwsYOMfT9YdkmDTyU5ATWVe/MaKVW8
PZCxqp7sHHVUPIwfjA3FHzrg74IE6IOxxhdMoAg3pSeXIWdBU0m9NxEVmkukqEcYVazY2mxeqgZq
gmzmlVUlizj3RWwgjZJGmQ1vl4cyBmB7AkWjvecHY6vThbBL3xkMx/qi6eJyWJajPL3SJClaPtWc
gBZ92ZwNC3/kokACGRht04mlIF4Wi19w8aj3PrQXd4Of/WjwADRDiwss5Jq7HDmBPFBO7H9cXDb0
0TA+Cg4q9qmJWi95eyPLmhKeZJJqJmpPM4hw4z6xl33ZArJ3WKhaan/J7SgupFh1KpvRVHMYOg9+
HJbeDDvsS6FcrpJHyVciLcwqa+DHWsUyGJSzwoopwEARfhdx7MjefF8fNzAeJBR0qp0680ZMwgnO
gkdwtL4/8YOIyq+ZCybWk1XOPw+upKik0M3cLLuphq1D3r6QuSiW6CbaBlMDeJUsWw9UqK0v66b/
RRsWRsBq/Fz2tMAlx8vbClGUtQv639hsXJdc8qybvdiBve72ma1dQeks18KHN5QEQJsDcRJMgRLX
6ONymOFny+PEZrw2j6wAWspiz10a+wlOZywjkopWDKaELPjDNKCNsGl72szGhbYsqUJyXIlzRbuO
6k1YdJeBAtM0gIurdfMWxVYL4HX5TDO30wyYNTlUe4dne9s1M1rxRRyttrpttPI7EUNEmM5WbKGg
hj1/eDwps1tH0hGK19AGSsPo5yNmVhHA9s3jROwS8V2a2kWf2ozGR9zv1Mzh1CXg5OD+/772eTPv
oKBo6nDRxrvxhkwRgDhs5cplWo2htomdoRvWpq5jTdg9Lx16R1WOUdW8s+iM92KIdm0uvFMt68Lo
+kwcZSqSMZE0VjVGJmTA46rtONba+t22hi2heb7/eS/amK4BX11pSrFc2q4LDKHNFfgA1RJQLF+G
u91tMYNuNFtv6lJZ+j65VHQIQRTOE5raM0KxI2sKKuJOxs6ROrfOiQsMh2+0j9heX/2wsNaUR7q0
VyNEth0ykuIQQWSO5iVaKEk4hKnPwOBtAghvF2R5kAinxgvTe3VCPoF0ZKKsVQZsvdV4AViQR25r
vdBoSvWQoLWi5H88EG4k/KAoPd6sGsQF11QyMlHTv99AIkVAMJD/dyncFZWNVnt5DFi3zjihu8/x
N3gkZ2CsSQ969QY0x8UJyVx8+x/+IBCsbjfpNuJxJ1mrP9btaREX7o+5XKtcaET+TJGDJJIPzxf0
/4Wjjck05rNQ0+b9DFJqKth0sdRuV3/SLR2SR4nLjym3c7zJNYE9HB9ggDByswSV4v0eGgmeqLPG
S43S9Kp29+9kwnFLrdA+HJKJEIe1SSP+DIHouWdPDM6C3soVdfkP5hk8kb2P+c4hzNaTWln/LhHK
hoQwuyMaiORwC00WDulj9i3W7jJQN+8ULp9aCLz+cOh3JRl4ur1AkK+oxSwHkbD9tTK+syMueXZY
PCH+2cZAs9PEnGcxWEkvtfEgaOqYYF5N9wHqFDO6z3NXL/1+Xi+J4qB6rXDrsMxcX8K4O1DTpfiL
wmBWZN47vEnaDHnFMccVQtSMhZ8efEvnxx8DpkkxkT0Dtnpi88YCiasM5vs82SF2O4AgiQLXYsag
2WeNWDRRlXCadbyvPP85tWSGssZhDm69w2TOaOTDWLQjsGriGPl779JfAvZcC1T9BKwIjWA6pB1D
M0uXLsb9shlejDCrV/NT1YPEKmw3PzLv1Q3ot/Uj/qmX+UOAuMPPsuCNwV+xAtazc/RX+KymU0w1
W7IesJ/9W2SnAaqriVtT6md9OQTUiHxeHbhQAdQNJZn74zLVq4CVsyOhtoPnFwke7/MOrR110698
kIzh2y/TFDXmrl7/1zZuOuzIF6wRTkEUUBXfwGQAzvqyS+0OuDnFws2z9fZmKO7gEKObKEUlKDfj
lSxOviCSaut1CqejUN4W5ciImyO2mCfwlbRqZ/1ct6p5fF1dHIAH+WS+78E7D5K8QOILZ/oHBihZ
gEy1WgcpvLEjji/kTOgKmLwrbmy7m8S9VXkgBfeMYWshZvqaPAyySRpOYwTftJN+OLRStmMQJvb8
3uRlOCzV3jVBNbQAtTyiWMfvrYmCVajKUjfsCkCxNa0rvYxkhxURvX9fzswmRza5b9sA33j9XPTh
J9xqhMTU6HsdJwypnyw0Qv7kLi3nJbS6KBeztTs9BPG9levMJrtOQQT4hcK1ta/O+mns2IPCsBaE
lA/um8BaxbvAJ7stOtf/qGHU/p85Nol8j/p7+f4vKg3Ti34tuOip4PMdG33cSQBvGJ8xUyrYMY+1
38Y64qy/Sfi2UK7vICRTQRdxEAxfglKFCgGuWDFF7GXgjZ9W8D+3sNMSS2SM9J1SG2j75Gwj/Stv
UMnI884TPexgpkqg9EuNrswFyRyGSBiiJMXvcYIKtg5qlkjG+nN7Cm5rVv3xS6xTnvy4jVJV0F8o
8Ek5yMLnPXBbyu81aFFEr+J0bx5qO89w3YQ3HZJ6EDHMknKCl/cCoAZtIS1WdJx0nmHWmEQKuXnF
cSHJNmgZcrzu3XLuDpMrMIsPdgYQ4WTXALLaOzjlrPpm7QsqXqimyyTpGXNFytLl9lAKAL9uhOpb
ZPzPTtgln8tjdw/dmV4o1GtETpBzGrBFoLux4HB8FJXdzxGTsVCiukvBMgUoBaFiQ6wYe7lOIxJP
lx1pbejgQERk+v5J082xgxGuaUIrqdB17JJ74gjfxb0nsLqmv485KVql9M9vRGcr28rFI3KlX5HK
RCmfuNYhzOvPcf/ZOvs9Rk7nQD7cYoW7CslMmujTSKoJirV++quga0kc1yhFDbK4imRO6gmfEOvf
RZ8sGp1RJWLw7xH0YF+DuEkSPTQpx7eU9dIpzyr1qay54FSiD7FzwTEtBicQgbOQ2vrDT/lGhcEc
c7XA5SMv9wWJaI80iP384mzu9ez7DoMqt+8Fv0oxaWaYxWOHC1i9cHCZu8ZkLZ4PXaV+QLaqkaEc
PHlTkgNbTqlIPReVA4+xcOOBwqA2VchHj1dQG5/viujc10XczQ0S4XyAmtTbbrL3hh4h0Irf5cS/
OetF6lLYlkKviqgwIJRt3mDkGvuQDMK4xtwnUNzvF5qGU+UgLo8NUnlCG7XnIw61v9+Rhm3+YrZr
AbgTH5RBFC9tfz8v90SAkdlRxtTKARxh8yqk25VKHXD9MNqUU6vvfQ4whofe1ltWJ3xE3d112796
FZTjI2g08bsZOmqjxyPsIsjFS7rdVJB0L7W2rZrl4Iw6GHPOD7e0fA1EdAbIxQTKPWTeTczoQ2q7
wVs6sNXabNy9wja3u5iXEAeTMNbCIBOWUEAsm5PmOnktpZKUwtcfXAdpbSqnCPU9uLCSswf+lAqX
xUM83qY9ZTgvLcbyM2JeBKayZTV2r/ZbzbJcCKq4RTyGQ7aFq9vnCFjNrOoSpW8d93kFYy2QBSVn
nulhn7Z7JBqE4XhD7aG89ubTYlTni037VM8NAawSxGoiqA3aOWsoDj/QTx1hqkxxIOuKx4Z9H7sg
QFAeHy+eFladW+SjqNjXyZWT7Mb23Tb5ekxxsEZsTRIzOBmtOtv5YwX+QZP4yb+C1dkx8tk5kBDr
EuzBao5QZ4bezEkNhe3TTvuxRkS7a4Bh937KDvCvyPf8P1zWiouvo+yBPgd10EUJACmfiqZeogfG
pyvoKQpxgcx1f6xxY3wMc5AViwutq2a9slPCW4tjwKHqOdg2ecE9J8VQZ3UuWFEVQ//d4wgJk44l
wW1zX/mUmhpvJnUe4vVdsqCKZE+51l2BSO4XX0LRqUeF6XriJqORDFic7udTuMYyw8rYKaSY1t5f
QWs3EKJ+tUUXE6Kcj0F7CPhIJI6rc6AXbF7Ul9cQQrXp8OxuDqGO7RI0zPKVW77wWpPE7sqyUxOO
xLnmVPXJPeI3cAXHTVkHx3uTG+HmFgEIzupCFW6m0jnDLaqoNUUzlVO+YSHd4ZT4Yh5kHA+gXRtJ
fHeFkj1oUpHS7vOPIL9ymm6pA4OXt0UTIghBr6vpnuDQsrnaxWN50P9ZwJKUHIxcGcMFK62xdXVZ
xtsWpTqpRjGEltMf6pXA4tT+O/4CmZQBuC4e8aGxoTlhHIZJJ2emio8+yRF0MicMpd8s5bEoxBnz
1IMFlU1PmThUDzIzNCBej0piSPmRxLHX1mIGDSeaVihRNDTlj24tdUhJ9IxcJfwVccQjWKQT3s7p
nvIYwqMK307fW9FLkGwAPThy/V7r+VrawMlIDEK1oBImg1IXv52f7XYTGnK1UQ/qbCtuoRhcpODo
ntL2rfZ7D7NddH5C+QQLB+9PShX5bUyMywCZnQxIxSIMLiPWSmdh6zoPP/Em3dY0k+Fs+omV+Tt8
5Ri30jM8CXcDegKSprImzmds/boSHGgpxEvUlJarT26h/MB91YovlNxVOg0ZBudYro8j/I/FExTM
M5c4NOyAjApB+stBj2e8LccvmW7FpILwnWckzLzgXo4/KGXdGS7SqBXWS6jYMk8STo/TTb3AMg2g
D5Hqv99ZzHuW9i+/u1XJ740bPDtVD6OCBZ2EWbphrEK3Afx2uLYKGMvWhPJ3oaddI527e0UmRmpY
4s5Th2bQt5g3gU/oTW/r/nX9ReFpK7Prj2B+c6Tkc1KH/5DFp19YyoPNKUUnSw0w44jI+4uTq4gs
AthkAI+setFRgSyIC8TReSLDEPn4GKBjAJaf92ZACZIUu9rgHCDVDTGe8pNrLyn2DqPCnALtt1ug
5cqvRu+jzI5AFxtRwWASL/X63+ivZSuOJmdHG4swdOyG6xHNUlesA8UBtvvrp15sEmfUuPtzZL4E
dWjVzmfuIXqbUawDaPnxtAZg7YaR+Kpdm0BtVgpfOyBgHcmrhJcgMRn5XBUJWnUorjhJtiZdd4CR
2kVZOfeeBxv+u/cyeGGc0RAIloCkp4AZSSkBDM4g8m23xavYOkzhmtmFVSJIGbXjxrnz6GtqI1aN
51CuhCOIARFPpSDPr/Hv0MDGuztaCLISm0Q9Z64jhp/m5ugmLR3b6x15UlwpQTt4b+zIhW/RlYP0
JlZ6VESq+WCVGQg3vA1jIOXb0KTX/0cOhpul0ClJD1bQy0fo7pzSQyc0c5pmgTKry1la9cR9NzM9
ia3ItmtNu7cw/KZ83Ij/jHfomlGmBlklhteVGGca3uuWycuNq7iweDEAU4w4BlMLkUDwjuFXFsrF
+CAimTU8oCfwgjocwRryDXk3UqZf5vPry7nkDsIuxPuPNhiCK2VaC860vLoZzZZwz1Bv2gJwR88s
6Wn5jXe3+l3nSMnAof6zyInB2YF3BbpYtML28IvXlqGT2HYWg0GBy3S4BvSKZiawlw1GQSoAqY4u
UhDfNKxdALXzyxUVM9GDeeNe94v63km1Sih43D67j3XUacCrNwt6KdLhUQgienk8qcKWkWU5iTK8
iyZgLBYkP6bLGz6ZrKBjEJAF6Q9YhTtTwUv0DkDcDMmxik9RdsmxJPqt7YL++4twlucOsyExW7mT
KGkQiyeA0Ftg0rRpLeCtRoR4nd7DRHLBaB+xGJVZKSoR8MBmIm02uwBrfSt1s8bM7FcvdWe0xsy5
o9heKad6yvxesCXvnhI4c554xPcMjAFwBfu28TqQWGL8nS/UpAPI6ThBbvQ7fIczfRkaN7vFRdIK
oD4KcGnfqTvMyS2MUbqi6gDQJpFUdF8lANcvtEchh0/ryBSBpzv99lpd80/aR6NtsFpSQ1TGjbLV
OJQfm0eSMhgGeXaEuUwpiYXY89TrdpsWc4pcHKSobVUi4i2mM5LIgac/zcOmug8a/IOP651q7veG
cSlRQeQGOVZA4kAX5PIhPknu31+j2WFfxdEZGn+88lIAMxPjMSLAfa6VxnxFEzTfQfFg0vt7193W
Mpp7YkEEzOcZEqyCULAxbeykXbzvlFv9x4KLxkB/JV+Nd3QZb9PVaOZzLBMegLiEmvd8GUYshl9Z
zbSquMQWTmGvg+WOVIcG1jKTfByui9hGwF0KM8GEISuDmfEyHGBDxcqWboFqSl5JeVai0H4OyzMa
hmbSza95R3y7pn/3hET7rtVVrqSB7VrWDA1Jq8jMQd9/YyyedLx8MN8GfhnEWztaPmKSQ2AQYWGz
SMuSVv/EsD4blSEeWcji8RSGRAvFtZeTNywdod7FyEMo10NZQJ1uqySf01Kgewk1Cn7dhOI+iL5w
WjlRcc2AhZZ7GA5msRxYU8a3tSJmNfp79Uk4nUUvL1fyB7iKX3w7O/XN8cIkF6uo0/LuV9s4fXYz
JJL+es/4Y2NMzbv+ylFlu/yD5D8R2UE15yMLUgbJIavLqArtrfCP/OeYmqVGVfju3TFhquAJMmEO
omHXOaNdcPkfrdzBZTwSWUq1gxU/EWft0WGp1gg2CAjyome+vaVfJLypbYYHP0BNmdDPcF4kyfvj
Eq/YFeCDOsp63+aXgVnO6bs4jHjiETF7GUTI9ksZ5btCRIL5UtHGWA864TxJIObgjwxuXop4ILFw
Nhs2Dwa7ibH/P0nGCLQm10gwbBIgrTimg3TszeB4u6iTyMGrk/1iuYumyixLiWR8o72u3WZpCq1K
h3humS1p/RElc6LvaHWRtpQpwsMOCI05JUXUcH9ymgBbr2I8QyR6NuChvaIfeb5TrT9yLhR0k8nH
2VJS+/GEmBuZ8glWLnjL6EP+PfdtRcqFde+EYwf3ijMhWC6hfUIimSuJmknzMaT9ozjebUsjzAKn
EfVrzLSQwnxrwhZEij2PR8wghvQXjdtb4Ncxk9Loi918t9C9pqbfSeg+skq9vWzLkFzkeubIvh9R
AeyVvXN3191eBmM5CeGUoIoMlPLGGxIQpvvFAojBrWVemn5QjAw0VGNqxLrxXZcLbIuSo1qY7Frx
2kj5tY+lqNhRlFGgJUqHHu10PR/u7CGCza8qEQpbVNM4IjlieuoqI1nm617JL5aiMFgrjDPJVV7H
XhOvpGiOxDRxuWLFP6Ix5NZ2HLIxFegatfTQJUsiahdr5fbqcMZH5IUWw+/J8uQ27goFB3Fh2mhx
gNpV5htIJQ0JWqNDaBcZukBT3o1+ud9Z3qS/AB6h7SSht8uUxc5hC0ipNWGRaDeVcUViN3P1xAVB
8FuQFZtFgURGK5hFGTthWvtMzGFXZr1vxpSI9V7UTd5xis/J11X8naTvoBOfzIRwBvMsK07OC1Jx
/CkyTR5BlcFlwc/2mqDAK+fVLs9Q5An/jae6NZe4cfTjpmt5gpa2ZuAhsqBVcGYVv0dZ+e29WKV7
VhMfszt6loviBVt66sARF3PGd3QBLo60wa59dLmu998NgJpLVYkzHyIsanCN+t7m2VD1zz7ZkoDW
pL5lE68HOgvYnXBLg+kzEaW1hrJ7443rakm40DevdFDEq0eKWASwa2C5FTN6x6sXMjCq6Nnxw6B3
xAAzpf4sCADZVyyApagYcdFZGsKJOGOsAAmFtCI+ORmVspUu/Y2QZVJIFa7ZeeQXGZuWVsO+3Jri
d2A3CHWg8PDAK/afBvJqkEu8tdcqIrWd+T+8sk2b5kE0QAc4qYQY6MwQSWjwH3AVnUPb9g3PHhX1
ghml9b6JX31ncI5q6nCMQT4LHNFL+PH6ANKHGm6kmr0Tukcj37kzxgSJDQr/MeTDZnBQGJhQPlvv
8Ze1AteyTdCfB4E/IBhqxrKXhry+YyD4x+oMNl6Cze7DA1y0Fg+svgpNz/Dt9AUWMiu/9FUHAD0t
22vTB+o3bxs9oeJf/Kr97TUBrHw+hmmUql1TNme0xgMN6E93JvtKVZO0d5O1GIf1Ih7/J7BJIybM
WIEOpOrJGYbKDFBM4XFoUec5jwOVGtb7V9u6MZLpqVIL/d8wADHL4w6yo9NkXX/ePTuB1KttUjeJ
xCk+NF7WWwQO296tFJ4cYLxuESySqWVpY/tpKu7OOWNhQcwGXW8xXiiavpn9uXcC2uUmCaUbkhFa
jCTgyNX8IrnQm2ZK8aDSguwhvxDbgCVORh3eY5FOxgnLmP/wYu0gC4fUXCjCjCCJ0WSVlOyPuQ8R
SlgNDyEKYiUBK/5MDurytbexUhLsKLhQUTkDe/RXlCAtmSw3blwVQcZaEhDun/bAKFJJvUABC9dR
aUkUP6RFL5EwuKKtAUdzWMp0nNpEIiNYLhU8YWQatFyEnh7VzFQozhbfPm6svR3Z0ZL0i6HFlw8S
2hDS1vj5DG5kDMGT/wfQxpUXbP2Xqa5GAZvjovtmpBcsb3xDVt032C+WVzQAtmX8X6Ljynj2kuCd
jfVehDqFymFpIB4pm4RysxkzU/xfgTKMlxTv8fFRhgA9vcnqF8nz0Ck5T4rL/3DCUxuj+9SM61u9
z8p65f9NOIvJIZBLYtXBwX2fkI8it4BTWPp5VW/ojIyE2HT6cavDMOKqawyw5qxJPO9Ghbax17q+
T99x9zf6TfzM363pyjXy88wzcGExTv47ZUWdI27fVrsPfqBDqbTLv5h7dmHAuyJ44SHBAoMvJWPX
XMYBmPappFZOyFP8Bzyq/EzstVj6x9e89209pHlBD92BnCQk/59ZBYGaJ2fVjuRSHI0zLryUNvhg
IzWOWX+njyL5wZPERjQpleS4tsTb5Uuv9CjAgOG3lSupG0rnfM81/YnRMzlWgNW32ud/IEiLmF6L
lpGUJ1yWT2gVbEfml4jjAD+6zGpJOr/3+t7nGx3dRj31NjKMnVW7KAlSeKzDUKBoN1mjjHncNEYT
8OV24ekn5CtJ2C1sRgrvgSsddMUfjFEHXAtMcWYss3puD3hXRjUud81kBla9p87NnENSq+tiua58
roWMRAS8mfSz3gJegjt8/HfCUjmOi8FAWHK3coh3vRT4mkHzWCpTQkFe3Yxo94dHY1IbR8zlfbG2
NhJ5+xWLUX0w9ZnxdzKilIDASMIqewJChsJ+g36l3jR72tQ0tkLetgKyG/e/6BXwB76MjVQpF6a9
QHJ8Q/XnRscyL0Ixsy8pjSdxUNxEkDKBGtb8+gWR+oi0bghkCAJy2U81pJe74Qn67PFyJefjCY0V
DbcqqtbTNRUr/nbJmHiDjyoxARSGLGYedbkw0FtU9/jkoRqSfusJKSqGZU3uFV/V4/U0RgwOdmCT
KH75bb/SE05q/sUc0RivjmQoYCSxGAc9nKf0Of1Bgappa8hQqbixqAgrpuVMGmdKAdNrt4BuOzVd
qXaxPJOHt8f4KPmw9Hp/sXM0JHjP13OQBveM+Ugnu2isQO53cFWbv6eAodhx6wHf876zqpSS/lZo
ig47z8Vc3k4CGOwkCw2TfUdlyB/uMM9utAAJ3bCYn3jFYuvixTxzzdBAg4QzCbEIrXZHdjGAImeF
f+gLsaE04OUywHgBZYfucGsMffxDrdqepA8LcbwNNct4vDh6QFFX3SnIihefm1HDmgP7/kyWW/eE
Ew9EqStpq9Bboy7vtSZ9hs0lmHUEnivD5W/jpCkpq4P6tty0N+hGuhU7fb/7KMFh7SmGYMuhi5O6
88279T4xXImWhMAX06In8ue/TwaFAQ8mpIrHrvow293vlOayEPxjwC5akFV6WoQsBhkvfXzgZq0q
oK4f74jF48iWTagaEAVN23hU3atCY3BCRW5I/Nr1/Vmjk2HNSpod0h8J1WWpmbkABbb+5E7+g4QB
YsWh4pm4vOr1XtbP8chyceajKECNjnVXhSyXdH62QvEKp8TKephn2YSq/oPRy4xeBfNcnggr9Aki
UGPAk//qA+eJJZMksI4FhHTT2Ib3ZaElULHQC7K0avUfwci+75C3vIv6TSoQ52B4CbDURu2iT2Xo
SWYPbg0taDMX4SyPpgwr8aNQFR+peTC/7eljao9nWQUJV18uMVfi69Tda5LViDGJtI1ybScJQ1sZ
V/AdyG9Qd+USs1vEnZuGXCaUmSr6Jjg03OIgYyNp5y/9UvTGVpsGMFH9HsxRsP7bbk+xWMRtLU5l
ZkhIIX9b9EnnWeTzDIZpvPjiGhBYqNV6Y+ERaK2mJzfSFvO/WRC7WRigivQ3ZuhaElhMkowVg3f0
ZCfOQiYhLJ+L55RB0VUF9sLprWbjyne71TqVtxgQfgdh68Pl0Scyts4ujMVkvhz65ucQhmiaPGeU
Gl3KYAmif0HxSf47+dG2JCjr7MCoBu2xHYuZuBN1TZ5pNDtQr68sCercl2AZx4nZm9L6KuTj1uLu
1vJK8q9KHkKPQ/l0wGBtjAdO2vT+RL3UfQCDsiz3wzYtoA3sK4rr3tGTPhy517P/MJFHd5eYT+Hd
tVSaSxmVRSgTcGZWUuxEyroq5pJqRlBX9QFjJIxtCz6vkErAJXoeR1UiAU8M14g/ghPx46Qn2b/L
UZaAl/QREcuvD1TEvH1eu+/5HlapVcdCH5igStNRyyKArAP8zmdDMESXr3fXFcqjqmUDYiyhRYzk
TkDWhWBsEIYpAPoMF19alBf0LM7kZH2zIKQun3YzsIZZrh0nLCMIF1sHh2z5uA2VV7HfJHfnz9sI
M8irg9qpOQW0kfLEFbtJLWt5kHunDHK4IETfN3Knnyw+Zav8FaG/EkPYK429FJtgCKuytdRYv2oF
ygKvvQ+YSAh1oD05Q1HoaNN4grbOQtZXceGQD3EAh+Qq9cl29sWbCEGWEd+K0BkZEGFYzW+M9WW3
Iju+s90LhzqlaWWd7I88lHAHcvf9BwNziJd7/P4/DYrwRGQNAc3kias3ZwEGnWKczRvfwUC/+gnP
iJLjMN/0W+xhF75r/ILVmudyBthkCeCQSlT0VPw61BwHpQUU0r3JgumIcd0AMzwGkLCJseap6q0Q
T17EKEI8hy8ChcBkP9+ksDyRp7ovdFmylkb8PwhRuh1UZwV3aeFEZQcO648uxlbGHROsy3Akg4er
7LcxcKe2J4HnEQVeCXm9y1do3AswNhb7QUEmbxO/qpan4EV4FTGPZbwEIgpGJi92jXzzb0ton5On
fR3ftRow0HmmMGWzRg/4zDJC7uXCLfG2Txgr/r6nfjoi2cQDMx3Cf5guSXh25ia6WGEMjtLibnV0
TQgyNdfjI1DN6OE4imNVd1rMaQSpqFzdY42X7Fy0xrYo7rn+TPoSOdm8Jbm7UufqrXKdazjqKugZ
R9S9xvgKhAKb71jgnxr2rFngbXxYgYL5Igp50/EQc4LnbbpU2fb87LY1kJjsZy+VY6ZHj9vVGwfK
MkV8CEinjQ99FOb5Lw5diVCq7nn6s3THG0wAi9/tS78bwG2P1g/RAm0ZDxt0pH9Q0MN4I23NiXDr
F6QjL+LO6CUC+KRSzT/AKkQcP0YZxwWbvcFD97BdKw91n4Pjp8+S3R1AvPP5b+tK+jzqD5dXBk4d
5CQPwvnbEY1+PvtwlF4Ed/+35PMDA+yvmrTElkhB+H5cw0XDaa6fvbSYp5fVpQUncslaml1omsw7
hJaqtw28IlOPIEjhNppFFkku0ssZPrw0wTi8usWyZIqs1XrLz3yIwN5Mkml4V8C45THYXdGfkCDQ
JQNbkmB5rt8hzZeoFMOR0CwyGMsUtOLa38WSznil8unLXd+k+KgDNSJBfhgGGfM4Z5rpmrYZJzc+
Bre2nks/C5D9jR6ihfPBAOb0IF904hJBLzFhspkD6ZkdGWiZlKuaEe/qQ7g8rKr39ExoKCvfqU+L
+NmAfkDybPRfuMI7h4T5WlMApdaMVlAO4+zRCV688tfyY2+SzipgZUunmxuPdCnGIGthe5lqUpVf
0GQ078fVugrWqPuYu5emJcpSaDVPDuWG6fFak5mb2ZK3FqDfbXwJIzIUbJGtbN3YEjunSAnAhUDg
U4hz+kaqHL2ULa6REIpynBJ7yca77C4eCUeqJdUT8+4BN/b6GM4UOusGgWJuIsxKJX0iE49uAm7H
eqiPX8cdahFuyfVIcZqbzoOMuvOa+GdvnQtJskN/B6LAGhLTwBcaABXqkVDJaFog0BZWJjhVeR3r
eL/JvpiU4MtrOxBZcqZyBNkiG/DdTwyF73MP04O20vnseryQe0RtH9Dq5CocJeI5ME30K0kzfYpS
HLL9XxL2TVI3Gm/F8Y0iojpfBkcGDGLD7n+C5IC4Ae+vTg1h5R2V5hZqRJUK4DkjzIxufojFnvTR
YcyezZb45x5v8kl42nLS5CsBSuf587r9bcXBkMnGAdA88NEaaTOePwf2yN5ch29eTeBC7s8s+XGi
zQ8FrYqxmOpjE5BmM/c9u/KaGesyRcrvWF9RMZepcIcycWcBawguX5cJS2j1erwJ6VZw2NWqfKXU
np+IuSu5gVDUz8H5DpZbZfV4h/k9nTiDFFsc7q43syR9Zctz7tC/7Rs0YBeSw0uJdxQ5EaQ99eV4
IrCJC+q3eA0rRPDWMB7F2psmNlFDCcsEdQlCyXRyxcQ6U2Ate80ba69Oo4/FY/nghfWlm+3AeOkk
D/pIOJbVF8nzneRh4Uyf9oycIWsj1DeEj6zK2qcniZYC8KfhzJ03nEAQfRwbnm5BFYUjRbQfz4zf
runqwRxx9F9BmxfFAHaG2xumZG11Q03daMgQ+hhbN0Mw9dF/UzlzRKvYu2V5jWeBUiqoe63MjkGl
7uJIlpmDYAfC1E7Qyso9g+Pkj8Qy9Kag8x4FjhrLR4dTR4hlE07EtshtrtjE+tAkdCSDqJrYllNr
NgfiYbsk6CpgKf7Pe7Nr8TyjUpy8f4Vej7WiycYDgMrQ6YeTYYZBi604rGmdePdf2tM815dgyXkw
FG2b35ENQUHZSxUhrB/uQyLKTeEfXozqsdFX8V7pMHt+QV7IgwS2L+HiaqaxjuvmcwQOsKJfazFz
UXcOKFTyBsgHHbZfSNkFMGRfqeJVI2qbnxg6pas4lU6TfwDOugucQ5JVLDZdwS36Xsmpup6MY7Fu
ImaTdrDdNuicDacVrILDgpckmv/+JoCqAraovX/aO4qcU6vYPO8r/B7T+Rr3vevGY187nHXM4K1z
HRGxuYr5IgNjlwT1TzPBDLP4+Y04brPWiTIt3HNInW/X/YGu8m6Ia9J7CT4A7JzWvH3jYqUem9e7
rwVwWOE+pOxU8AIJ3P+t/KlR0wQwd8xhgO1tID7vx9nr2ARnFazr4orsn5BuDmaNsFQq5exb4Ivl
5I0I3UNEhXlEOpyopabj8dENxwu/UaQ4kIi4pPCj+txUV6X60JJaQg8ZIu3ulRfnjl6pqMfXS0E2
b2PLLLe3+GTeK9wiBWBkZGHXvAKrwxbNornWZtBLZPmi00/0fd8hzGKNH6lJas5u3tcvkLphnKDU
FkYC/kFRCMPX9LkWRGX/5Qt7E8ZY1DsWwxsdVsTjhfoOqeZVJ5DgwZ1RyARDMUAQ5TUW4JLY6B1I
ry3FwjNynMWMut+aSEXeowt+Q1Q/7wgkTtXuN6RCqZ4Yv2TjFMObxD0foj32UTmtDftyWI7uiq7r
fmm5NSwj8NamdPX/FeIIE2gQXRGtPNbIPxHSM5hyGrovugbx4hWGM+19Owa/Z+8aNmj+UJpGHoQ9
RmPjzX2IjP5Ky6ldGGnXZHKUfLHS0F39LSNITq2TjD1/B/ovYpPBW7fQHRf01ugW2yF/gKDYA5bN
oQcBh+bDvT/+AmgBPDrHX7VY7XOzCkBrZXacIrk/z+3q8czEky9KxejB6tbaUTcNnrXg5rkzbxkT
h8kYgIbGcCIO9xH+0upAZkmqDJJ4sD0cbyjmrFBYBH6okK+X+aTUJ0UzUnIkbOK2iDQgIkix7/FK
t5mCk05hb9WfShhmD9xUrMqNWaJ97Ws2Sf6NUtTUGzkxKUM4DhRmMJQ5FmyZ2XNjqflmmee7Yj+T
IjyAdwp1MdB13CB9ZnzMbmvueysdJcf/CgRtIJ5obLJnp6u9cB6m6EPmxu46LkIVSwrGtWL+berA
01grMj9rDGkIuvkbG6Y1LlbmrgbDQXiUJPlbi/v3hx/63EiZaufWI0SOz0Qyez7PtZXNGMFI9xvz
vRkDVgA6F+L6k6WGSCcD2aBV37r6vlf2XAewXDBRKtrpqUK+4pORi+ekFWUTMgYt+JQfjgGBae2b
sk0Fj8MejmOa4bev+g9rPvlIIkgC0gZ/V4mAfvr3ah2CrDQYQKXT7uW1d5byR43L7/P+/s1N98r3
NRfx13jmIJ7EjFS92w4PSO8QIZMiG49TwzhFQlE3u7SisFL/lazm7gUIPlP/iXNkiP5rMD7ZXxUv
WKAAf2IxCEoulAd9VcDnmoDySnezTiuOnbhEhYr7UJOR6kkQZdzZLwh4oC5btIEr8Kx8BN+UW9uQ
mhUfwwMjw+3r/Z2C5Pj1WvKCckoSp8C9jNAZ/PqjZjduXFEoxYeLkglQ4RvPk1VMUuxa0jF4I7DN
rhdzchrWPUaejGYJgIQLRA0gWG0sYKp1OuWsAD6V2mg5Cr/dThVBPnLA3D+i98bUIQ/UY5iKUU+Y
GO6jI5XqPVECJ5JhDlATXL51qmhCeWWS/sZ6FZ0W6w0Lmmh/5Vs1XSnUJYP7bg/SSazv6VvxuWU8
kPgPSOkImzgS0ktLC9nmrL5rNN+dYvFAjVIdrda9L1yXFZKaB2n9mRgz6ZDFARDgzYMXEbf1Ns2/
k1cIxabRBb97IEH2oNMz4XnUjPtqcKx8DrBgQRmSUK1kgbrI9lr+vZREBT3dyQXUG29rSSBah60j
jGqA9eY7H0OmZqlDp986MLXfcc/NFkps17NTejlNgOvHovZmhyT41jtDWB20LgVWMU39kl7uw12E
OHe1dopq5Z+TkkollyGc3RfJdITf5YEVhQuD5c39Qf6rkwjVR2ATyAZ/q+Tbl6Aa/mIXHMRthL20
pMtwJf/VWrFY96COTd0cpj9Qtv60hV4YVR/oUR+r4R5dxBq7p87w+8UWHp4OAAfY2empzwpzKy+d
/e+pHYS3AJg/Pw0MAP2VCIlePymDpZ0DvbFgVF4TAo1W0XmZ6gln/+FMFIND27+yt4bCLksvpI03
qEGmOp+Z/uGpZYdqDajL8KTtqEPx3ilkqTJ05bMxYi7U7SzClD+UrGSdDMgWCZU49M4Rlsd9qbxE
Y2t4A4RGTz6l/3UIFXQqhiNjdZgAsTKk9Q2sriNt+yz2Gthopbmg8u6pOegunGwf4kOa199nCxYS
F2Z9oh39zvYEYhnV27BezYxQ3jBQzdVUSD5szkNl32vZePvh89SFyTCSc6+3xas6LO3R0OV6+DPt
PM8VHyQK10VJoviR2jyUKIJDzG/ttbqCm3mcSwJvObJZKcQEh8jdVyDYrR9+s6xv53mpOncdC44/
uRmqlhBKKq3y+DK16ULO0MwrOiU61oIMLisFO/XCO3wBFSrr644SOU8a96ELSmL8dRh/A5PcIL+N
WD4UzJ4TWM3KXxG23H/FxqK1Lo508MlRYQS/ogW/rr6DuAP6nW53sysWQAB5z+4om2hqEQyTzHdh
H6r/5ajv5brixdAmnbYulBX2NGy/1mJdRkXkFcodtJXhduV1j0CbbliEp+dgqKatlj3UV81QmGrj
mGYs+i1TD7e1bzBpDKBn7UOxankL4nz74/uRkk130t/X62Y+Xw9ucMwJN2iQc4VRBK7jp/QEbZUQ
afcEgWyN8OhNqzKp4PBil/WUTJKcjksuRXDNTBBK9Lfon4seA+RiDtO3akfoFpqOThmiBXNcTOeN
HiJshM707is8+ulTcskCWz1+nHLoRnep9bt7urZUEfqgkNPbqM/w+OWI/7J9LUKGn/NxUhqitZLY
JbvQ50+ZwHzU8/cg7ArFjTNR8rzCJVBqFylWJRPwlTGsw4sQeyHuJPauWeMkBXmGoayC8qrWDsfB
YBgjR0CRBhJB2MKFmtvgJxq9haLG97xp+t5DxAaPXc63asyKMvj08dk86ZBA/LcW4NKRQlPTv9MH
trtw4zWAWFohz6zmyzWNIlBi149Fh3Bt4gwOxvUHhWk8grX8btHFQIbzMOpVw8+qXbWGKv2xveKw
H4wIbfy1LUPNnee1Ld6ntUXXsyMG2e/W/a+Rr01rH4pALg12wX5wA7kA5DZTWCcSMy/UQpgmT6Xe
ooyEVfS18KDo13pzdegLi02zsvw/XqEi78XS2M6jYZhVFNDZRF35tlTeU6VpgXKtLntwU3rXNUd9
De0cHM9tl40yM9DEW2FzLen37k+hB/DFKdwH/73a/OUi92adED8k+zqEtl52noba5cJxq1pYx9u4
kjp3cmCXKtoHnHDC2d+mNY4yBajcR7a5mpVQQ3Rn0hsGcALQYrek6n1pSujGZwMCXPrITNcLgLnl
qxEkmxSBFe1i8Y4VTzkPEgHNtTzF4hG9t9y3c3khKU1YWuMR2l4GIx3h0gDrNNLO5Ktwmp/5DvFb
wchxINIBzNhVs/B4Rvwt4Rd6qcaipd3c/kdjGH5a4LNDW8+sqBmbW4kNXRKex4BLdq5NvjXaVX6G
jcvdmXng/IJP9sFIYs72U5Qcyuy1mnhcqM2wPYxa1pZOvwjiwEyj/7Xcq8n8jl2HyhSuB39oKBvG
0rrZ2ykM+DVyfXVt5ahJtkvUMHHBN5XxXDHzQB+k+5MZLD37ay4zKNC0WtdbAtXI+IVPWywNYAo0
nUO9PC7rqanGKbRfXa6OeDpLvgQpRjDMY+2WKzWeOSvm+p7I5XKYJqXqdASCdtQBBVcXA/xGWzlL
rRg9fVRZ1bfEjXSgZbenNd8Z+Ef4Y7Olbp87KoCzaWZXG09KNkvt0PbKEvpUa4fiQImofNJLVOVX
cvK8fA1TTQMWimwSBJVTfULcay7NyWs36W9r2+zZ8YuLWfurTJSpDJRlDbpaI50IkWUvnDldpGEw
1AiT3NFghhAP2BbwBL//tsA1Mh4IL01PKJPGz2KhIbKP/OmioL4ES1Ei5NMDVDdu3nbjiWi1WoaK
iFNwHGFfOaJ/1MNsnHl0U2Adrr5ijzSMGYxdm5zgS+4y6iWqzNrH8ZMvMU/8bCT5JVasdcaGhIiO
gSyo0QlG9YOo940pAym5960D6lETgWJl4Ki+olH4HozpNDHKxmiQX+5etikCclQGpGgvq85a+FYI
Ix+L6QTkPpInjXATF1qFOtTf8KEX+qmXwc3fdU+l9qV6eDHflXc0PBIa6dRrVfpBbxylPP0pSDoq
Rd+UCO2nJboY0TySEyXhyulxjz6J83jEddluIDMqM3+wzBMyFLUKlrqFn5FMfuFx4a38pIQlaiTu
3Birbph8rv0QDpxG/PzEguWylkf9m1TPzXPlcXejoC+uNdJAn5EQCAxqYK6lFEWgh1jIfnZOsNFy
YmCQL3V90be88EBfu9LljtnNFT9ItKDVo6MWTOYne0tuPuqws2n/i+MEvFDFnF+YvlqjXmg5rx+5
dOkMdOvoKiaDWZ/38sB+3fxwaqJCGOykr0JiwvN+oAvtd1x2Kb14BMMV9T+ecE9aUOdFfzSn3Wfr
EKADAMfb+eLen6vccMk28wbtok/uDPjGb3QyG73+NCX13cVkIanmJwOtlLeJmYYaUSyHrn35wU75
KmuXqkA9NXSgEVIum/ymcXWT2TCHHZJMO0Ilva0GTfIW4K4dmmQbkZTbxBO5t8hMOwco1dkQvaPL
gpaMBeTgHf6LdkS59Tl9k+AA/qKUi2EGDMs/Zn4xC0MxOjDqPejTfUhqipq7GXkp4bgI2yxh9I7q
Ote4T7Y4eZKthU00R/Ft9UgkkNBZYv34cVI5Cy4LXygBL2uODHSAg+pDUHpK2cxQsPbxso4hzzMh
yiDJNjY9RYivHsXX8OTMIXN/pI2MfdxfK8tRRiA9+sQbbaHnAl2a3Wow6aaKwFlI/6Du110ifWlJ
YeJUX6vUbc+UHnro0bi3MsMqEwXECR99OfrXOQymK6unhfdPomtGjZsWuF2Iw3u7zCl2rSFBEKst
Jg+D0TuGHSWzG6ws3w3cqBjojpyvNXoXW/kX5w1dvnZYotWEEwl0zmIaFoq1svud3K+/YQFK0/BT
5qpK4QKc/ILeN12bUxlMbrgZz1Tc8m+epcKFJTkVPhkswcaLBIc5T3eIHZljp1dvs1zOId4+WOrV
Hxmm6yAiWW11YcYzICmZKSOJEZ6bKgHUWqIZ62leABU4lKNlc49aynVTKU50WNmt+WI1f1pQ+4qy
HnF+EZpW1YG9r6054fGBcPjJnkTqioEDEdGF3zwEFM+XoXm0yWCrWPrYG2VBiJEhvoj3fzHboSEp
ginlr2mtKPnZpx3rhJRMazWxv51DAFzDcH1j4UKwToafIXrE/yo0ND1j0r3gXJUIwxI5fI+H9HiE
w+axAFE6sdxBzMZslaWb0F7+x2qX0+Wi4RNTi0jKN8lSCUy5FNd3Tso0fmbrQa2mrfGaFDag8Sat
RfUlLPNIqZ+L8Fjgu6tWtZsO0SHzS+GxIFd7ljLT1TwiUjsa15lMRf89cs1ZuLJFXoUV63sOT98q
zaUxuOVu62XPT3GG/E9kK0/z14O+m21RHogd6JTvkOTvkDc2H6DBXW9rIrdw4EPoLaojb1oVndZv
i/8zrkvU7Xc76m4fpXB2CjdXUI5MC1Ko+PC+8sk9JE+4tyaKE8hWLK44N5o6P2aT7K2LHfYKuYwq
gMHxz+yNT5W+iSzp1QLU8vDsoGJoH6pLLugTTLOs/s5bPt+O3kH/Ukx4injlCF9RbfH0jAK4w59u
A1bKiMukderJx/d4wgdKCzWA9qrYPeUX5V9AmW9i6YbZibU3tOG19D31CeCZqI8hlUysx5CGyzcf
18TCKslpTHGKxovG2MQ50YF0NPkozcJtiA4sxKlm/v7HPZWvPMFD4bvaNzfN04r9IPkP7c0I9ouM
YTeVkhSWsJkEVdz8NmeFYsy+tD6itnCSX/icqvoQiTbuzIzW9o6YBh17BzGAnOaLdB5Zqcve6rRn
jqPv4QZbtF0xPFlkG84vSWRc6xi2NdkfWcKcAwdLTN1Kv599Y39AYQLqhQGsOuR3Bsyjb0T96hxg
blhQ/U00HhH0NXVVs5DZsdRm5ljb8Oz+DeF12dqiY/mRwut+c0weYcOkPUReWRsHzxpV0q/iyuVN
17a1FJwBORJsU3j1bXJqJfLfZgbZGcdwaZd1xUwFdSQxfwmCdzeFG8D3yKYXPoa7VbgIxU1GLsy8
ud731pHNRuM9WT0Pu/Vz5F7oDhqci+8/lvoE7IOA7grCo+NNX2aOnjSRxOjivI8ZoOld2tnd76i4
iGT5T83VAvqfo+cEkjExI6okDwT3Y7Ej6/YD9W811nR0duzWg54DMT9tz8h+Zg7Ncu5NVOpJlF+p
P/ykTX3+itWHiAV1R80ZiXBEYoJX94fYOy7xPdyWjg0SjU2vCNTGi5AtIGG1xyxyWrCqlENwvCAJ
DKgaBPVe3nOgtJF9Pz4DEgg2cuslcySZPnPP72m1cMvkYs7yWxsYaSENp4QEuGqhzb3qw1hdBRhH
OWvI5tgbZMtKVjTfi2hB+6qAOfPPZ88D4S0Biv5V7a46x5CDjAEf2krGa+dtOITokIdiFCRzeOM4
nahc88Rs+YTSa1/yklJ2a51kTwoPZr6tseIXRRVOoaXffPT2JNVPkEcDGTRMMYugSL3PyEWKjIsT
5GCIHPbpxVCUkofB2qDRDSKOKFwoHpMleQl0/QzEs6RLAesH4X4uyvnz7AtOSlPXZFfzih0fSTHj
DRoj787DB22ivNCkussNVVk3XlE5B9A3h2l7dYW0Qre9qkriDJ21uAFHn+WauPIrkvCBhNBfVBu3
raAjBbEeaOEGckjBYsNWpfOTEs6yJANo2vZ5fS/e5eT84xxi4m6q+d1MKEetu72zmJtRb4DoL8Uu
UVxEGUEpl5MqayaZhbBKzEuUiZy17EwDZ+0Pzbhv6JgZz0lEnMLrOh822aWO94oBsILIiyPMAOyb
rRg9l08ILNs7aLAhpZ7t/iROP+7I0avTV6sDv8SguWeAWotakTYHNf3RhoMwDoJ9I8pNVsndErGp
s+BFmgnD9scJ5ooim8qO20isxRUvVh5qLnP9JC0Za12rqOGHczKZ3hbQqrFTX996DoCTeEzsaFzk
vmNCDbiTueXME7hMHOQEZdzUbCXqyiFWt5X9/9ZKrZvCS0yJ2zST9IIEPpWjQ7BX0BdGw6MJVvvm
OutP7PM9b/7zLz2+8lSgImbWI9NTP/Ua0bboiHjM9dssIgAYjmTpmL1VmUW3dyzwN0rp4AXPKq4p
JL3RbOICYd+oIGvvukvZmV1AMRDlZk6MxKoh9d8u/o51ZdDkRrVQYM4S9RS+t29O9EjKQHvvU7x9
nS2MIohVd8RzTDXjdRk2n0euk/IZcktjwHii6GWSeNCOaqepXn7aSzamKnG3H1/Y4LryZeycy3JG
JMBGQn6Hfr+DpRzS4ge7rHAtZp0V4AdneUj05eDt9gp3rkOVu+sXuUeET3H6p/gA2U331B/UZlBP
eqH3m5bccJFRW621zaRdb2Rhv+VuqyQuIvx68p0s95iY0K0Sid/FZpXnkaNWtP+7lUma+S9u9VVA
lRFoV0/GnK888/A7My8nx6tAuoa/MOHPLC38XoU2DrNYFNmWBhLIcpPhKLlqHjDssZFi1A7FiURb
K8zJuabfizlNy3gRSfzn/WuPVJgCuOf4JzgdHBI/67S0NEF8B9BV0IQY6BsGCkYIq3qfns+EBuyG
bo39lemwP5ctROl8MKY/ki8iYQUEbu6LH9KHWeNu9ir/nNBRdAoCdUBc6e4gEqOINXBVG2oywrn/
3SzIBcxjaF8drcD7HsyhH6h82jRXq5VWwekfYkpSC+VEpZGQaq0fbtQrIpkPO1U91K14NJP/wTjL
ne4sMXsCTH8i6aCSy4y4TRiucspApJK2hAE5uMdVenchIa726P/eLaBIyKusp14sGzQGHhFfFGE4
u7xuUHMHfBn03juqjprFz/C4nviaV7tO2WdBu2Oeeo/4UQOFckSG0D03pv9iAs0NfZUL4ciy0F1j
bf7oyl0ELrznBa0Nar0wsvySujC5aJ5W+UERS7zUvsApSz7NBWoKjq0CqgPZC1XWYOyLEhGUAjxm
NRtYMXN6FiPXzNK8GXLJTU2S3IrQhXW/HP/7+UVJ7x38n3Ib3iRIptu7xupdDTn5hHA8tvpkh1VN
64RtEzVTgjFXX+KHdDHHNNn61XNZFQcCRSSOPWb6gNUbqgI1nXBUX/LwRfIeT3jszmejVV10Iac+
kR/w6iD3ZPW7UKsG1GXhT33Rn5iA9UjQBAB3/XVOQIlUkY5xvMg+0WlYvnDrjCJqZfIBQi7M24St
g1aDiM+V2sZ46r5fjOWwEalfzXs6ZJzKSQnCYoCtAwOBa2l3TJyRVRhdoAqOfOmBiw/D3v74xalU
+K/sB9WEvunWNp4Ld1ltG/WP40ZCd4iTLcOSZTn2ZFwo96cWmynkAtLHOSpnQGkCISKry6HlH9VG
GvlYkE2IJNQFGgbrlfUwCz5QujI+AV+Sc2kV3yeYHAyK62DI9G4MhCGJVZCpgoVOW8h6xLmvDMCG
KkknalGDaUYFFVZrWE5Tpm/8pRYUQY+to/a+mA0dyQZkA4tot3QaEWnXMPjfnHDWGalgmr9QrBpH
99ICAVL82zkHjsfzGkZIPAbShlUVLwDFYhdJ1qHiVFuG4vS4RMCnTLhPIMcNVVJaffpJqSJNdJJ/
/h+G23JMfgdSMe1G3dgRdQBU5TszC01GnUn79UzP/Mz29r0rlTAcT1ncZTI7T6KD1qspnxHrCmRe
SoOdr1KiDkxCbZ6JeCifGRhOBkj/UE0FRaQq21nBahsLegEJzYnlJ+hjAL7Qatzk1FfR9y0dm8mj
RkX3fn/kMKctqfmt3QD4G/MBdiWJPBbEcj67Srb0lCTw/8Zb5gnneSS8Q4/T/+Lwl8m8Y/geKt6B
Oa39BMNW22cYMerIlynlEQoiVfPkF1goFZjuQrqRdqqDxs0cWOFv6yXLe5gc4BivUBjtcUbXfeZl
csEqedS2xI4AfHqrcI86rHLNTLSlXW+jZwCIEONWx+RWDt22kWCfyX2l92jNxgRYC0JAJbLp1tf9
UIP3qAbVkNSFUzRtofhldyx3O3quQyadFIChNc6tEPFqbPmTGIR00aUOTkq1cVuLI4hijMPSK+A7
lFP9IF9bAFzCAx6vIZ22PZVP+t+hAqaEXt5HsE3SY2MiPVoS0i4sGDur92JfpqqqhW9sAMSBaOGf
a0CkeuOQfM5a6PBLdHtGUehY2HnICKvTsjlBUKlhdBgRSXQQ6hNo2lZPuyjHrTR78iiBsrsSjQ5s
i7z+mrbAKkzIcwV/RPKszDm8J23mA3Xyprkvd6Ptikki0DKdbE9Vv2RXA9pFpzTt35X71yUoZ9bb
KIJjVjyFWfXFIobo+maxsmk2/QyVv8UsuO83m0eld7k9t6nldUjv03YgbVgwIjZT6W26M1InVnXm
YbESyXhLOYbwGx3n4Homty8t9Wn99511378X7spreVEUUpkkFqXaIiJH3R5bPByVxv67rRZ74Eci
gPSX68WfLr2rWxQjKSgaDnFQrXJNtdKUV4JFXB7r4i4nGIJuYz8atO8fKOIunQ8n/pFdOTfBay4A
o4jY7X7JyFA6M1y4AdQVRAqBiTw3MsSOps7iIqr3qRxlKznL7Ovc63pJsXGJIm1cbGZevBY7Gak9
GMNSnupAPLPAXtDOYs4desVs3epIUgNkFa/KZZJCPAJm2hWomZsCe8bBl0aeD1zvzgVy8r9PulCC
KDPVcQtHkYMeXP1weucmZBrUt1F/mEL97Kv0r/NeSAKiJHCwnJ3iUU23bWISDvuiwFZp7OBZoTb/
0pS6oOakNAZ3iZ8ATgn3Ay1vDNSru0U8mc6irJzHF4F63UYS5Ke++jrbAMX0toCyvWsJHJwwXbak
/BubNcrd8/J4A02xhlITgM7X2iSF6SHZKQty8fP1hjLfSYmdtPnE6+/n93D5h3qNM06YYOwOQiwT
P7bSNQeKwTbBBAd942AHryx2mLVs2UlgTZQk9rcrOMDDifLFqg+g2tcBN14OPFMl6YUEzN5a7aJ+
s9h7wkiv+3ARjHArSbM1NFSBIkeA0rXn/fSWqcDhc+WXZYh2Ptqz+5JkQR0nFvGj4t5OvqTjH0a6
i/uBmPpwM4OUBRFlgBF8kQsgT5yHDc1e6q1ruUWopdCX3/Jz1FkpkoEvMADphaxYj+QEu6hYN19p
m/3zV4wrs52t5sWaRBo5hkEmyTs9zv+vhtYBG4daYxUSDXxY8iudwTuClSxPhlPqmD71iEIBbyhZ
Ab/HIC1Ug2Q5XCXc8dwnQL5lw6h3n/EuJvZB6AURpig/6Hvcl8cp5xhCr9GdU6kYX+oM4NvaZdCV
1psP8EUZLJhd2bkSPgCNo558UdNl1p0UDJsMz+MLqqJaxV037AH5hocXa4zJnLCwaGO2DiAiYyfp
IaPyamP8wbYTONswJ/yQEdxNT+GTwKs7RC3OSYdw37OuGwIOhmvuYJzFERlMf7AJ1LMWgG9TnkPm
GaGChv3eNH2BOy2LPQNjzfGYb5Qc/WcBAKP2F0TCdkHuqOKzAHc3B2BhVUZ6eNv39908f9ZoyN+W
RxQJCmt4Uq/bwPSNBPAm+gaIxZz0sKd2d7ufmFA8FpG8AooO2YEfiPxLsqDkKnLLoYQRdJU5dmxd
2MZBHf1Nia2thHIBIHDxSQUYCX0MtoakXvcFp1XyVXglZxLayDHSvqrKxKsPVRvPDrx8d4wbI0Tf
yfFshKBBBXZnQ71SJTGQ/4GwPNES7rooZVYbEH6bRAGS7g08j2yzKFcQJ8YkNR6THyJcMTKV8zr5
rMPbjBpuqn4l+ET5YMIaPUFUgXQbwHUyYhTwvZjeX2fkFWRmxEctKlVTnkAC+PMF68zzZYZjHdla
zmPHYQXHd5wGzyktbb/0s9gZ0tFZDu5duKsgiL6um3ar8WobFKGLXu7/AiB+2EtUuHMHWlWLcrLv
5DuhLJ4LVMhAI7IzquyRzVYonjh6215hUvjDT1XNFYTPCtwURG77FmprDJt1dQN8QC+fUH42dz8s
Oj85MyMkguP91ihrKkxs4cS4UNXV/3/edn+HtD20aJNIL00TBCgoE5IbXYIw21gocDmx6Diloc9h
c/A2omIuAt/sNG4QM6rrEBurYzW3ep8UjiNbJfoiLkkzjPKjO1r8+zAxL6UZj5yJuPpq4F+2DPUt
ATGItsi9ju/7yT1qMw2CAK6igVN2tzfN21kkzqDhlaMWQPz87r2xdLZFCwzpr5BL7QvrCExq5284
jZgQsVsQkXHmrbNIrpQXA9p/NnYTcQZkCw0vEyjx2LhwIsl+7m05QeSegSGcmYOZBIcHVs8x4mGu
AfUff+MRZHiBN7UZ7j791xD6HunZXG3idsf8jt4dxK6UfYh9rstchEPjrqLnOYMFxYn1Q+HJYmD9
PCSpBmSQKGX2rX/Ti/R0a0zpzp/hND1ISQB9NbneuwXm3YhFbIiCOLTaOzepKWR744dpF8nHVicK
xp847P50fkGHVc+vTvTwXsOZrO1kcDWdLwTr8rWfldGPIpmONtbLjFA4oAR+JJFCx/j8haPjeCXO
qvYYrPeHIkzzc9MLbOGHzq7c8ElBn9E12mrhj1lfuoKxn5uzxd0XgnB0fq4CROXSGF1mdzxR6kug
9UKq9mAghdNh/lTVHaiWAZHE7um24HlpJyWj+5ccQKx14C2Xy1HgJDsvgqJcfxCp++xyzcMwqmxG
mQU7iJoyiCYQtYwt1XpYk/sdmvdhi3NByyuOPdeelALenOPL+BYvHaUwMJNiXYX18vXDwDn0/UMm
5BSIa4OPOaEcXspirHqynvmDHpEw4Fn76AkBjmA/SPlC02ew16btpIVpTlz1IypvDypIsNXVep6m
yUWdnWt4efjgEnOSzY41btxL8v7e7RNpxfjvok2JnkAbB96SaCQ5QD2+Jordh+lVrugu610ECPic
Ty3xbB1rywppJWwDiW5xODUFrsyidRvzrwJ+A0MgitVbQeBqQZjMB0NH8FNma+pWYoEyG98g+iuh
p8lHnXuaKpetFCiRZ0mD/m/b5GjlmVDy1VEzqIsBnptuY/ocNDS0TnleOw69nJdprd+tx/OwnVbb
0KPBK6WLQe501YqeNXv3WgkT22HgNvUWmbvY4CylzboH4/svYPHGbHU6Ip0YEVM/B8L4WgQ76XfC
bTteJUlyddmuZPUb7uwZc7L/AaaZoc63pkFTPIdjocuBbNmj3zljNb+F2g/h5W4qqqthY5nrs9Ll
xqeO8+KZDFR/Dh5OIJ0mEj+0D2ir5idtzvg5bKgdXBPCAEDjgGvy0jljso1chfeD/xQKDQBHZ0ze
wh4KMeLUuY4DX1q+MaGbLpPkwO39h80BKnUvYpwA2KUJQGQ0odU9/yEgEQzAdzCJQgx7tf7A9oZf
8uePhk3O0/+36UejdV9dRYYPZgNf+ubwY645SkmAHBtqpNPGWGhawmM6QgKcPrOcg9quQH8aZVRp
HCGGitAS0Mj2K64F1ONllD3n9C8vjJoUxjnNOe4CBlm2v4M9tI4u9MLaLc69ScEeaaDjFcOoIMoh
x4hWrqnYb2gqVt0oS3NmrEACl68kwNmtal8Jzx+xWCxV5Gna2JL/ikIqrFOQJ6+rK7DZuWW+YRc/
TFgMhT98AGBVO3FoB0k3+CnS7hLZL+VCe0QiCQVCdufmZeOulS51ZBFIzcUgTL0MEpZdOp+y+cqL
ljPgT78S+yFLbCQvlHavyVwKKH6psRhQq7ymhSeir8QrfpWmYvDRLxugQAqzXZNymKXiz6ATA/Bj
1/7ofT3KQxZq3zumawfBz9aNQHfJkHsDly+kUZwRuWLRQ1xJlo/kmFZNaVYO4EKBx8Hn8CJJfZ04
Z3hy0AEDIAnUTAaG5xSFf3QwDvwlrDZBIo7qHOgG48LLoYCNi26b15AaXyiUr8XsEScu7lckt3yv
Vpu805rf+i5T4BDqP7v9yEyoRGKmkUWRh2wGEF0/rJX44jWouQIATl7w9HtIj6sdplB4+nbkTvXT
2BKvhXZNIuSYbNjiBExLRAq69E8FtdKKXvPNLk/zCxZKwXM0tsPNytJzTkexzoQyIS6ONue1uGEp
7243WDETfqXCo9dVCW3qkxswhqjI1EVPOz/kUDxFNbKIGhwVyBivnCEQrYftVmAIN2IuqoDtbZ34
bob7LATrwi5uYGZcYuYYy6eVzFbBWwDCzliOGUhKPT3KVndONmiW12IvNRgleT0v7ifytBKZqF/V
JvmtRqss9Jgcp+2c8AQbTg82LH/NBWk9YNpwUa7f+DbNoRixAgdLSBpp74Dgw2T/f2bqySAIKpaf
85zSITV+GWIBn2v28TMRDTDCXBcPbLUa8x7+oxypRl1bnAw4Lu7iSw1OqQ44WF5eMMni4kwRd8dk
e3x/THWPXQfKsQpK33keo/bY8dF56D/F9vAzXI1UP2B947sow05YyJqBkCPC++u37uFA8xzliOuY
iTvAlcM1/AilDXcPRHlhaMdMx/SQtk6PrY/505ZykdFbK4nZWthmGNHFauxVW7qjQ/GViLUlQ8dM
YZF9Z3gNC+I4xumOdlT9Q46ST+b22PVjYMGLwn0vnE95AyhzgNimKrZ4YrnsmFe/61dSCNm3nuL+
QGqQOeQHJWOUdaUGVysRsCD8xhQbrc63jrojtD/NzT0epZxwWj8z6HDSX5MZT8NF9mnm0s/k/wEp
kp4SgtJIBVtDVE27WX9WmLuvUql7XDVTFD95LlVXRjymHYWpFPMo1fn65LxHf1ndBSLtxnmERN88
LiwTBCifYi2Lm2r2vwiLRvg/b7taANJpQsFvXgoKNKbP3WXw0Evao/9Co086pxIv0mwgNZL7qUJg
PRTEbmMtx8c5AWKHSIFtjEBlVs4PhJjWxzx/dDaXiwBQUUhnn9Qx71onVywlFb8hWc9Lz+3jiFoW
MppEDW3GQJCyPzlJGvUBufhZc8BWpFE7XAB8qG/47uIq5K6AeTGigCx1rjd4ZoVUYNf+QUnjNaBh
RrCotO2QG3R3vrkGGwuFUMfxvq703Oluw2MLgAVICwMvuzXP+8r1m4l02cWRB6ARAgph3lAwehqH
53iGuVQ7/+WXJJ8EXc6MpZX1cgh1aGV5E4Y+SWoLCQ6IEnyQaskJ/tdLtgf9zSfnimIymPk+u9G9
JDoc25AhrCP3c9/ZFa7BCsNYEsjCS0tOK/joi+stbc5/xX28xV14iiDDewT8/59Pk2FvKxE/tZBy
4Cnwln7YelWMhsSDhDCEyrMuc+mhK9SMaEuPwV+OOmwdv26Po7iOMUE/+VPXDC2SPv4d3brxJ3OH
QZabcfYGOZlIikR+TF6/biU5WxYwYCKtfObMidYZpdzVxmODcGheORRNLtGFwHAJVH88F6kG1m98
/yBVmiNls0X49g7iPbNWh4JWKyoL9P+pXdWnXF4I7KEEpWdpo1Y7RnTu09j0wb3dMoNJB0c5eHak
eQEd6jrspc9rDnxdVTJ0IsyzDS7kttOCPo0zog8qkR1kXyLY7zKYSnw3DkxxTC6FPr8QJTL/EleN
6PV5sgg4M8U5V+YQyHoi4e401K7owTuHqcPppDCaj3ssYjtesNGN3R+iu4ymgK3KPJvYjMTdTsdM
fYr41Aqz3XTi5SJuDojaJul2HB85ePU6a6LxmlpC/ihnTrsJPh9cHDQHwFGxpaiZADuVPtybFo2s
ULON8Mkh8D1iFLHLk9SLhofm/i1IyrCOA7z91CC3c8rrc8+Vj+k/JkBV6G8yII1NOtYmMBKU4nIu
+3qx/z+aZJv+veZCom2bkJhA3ZvNiD3eeD5qrgVhrIY+XtMqV8NhDpjgIac9wAkikH7pZl/spga/
kD6OI/XsL918SzHwTOKwlL9eILB+2XPfe7xBa3RIIUou/QnE5Wv0RnkXKBuUFxQee/jM+YY8qfFu
kTLI6vd3+S1IRSJFsGQHoa2k5zqw/XfABh2kyrUAgJ2KjRk/VV7hWhqxZASqSQDscXdNKSQSo8TU
3GoHdNdZohxR1C+viFIBjlwKFTWsbncwt3K0JiVHSfYm/vKMYQ820hp/in7z7KqugFpw1OEyvYox
fIeZjy1YsNPLL13I3Q+TscFitj38V8HbWjNQ5W8PJo0nP1rcGPQRbYr+/gd8Hr8BiDOAUPTU8erO
7V7nfl4Mqn4+/nwEo883nQ2BLv6pwFP80ps0H/gc5tnRCRhgW89LoK82Pb3cDxUA8hgDZ9cO3i9h
NZVQkXrK4KwjS2J8LmHNMg7aqnXRZI/b2T57ZeJTyQGUODOQyKUKOIciOJlhnhn3L3Emxo0/VWqP
vmlvxgIX50hcdAj0U+51sWn9N0KzaJFRtlsjV4edWsD7u0Hfw/8im8vC5XpQkGVwW9OZLtwIep/K
HK4XwaQj0WPdftN83SaJJZuECxD4Iir664pIBuboOqH3nrL325W2iUwRpHgAP28oAbILuSfG6QUk
B84BL6MHOVMwDwqOFpYu1WNv8oxNY4jqCNUkUSwteNVNxVUitMAD3ub3vKlvVsCuv/NGYvU1Qlvu
XBn97jrFAd3Hif8qdVhfgLuDWTMiLCSqfIJGJCEfJ4tibTP/cj26kIR6OX22Q2wX+qLsxloLDuN+
TXl5aO4y4fNJGb3e2SU9R18tykYjGq4NdRii6gFsm62058Qwb/ubmo0zoZTENWbP2J7BYjGozAYM
d4Efw3oPIXFVVqEZd9H+v1xfQ2O5RJivbxd4eD+B/rZ51VhR6mHrGJJ/dQhyYjeOJvyI621zQvOz
B/7C6GogCNS5KgcKNCAC42yqo+Btcel3KYMlaNR4oihPEP10EQeTjrC2dJuSPtQxJ6A12rmtyWVC
Ccpl4aRQx1yEnik2146ftokUKTDtP5lbFr2YHjlhstpdfbZWqOF59n4Sfhil8vHkXaje6/vRCRPW
jgVbOYRivlsHRhmjJXgy1/B0GmaMVMDEKjZjFNLnO7UFs6ao1oSMpUWoyeCQj+JUZmrhRiVIf+GG
Ltbez4vllfmVznCHV+PchgMjw/2bDNctOi0kelenGxB8ifhlmYsxGkUuRMB3PzvozL4vkOAJoG5N
16LX4097pl80XpCzllo0UDpdBEkOYE1+WwFArKYy9zvg+n68h3Plb+nP5mTUoHoRo7+fY4MrNN2R
2tL1G/63z7DKLTim4GsnxhzoQPWTk4/+bhTrHEWwInR0p7UiR+HW4FEwuAgxZQIE/69UPh726EIg
SKnH2Vq7BDLinN533nT2eNzz95nXWfCghfvlqwi3k7prJ6eaN1r3kPcOt+jHUulfIEiLNJlpcEn/
R7mSPnP7AijjWi3cSFOLNT9/IyJch5cxAlgdrFJ46atMDvKi3e3CHu0LhJFdHVzzHRZ/Zg0dtDgM
Xw/ZJyIbJDXm8L+STe2nl86udgyiMSAvgDK2OxGXijGSqBb8u1TWVs+3qUHqmSQKQ8tZtIvWkcP1
DWII/tJoqKIic+Boxwi86VXB1Du4jnMLVWCfT0zDgD3cM4Ao3AxlNxIimDEBFq2hfI9lYlnlW1IM
uqq5oDpQSHKOM8OLnVmXHgIqYR/ZFaBHSDsOdUwLCh63Sbu7P1Ig3v0yCbyPYOw3YanKKamk5jGR
tbdtca6imQnTlN1Fj+EYNTkVq5n9nH2n5PhUThc5rZLpuxjLr8KipxSiqALp98dvSkI7OMDin2Hc
8J4Oi/CFJ2MgPUXCa0J5NDn+vVVE+THqfIYu528EqrA+tMmuCb3wI2nhQQcaflQoIYjYJE9pGWfm
/X0/dy90GndG3CbBvYPEuHw74vhXfaqpWnIwd6CkPkYWzcdtPyXCgig0CfLVDtO81/Vbb7v0SDmf
k6/S7C4bQARN2uAfP1wbEmc7BRMbPAKuVoXAQUVea2qNbTtzjZ2MSv5JdFxgWpogEIOmfreB36XL
FHfrSqJMpMetlngzVclF/U/mrCnQfdv1LIV+x4JVFJ9SMLeWlYfZgmBeYO9zZ0Dbh4mvI7CepANV
ryzpZkABA9R4js41WXe8YgvDaT7NN3UYNDEAxWCMaFslQFbE+4svYSREKn1hvbuLkwyis03zVkg2
KCW0YUsYc1hnR9X+eG1W4/GHSNcgr0mQM6jeSCiIkFzSDy8bESz/6kOd60J0u0w/+5PzgSr/TWkn
Z3vxG1eP7UDXJQJpPFHyLtdwo0wmMJS2zVrUUt9l9u/q1tRTm446zXfq9iwIpAX9If3APoUSzjgV
XBFS2ZvccfQxkAA3ITpH8rKBlv+FPrO811voghYGkDyGmKYby0BWj9/M0nDsjMQwXYvnkxq6ddJp
UdYx6wnL8Gm3wjjWK4PtBXnaYcFtjhbelQY9w0IKQky8hC+oiZquZMja2gfOpZNMC60X7Vgdemf9
5KVU/Z4a1Byd7XZ6UD1iD2zPP3ln1b56/QwITNYXYsiAafTCMUAQhDGAMoSACO4onc0n5colfAZb
vjwcGTHnLcoq2J5VouTNr9zHdZ3JC0BJKM8Tn3/lNdBP9k8QKeS3hoO2QROkiVPuQQAZd+2CFkmh
xallN+iWB0szjdF27SmAnfN28m3vzcT2HjYmaCiubd3YQtvQ04V33NxBaIT2W90U1+EEMn23ssFW
4XrT6hxthhxl0VXqCbLe2qasdL3m5xqD0NHRQfHzUkiKmaBOI5UD8nGwn8+UrEGR04BKyzPSzEZQ
++GxYa8WkURMHIF4vg4+qQ/l3twV7+MCSOOmfBwv/W5LkwEwhOVc11xI4MlHwT7UxBzG2YrKx/TG
F7Z8qY54iBemw4b8z98o89QRhLGW/Vng9SvTcDe7zOlYLulzRnxNwkB7vAT8abUdVsCIh3bTZf4G
u/BztVlkZ8rNPPHOu72IGs/T0LKTXSJdPHhZ0glFJMDnunGXlV/B8QQet7w/y05/zQExJm4yuyAL
oy93GbVkZW32AXYmsl7PriJVoV9c+cErMZ+GsjZfQpFsuYK8Wtb9a7fVnwdRCWv2DlC4SAtlhU/5
bfTYsTMcfiuA3qvsVF7++oTPvsU1jlTWKcXT2Yr/yPbvxaoEiNkWe9WONXJa4sGVd4iQrDXfz2E6
RYOw9E8IVaVmjIlJ3IvROFcVSvCslfoLxaNRV9Co+7ZYWscW4lrpekMywXB/SYLSfvS7xIGuuTpz
A29R+X9aaNVvjWNl+E+GQUT1VO/RDxmd3Fr81nWXyFuNONwqC9MS2U8fZqznoLuEkJIQx11X9/Iq
aPMPrRIevsA64DwW6u1x+k+H42EDbOGQK0jSaaKE+zY8cxYzU+YDFxnDpgp0m4uwBQ+qg/cWZCvX
nweHpG+XPexyKsO75s70/OBgf+Eb61sJvigEpn4cavu/B5j/4V7EnVCW6lQxAPGUCpDkm9+2uOWg
lF8dev4a7Y+FjatVOX3jbbngDmpmxwCFSuwuF9pOn6oHfMe1AkeaiYOVUl4mkHjMXEIYBm7LemcM
6zZw3qfKGKvenLUnzQe2bXy08cSCXosA+7m83XD4ZuLc6sGrNRvRBycOPFJ+F4LdpgptwM5kNaZR
5pgLnyx3xlrkl8XWXB27j/XWJHHw/Wr8TlTKfCy5F7bULJVJRB0wQb52hM9pAxE7eiLS7O+JRs5G
MZ4iAh9uSrQJhqHeHRcvVzJ1OqrlcZGG4Sn8lMugdsEZM4xHZZUsK2rHJxWCtGD6FMukdC57zWEn
qydHG4vVxpTSF8Bab/cO+gX7QndkhDqMafx5vfQho0MU3c9AyKYD4QTnb93oNJprTsTzRn+Btaxk
BCisBC/NiHom3pCEr7D5P9rvNp/WC/us2WlZ1WctGdxpDK+0TrwaykA7Ah0pJX4eeXCi2dZ16i3Y
jdeNNbnY788V/qCPTMd0x/fpf4/j+aITAZvMedpmkddRVSG0qZwo24DpQflGXC4wzAW3dqcNa5vJ
qDezEY5TxOK3vnsRCtRDSqwQDCqFBex9Q5NsDcOB0NpX+Em1/aRlzct9qiIo2d1Ko+RZGok+LVl6
p10WE9j9T09Weq++H0Io6Ha6Ds2DKx38lhJ9MujahVwEf8ZSz7FDl0Q1FnyaBnvH06T23ncTiYp4
s76+3PIQexaHP3q99DNEEP0rbRXKNc5P/DvTb4CoJglgFmdt6kz7iQaVU7eGGzeIEXJbVsKaIMlX
oqE9yIbLoGpX62Um3qDVTv0nexWyMAHgQ4uJ5l2zUgGTIAyw3s7fOmHr7lGF3sbYdBEXFCC74qu4
iEHQwokBb0oAnZT+cdASuCssfCHAhQy/zNNyUqtGV/oAJjcNrQ1sweszSnWgPWMTwW1PnYnGO2ev
4DV5MHb4j6q7vtnnUu313xAjAvLvFvdtfcvGB8izVlnCpXllvgs4cOnl68OHBAIBROkEvmXtwULR
YyhIEe77lCYb+dMDUGES5h8Sg6plcOKmqlr6dkuy3NzaldsDgDZfretqZqjJDV1uHHXY8cG8t2kH
nCWXFvwGQm+hV0Zt2/n6Qls86bTer+P9S3ob+bSoHfhnMQd12aQv5dZpOe3GMZGrAwdIPhcm6K0t
PWbysZw+WyPsBdqKnK0mjLsEK6V7Rg6VUK46T5FjKIPWEl9KJSZAkog+SK381s7gZfktlhaqV1Jm
eiV7WvPnXy3b62xh+P/WLQ7IppJGGM7+rXM5lI2C4XvJaBI5z4BlrUMenmmioDmFKXcXqJ1oeM8j
vbgcHDXZwpH4K3adnpCCxAkj4XvNn+X0texGH+E+1bCCHnE1M7l+SUQuVcmR8mxYxe/NdfrjjfcT
L9zn2VAwftg4aItmsv1GAXEU5mwN7964ybD92tLuvNQqZNaVqFBAFc+CHxiKUH1S+txz3rnojvzb
735lGJsXwVdnHLz/AomevDwG7FeLWF76qdL2NiJ1tuziKd1fjeqcD1WILNN0Wy5XajQ8S/uo2+rm
PZlGRrbWnWxUwHD0ILIJEpdtH7mwtzYr6I0EsCLvUIFFi8A3u34Z4ohLVrgEh7zD08xYW5HSI5Kp
eqpu+syu6mRnujQa+cQdYxvSH4I0MZ6FDSwH6D08HCJnLiskBE6SHV25XJHoiSu80PDFrFtfyiQB
Mgezqc1qRp9fqfw9Ug897DP5v0/ChBrPebnGmHBxjdJ5SQguFL6NMxT2sVAVZ0Kdew5N9L330IhI
syXr+ycLBFJvMoG+CJzSgJMO2531i0I2xI35jCbmCDYLt/M3p9f8j7+pJi3r+DvVS59vHbA9Mcfr
LnMMkudk0lD59A29vu/Tn8HPdOYSJ2nO1/aY0qWrevH1u8RDUN+16RFqC46NOhbulKRyXZWmU6Tv
iZtBCWrbxUb9MsxMQLX6KY2DGzzNIUFnJqQZ0MkPrcUmmuw+Q79tB6hEfjr10+sYoni7L0W4u4Ff
E9fa9toNUM0DSI28s6nkobGk0Xl1SbwTM88Zm2Z8dVUIFuiTS/TgkvZ1JQUkZPissjrrHtHyzZW/
ZtCvKxjwRlQU9fo0pAFAXU4UF0ZNjslkuksyHw5ld49+Eb9iuQntCWzZFb/Vl60emJmRmiCDE3J5
Vc3WjrQ5PI8+fIpIgi+liC80V//BBI2U1yDmWZr+HvYA2gd8FyYNurKwd1eZ6mpQ1oEFStrSjYfP
6qKbUuEFL2o5JlD9DfOwWZMih68yaoRYhHCb7yeRbw32y0HqPtWB10BAVUn7L1fTUQq67BXj79+x
CwJo91Xdlvi+5N5Ra17Xo9y96UJKM/FzWNYne2Ow/2iBEChXTXB9pin+Ap4HKGdDVN0KQhPDp1nA
K4ncCgANFFk0c0AuvcWzt6REtuhWiwjfrZYPQmG/V7RetC8643oDuf24iezseXV0IKbHgD6mBVWb
P27zhh0VkrbK5fuPwig7EmUUNpMWF10YFoJ4IEXd39doPqMs8I2/VXAfnCDPN1jUUOPxSXfDc1VB
ogcU4npZSR00VEpNer62oTPHK2YVGXKjrAX3ATiVEqtXYsA7gUEZbtuQpSCvBNO/HH4GwtNFPcJi
99i3B5fKmWE8bUPyiMPi3jctvl+SGn00JmsYbN4K1K5OUqApeBeMNyyDTON7LENYWag1o5ix9VI4
JXp5bIgWOCyz3YHQkwDpTYSMP67TvLqpWVihasMnxLKGdk3giRNskd5/DyEstC7nFU958Qnzv7gb
SZUXIYKz5aPvy29HEWVcSY/l1+eimo1BS/pJgadU/ihAzYFo80vWJJZw208L5IR5F0wMca7RR96y
qgIIsUOZQqlvjM6SqQKt9Wc/TcC7m72FBgI5vdVY9QtJuGfA5W+0Owe0EkssyEJ34U/3ZQIwSyuB
3DYlhp2UfmbQB/YxH4OD9uk3PsYQv/YjClA26abGD2jxrvEqV9MXoKm1pYmbJVs5KzF5e6Vg1IlC
LdDsdaqkPgzWzBzuojYPPYk56wCHB8PHYnY7s7kjH0RRxl0wSe6zrkcKMRTg1HpGG+i1OaILZDTP
Qlb+A1MV8B9f24vtomughtUMuuGk5AYguRFvKi5OT6w3+f2DSmbRbKgqXU1Xw9zJ2pKV1yV5BDEQ
e3Gg1NqWlgv8FC60ulysPAdBx3yqbLOHaxWti5e3Fe6ZVuTiG5S4y7JauZl2FlJrN0Jcqa7wY228
a3slxonruK6eIPTMPqfqPWeU3xQdD1+1lUqCRdE0Tc/uUs6r/xkFCLitNRikhPpkDwFnOb/EGAkC
WDQrjbELof+puSYiXJhYQ5gnBLQJuN9fHmTAtvB943OvJw3zTP5+4Pb4ibw3FkZ2laIzPO39Ji/0
i+N6bOhmr2QWP8XVT1mQr+N68sOB7dQG8mSoUzpdIPD9OG418gC3uANTzOvWxyDHrCtOYQxiPq2s
rUeFhOUOW2BOz9dLFpdho2r7sFoKHMnCtMF7e4rCIzP3zAwQ2gAw6bV1Ip/Zz8tJ/Pf1PGRVaatS
bfkZqqwNu4cy8XmpvOGf6B8vbEIUxzET19STr7ety4bjKGX3FMdRfa78xjvoMWxd8CFvN0QBnM5i
CKVQyUgNIxomlSH0BsEkWM5Mu4nWW6OsAOE87vtKTBkL7PLxkFH7ZWrh1kDf/DS0E4bM8aAEiIhR
3+j/Fr/5Tk2wg3Ffeib3ga/yKeuM8P+0DDFMJ+vboM5u3hrsY82WL5BUkix4WKkkuaTY5Vmo5ZM0
JMjN2d0G+btBA1rl2Al7LHSGcK4xn8iILaU266PQYSmbo5X3UwE/mG8DiLIrIIPbPpBN6UZMEgjS
CQZW5C18rVH5tb7aEpjPTNtyB6CsPxeZK/aIqlO1lafId0WWhkoYwG+iMZ3m85xq+m3ZtjlRWI1K
LoBplz6X6iXrCwcC1Veny9XyBickKQyhBpBXxjN+mYmYxCVbMT9PGvV2UU62OKOargylAqLtnEI8
IFRmyY19dDq/x74b8OM5ykMToJcyITeDiAy1yXbeOIwxj6oSHnJTlBhPeBU8JKIa9vsqi333V7p9
SJFNj88ID6ppaPAe2xIndeSviFtWJy55d1bNCHxUzsu/pMy01dz6YX7yeUFftRXwcP9mwFm1Znci
jVr8zlwj06+7fCpjawJWo2+HVDE5Rb46wvt1H8g69NEajwE5Y/FI98Su9dDtajdjVQ/7eC7xP9KI
vUPEQyjRhGfRAIDw3U+kuJbfxxnAE0Nsksw7VI8VqoM28v1dyF6X2Q2OY8MXdTKaSDimgcDZebz5
CQTkE9z9kgH0yviefprn9qnHaUItnwf+1ya0ZKLdnua21XVGzB4RVJYGg+vazeofTmviir8IYxE5
29sTGOF4ICy3QJx31Fda1vIpUYKT0C58wuwny6+JLALS8jkSt8QDfWh3ujeDiS+t80P7dBJICw/H
kgHffRNRBH2xAJs0f8E4IxUIcjX+9feb6sPsDI9La0gYlPe6mUVEh60fH3v7/AS/dyuvaSyBGsUK
/7sxx7JYmIw2xhc7hzTxuWXxx4pIr0P4vhP3Obpwj6UzsykxJ4WP34tdLLTn18qh/KEKpEyGDwyj
8d51cfxwEM0RB3OKX7Nw712iKBrtqmXP9h7Q7cSzXcEPHIyTtocRBjq/criK0Zg6c5FhF08gPrlu
s2NUKEiWG1d+0gZ7/MnZoxn2uC8I5XlecanEbnNhpclX/wbeUnnusJ54+VU6b1uuuUh/aw5b4RAS
zh56gut31jrUxanMLLctT/B6ZNxgekBTDvDbH02S5ilqgD1kVZWyLolA1F7LpASvaAYKIINwm8AI
0Su0N/CD2mqCTI3tNDhIiHwto3ou3gbOWhhoJekc287ffjE1/XfkGjsDh0IofsjSTjE/TcjnQA6u
AbeCz7BCfHEu0Lp9v4EjyLp6n7syPhsdkvmYbPaB4K0qC72givI80wtGH8VXzYC5Zj/22OEf1tKN
OheqY4dzV6MUr9KNKP5g1sX6zORFVsQ0310uylMQRFLzaI0L2kbZswIISF9c8tOR7wXmwaoB5oRs
GWCwcNHzjIQuchJakQ7RaJjUWzVUeUE5paJf59GAj18rfS/vDG8mX3M8pR36cPLvF8fQgNwTDNaa
xaCUdnweeNs6YqkHXhn22vBB6PUE0QWHVcztXXLHDJzh0y1oEoe6KedAMCOtNiNpCbct/8G3K3rB
oq5AARGWOFpY7ytjN/nYL51Y6ex3yC98OtW3t106dN7QCsSbi9NTpZQXhx2rLSLn2J0u7FzW7hD4
rl/rIQ/xncpaO/wy6R5ZB3k1CsQjLkfIDSJ6ybIFCXN3biFDoPwBPmAW4Bg4AB08mwbQfNkPVlJd
FxAHyhQIuZXi/E+A7pdFRVRskAoQsiEtigeZjwo444JpsbQ/BYfwW7Xj9N7L0EN1yLoosIq1PzEf
DDzNIEjq/cBM15YqaPotznM9Cek13KCYk3YN2WIEximm79+L3yCKQn9i8b/ztJ/Gu3UWtzTkbkT9
XT3luawo587mFKJkWVQwyblR1xcOoMFegeTPMEstNMqiJ/HE1OsAX8SZI55zHq+Pusqv67L8n8k3
eG4NPM24buuyCNEocWa2NlBYamFuNnxzZhEZuRtqUuJR2iHMGUZ2Kukqz4GcEgrPYkb+16lbgWMQ
l1SgF8g3rcvQridZA7eeDKKCEDEzXqYBPaNLUA7F5LujhvvWKYh9/BkPpnTdjpWE1KK5zqXGk8b4
/nkXV7rSOnD+MX4CQ/49JZzFzk+K+Q8UQ72cEMhpomhuVt5RAD28swDwVOmcC9QNrfbzjmIHe13Q
a2SVnvsA6LvTrSVYCijzrts02dDOlya8A1qyjS1vVpw484aa8GLXO54JGF/btwdkjA5tjTNSjSSt
rnc++6rUykY5GWihoOK2vtHzSLwzSgIiEB8/hCwXiRytkUE0R+uMNB5YD7sc1NH0ZHrgNnWyxAyE
lqtPAg6zYiTSXTSTU3r386Hl80vBXaBa/pDvVdeuMDrVtKxitC7BD27oHgDSdMOQ275qWXPkW83C
jEkUaNBI7BoY8tZI9QZi0zQRP+3wF/kykNdMKU6OemQIlHn80q1AkG231hYl5wcdZlUtglh+bMZ7
XKEcueVeHMAnUtXrDmfYc2DMs36os6EemZrIq+TxCgNcMuFbA7FxjvRYYvBXYqv32ZTb9YuqjFkw
ES4b2wSATDbCrS0iXnD3KiL1gQYLgVQcRcxA2WPYUJHtCS0GqazkrbwMu54D+GeQCHLA0cGuVnhi
Wym5YF+zxKyXKBd9XZEoaSTrnToQAoqizA5aYv5yZ7TOMTJx8iJZRALlFwe/NL5Fj7YAZxJtcutV
zTrgXpRcC0cn6Jszwef5uFn1d2ot/6pIOcgvJ2UZBDHPYAC69XFswmni+UcHmuT6wvBwFP92QLfc
vKifZII6905FtTHijPdzd90okScTitc15i1NlOiZ7SCi2PXiFC+eG6p/qERg5qeq3COFtT2mMMX5
alKPSQGuZes6ikV+j0fDL0SLVAOADiXJUmPVXo6hzljX5KhlAkYbQacpUNtuF+HQf5zMZ10Xl784
8eUgW4+i9x41CFDrOvvbDvg6DEMX0MPr49tYOboF3zVuKQBKTMA74bdn1LoBGHXmRDBHqlc/dX31
E6dDN2rtIU96GLKsC8GUc24tX7WcZ27fxjQ7Nv6UsNIZYecbKlDsxn8tCGIyueAntR0LVqWA2QHh
U3It5tqUrANZBj2QwEsyD+6BR31nWdl3a7u2G72M24VzSQJF/VmgyiQ2ks3zGaUh5wLIyMYJ72FF
rfT00T3zcOKVs6P59xWUFuyXgtGafBhOCzqDVcAlEJVGA4TjpQ3EEf2hnA7+AjUs85ZeqZfbObNm
7xXJ8Hc/Zkz2HXyyCuTJqbBPgC2R+gfgekcX1RVzUuL5kpDY5+TTRskYuIwXSlSV0schWdYybMqd
WlV1At33wKnwcfCPM4gYhOzTL3bESAxpYtRU0I6nTyvV4b6N5m2WmiorS1VUjXiAtuiUWxHX7TJ6
KuD1SccWAx0ZLIAAOiELPHvv3i1fxAeXRkdCDgdGeOVFK6a4FI3FAvsbHqWI63HDduVfu+75xaU8
lTgMUmAfWfVwMk2x2e8SISECu+nW/EEErZmTIFmfcZtE0RsatUD17bow4QFlI3ctuMptO2XGevrS
HJB9utppHN0AIBhXqzUKO4EkFvXMVc6IBdzLHcIgBFcWpy6OP8MCLKWxSq9t9jATWGBUEVjFcvJt
xZwpDUe2MXf9X2eGSFmwEO7K3GhBHEmhCKB8LvStV6yWLmhSpLV8kARsOdN9HEBzcE3WIj6Bbl8+
danININk77veySX5hfxD2VUxEMM/BBiD81xo2RkYZpb3+IIodlP2k3xmaR7k0rf+DE2o8Lewg0PF
SC7CcCbMojwlOSboNig6NY3uChV+8ke/VQ4OBITcntcXgiSov30zvpyUdZcy0RM4Hp6Lyrc8odf1
ZjqC0Boyy0VfGIHnaDaYMCVj1hw3o8+x7BwM+dA8eZR30VD2+LfucF9i9E2zcqLxqvqO4dPvM4kF
2mfmjgqLHDWpAm1Zjvcmws/WPTwKwfOF/NrOiQEJ28bTWJmZnq8GFS8+MC7utNnPKzKydfdbZTre
4pHuD37orpkQ1OhjC5+kvP2kHUvV3Dl9taU5zEM8G6VSkjD7wWlyD6RqvJzhvbJ1JiBjQRw+5b6Q
U7p1/Qi1V7DxRo9rLPVuLkjdO4vE+lZvxv9utlCjN2iZIkWtCuVr6b7w3vEF8Ok6suT3NXU/I929
2/vYRwRpyUleNIaMzIXMB+a1q4iKLEQJ7lxWkPQTd3gwV4jAdb7QZ7AuKYqqeuSsmb9VKdtqYCWJ
Yw5m+5MklQuSR0Uxc3gvV7WJ/dvOUDFoKlWUt7w97spKuxqVepfa7Ncy9N31cge0LhD/SGBwzvWp
v5AhuoFkH2Y0S0xihPs7G6u6N9xxrAI6xYlTaQ7xoFtl2R5J9jH53b3bCBXCP9Ruyf+VcEMhpx4a
9cXs81Njc6HqfuBUemG3lYbXZd7vDkhLhu897LXknlFtWQ4Zzk9b1uKvnVIDlGVG3RgYkzm2rZ8t
Amh/vnp1AfgUp94ofiWrFKzytMGYKFVHDH/sV25MmhEWDr95hwcEEJMN6eI3PIr1E6Kt1udVw5JI
tY51zqLU1vJFyYvrXZVZFFsmE3yzjMFE7ZXZVeiKkKVn7jSC3+h+wrfRfxNVa9dIN1S9nRLE39J9
EeG46nO+RLn9upOd3nHdgl4tBOqmixNsEZVeFg7Fir5d55Z2V7BT9rMAAutPVOMmweqE4QcQZ1bG
B+5TV+aEZC5ns2o07r3VfZT2kI3U6NMyAP6cBawFHV3oJ4DQ4jhZKgC4yhJhebCAaRGv/cFrq78n
N6truenbSfflyPa1QjNWJg1MtJ/qDs7+BL1LJwXkpYyNdxP/7YzOPnxkvkmBg5so3aX+0pBqyBQK
T4KRGy5YfxwjGADdgUeDmfX8E3AY9MIdaUC9h8mKMLFkYrlKphCtwaKYqfZAviECIOKOLFxe5ezO
6wUxrHB26uPFBmNeUoR6LSWOnmsLmmjC3xJgb6BghTk/fVPoG4hHJud/IShfg2HY9E9ze2SsM5RK
E4aR7CZ7O4k8Sdln9Qs5XGNB3HPgCjCaTadZODUxOYdsURwL6bUnOrE15V6n9SqqNL8ADUmpKNh1
chLlA/TmdBikfQ0m2fww97n3RAyouzj51iVJWizvIJR8hH85kx8JB8ASpnLLuerarnYY0IqhfRCg
pilvhS4Dz6lcZo/6RP0tc0Cgtrl/ztx6Y3HmWUTz4iZm6ib7jJ+a/xUbZ4cjNSCcWta5fHVztp9o
ULraI/PJL5g9GuLwxzipI3gghBImF3aXKDpXx+OXSWC01pAIEahw4rzLgUN+wwV1qR1Qgoh5q9+E
Hv9PdxIYTjbaB+YMR/9/6/lEbSTAOjbTY4C0+c2+lqWdXR3XgBRq40GX5i6/z0y+Xi1iixbxR52W
QcuK2TN8ir6+GMC9/W1STh4444/WLga6d40XslcE6RHlanW4MxSX+WVt7faeE0woPlep1Z5uSUrg
CkurdYybbRs/EyZ3IgxlXEa94s1RWeXQ769NBkCcQRjKybdjgWa/j42DLzcYdAzvrej7roNFwkFQ
/JLY8zCbGCJ93gSODFLhvXdzXun72Hu81HsacpMvuxYXN1W533JSpmXtYyzPwDpUxZ03UqM3SPSr
2galQnPUsjE+aFmWjZecrgbK3FR7UUHs61wT9fcAKvF5rt8wOfPRfnviSunQjRyjOUxnhpRxG5C2
jh26WJtK6zxvbsYTQGSBVPBTfwBjHZ+yKip0/8Vf47AwKWo2odUsDFiXD1wE2rIi+3dhjRGE1OMO
U62K5xe6SgVh+UwX+EdBV9pFzBcE3FmQhV8ONuLIgpajBJlF77Y4ORHoQipMQ9aYMjFlRWXhJhmK
wVSNpFf/krsSarDv+icWIqrJgoyuiK9tdWsVpgIfu0oI0gNPaz8ZMqQWvbGnDdHZsycg/RGYQbY2
u0p1fZBcKM9o3t23WlfkZ8pkPbBntd5b6Ib7X3IF38hE9T2+NBZ7LdMyrMki6t8Ps/JO8Ndslezb
ohm9r/X19ctvA/Bk4pkT65RSu2qAY7Kc2ItukFwUCJ0ISUGtVGDcydr/RVB1M5Yq3y2zp55gN3cU
LiLGtZ0zSRrUp9jOoP1jtPjg1IXk09U8dMRF5ujNH6BQCjpiyB6vBjn1sHFsoFg8UNtv7gCAeEWj
wkwabuKlnGwyIHgdcDpRWlB0N7t31tpfNwgh+RbqsMCJ2B3ia+U6yeqqHkKvDY56mcZDbuIzMEs9
EN/EMV1xj32itrvjVuzWZWYD1jtfA0RopSeaOa2mOF8Z3bF2DRWywBeI2R1aSGs9iLY34fQhxnO5
CvmaJg7dGl96xb0um32M7XlalcJ+i8CHyoC1lDezFTjvSX+FLHbQGxx/gRy5gNhsc2/eKNmg8LGq
FKuA9CbgdYUuA8DrRXUnlX/djDPdTjdTanJq+Mnwh7Pfo7KfODWs1bpyTvtk8FMtWvDRDPacWSEE
eDtXOrJne2zaTbefygbO4a7bBBXSetWH3Yrm/3X2O+vutaJqBnewx3HewMXC9EpxPkaop+Xi7Wwn
aWB0JghM7HrvE1S/f5Ye4oEhSWj/t4A/X0BmmWAMNmy8hCJgNjmwfESGzRPsebODnEqDJ7PITwNa
V09miLRgnAVmdoXDEG+tpMM0oHMpzXUjiByJQCuSlAoLT1tYtjN3u+hOqhx1Thw2/6D9PbyNJ2z5
EzjUsS84GbWxBWfxNjACpa7Z7wFKKnZSYhf8d4UChpwDRYHK9KMR535/qwxoi8zGNsDpT5vJXokY
gu1bxrc0vwRhZRDTzKo4tQysLC6tqgcyLxVYUEiya5g6h+Cnl8iKNPbbL3V4+8ZFE1cZY0z+oEeq
KwnP7o2NxdR5EMypz8cZ/EkHSZpm6Y1dx8HyedyHRUm1dIdhi0y13EdUbDm6UjaiXnkOuaYmYVuo
xCkc2juBAmVnpuK/5hWxCGdJydpPlUVKBY4yR0kIEffHV0SoR9eAnXATAl4f2nZUhZwKkQW53t1l
5zN8/Tt1KXHlSHwujNTcwqjE1sU0OVldbwDUwAtMayMS7yD23zTcwWjJ0QFp7ryGcV0+N6M4eLEo
+B7ywkgZRLGK5ZWOeE4gH3myNi1wdtF8OAbzMD2ZhK7huOpBEDi/cYdTaE+qmMPjfY1NL3LXgr+Y
DlXQq1i2ondx36amFGceLiKodbDv2dQs1CWM4s515oBR9EeF7r5VTIkq+OE7JhOfVeycborcMzoF
h232pG1z3QV+q7KN3sgvo79JwbDoAWkMEqEITopN1I20brMJZun1gHX8Xc80J3iuXc39Y2XdxDZv
7UakPosECn1cVSH1ArdW7amFw1hZFRWT6b+RSMKi+S0oqMR3oUjuUR7EoQQl7YODutQuQ4NL67mk
+aYvqO1QBsLrsPzYfIWgifETXNNrD7xKtRge0HaTn6HpoLtKArPie/SFupRpWzOtonghGPlKlFaO
ql29d0fARp6wP8OtOnS+OKG3JrhpGTtxx48sz5Pw1usBS86osWV9pCs0hW0oWatfq+ehUUBXF+OZ
kMCyqUiCoG+7UE0hRyryokxQoRhK60JBBrSpMOImfRm4SrB6u/FBBnhMjf8k2pTAeU+cKbw/1PuK
8/bQhPzD+JPVrLSC/DnK7Pd35Jq7NAw/ogJ5/vTvu++oBcbiKj6MzShj2OvW05ZbmF8XkaH6/udm
Y/XljGgYl+yPMfIF+7EdVBnZs5ql+rkfvCcyqgpJKLiLcoBjEjEwwGJnHWvK2PUzpnwhwe8x69pf
T8JGTqQ9FWeHZwGpA4vqnUzMxDa78q3XXbJ9EGMw8KdPAORtvuIk36ST9SW4cHD3PZRhQpVRcu+l
uOvUmwib13lcu3VUW1bKls5FXtrFqifnUYLosaVuqIsNzKkdflW9D0So3hxDJLFuHOjLf0Csjgw4
fzDFSD4bjq/d7bzVKguB/vl0q/myZMiqvZODedwbx9j8h8lOpx0DquZTJuiEPxYkYgvkhmXhFDiO
LGHEqA78u7zbYUIQfKlaj9kF0gxYUm62I++ywvUDg8D1WVryALALLUZJT6AKlsKHnuRtNi6oRPRW
LmlaAMWefE39Oa/qynOeyagE8EeaVPvTIUmpoj6FbfwQtRUVyT29ZiCP8L8BEeiDuRE/p2r5SKQD
W1sheMsX99bHxMDhUJTv4MdIPFjNarOn5TfwRaOzBw+DtwQgMPY/lU/iXHa1axzda4OGbxtVxMG7
CRrL+WqB+xw2Y4mvjRpgNIchllWgQWroLZclBq87+/wvX+vvcGztPUuHTjYyZdidrvY6H6etp/xL
Mwn5qvC3u3mkCBUBWWjRsw4OaOalFrujRW+CbgGus9QIiN4rjK62PHW1vnX4vlDn1B/SdGmwzgtK
NpTZJl3ZhXn4zBp+uHAdSneEtScJpcdsyuOvuC70Kn/Eh4vuMoQ7InMfs4A+LLxUiOQ/bELnhisR
2lf9ZbKbK1hObvwsSalUyNRZLhZzvxYdaLYiS8n6HvnZKXB6VJ9QbKHp0e1IeS8Nn312Cea/uqTa
7JkTrcLc1rd71mEYNEZAfSv0NM9VRqnP2PfrCBqUmm1AQEq70FjDdASi1Rv5xUTkmbloLN/q8QEF
bcf7+POFdObgni7giUt1Fm9k7E7JOM+waMzsaqgvlZ4pshBr3IYuLKfrm1Bua+Pj+fo4rUlzwaNN
7KEWo+5Jf9WXsGXKWdwgF7mlaKRP12FinmgkEIrj99qdJbS3tWeiIfhQPd6wNeEuBUt7BXDabAsT
K/IVZ71qDb/yvxhrwqGw6fj83MYII59aCE7hk4c8lB9tIKehHWSJ33q/WHIFC5Sa8HUK2M1FSXoh
v6nlTVdkjDRLtsOE+rDocr0O9Ymk6tboEmLXMSPbxDuBOZCNQFrn9oLqqTqOV8QvIetQ+GlmYtzN
ihoK6Vtfsps1gAh4ndouCrq/4JCl/+A8h4+N4nksbscmhRXK0tc3ra3yLMiTYRJU+e+RjHbTfcoA
OKbXxUUOGmyLOC8/FMKPz1H5ju27Ode306azyBnYZjUz9/o6wMKnJqAv9cl1/oV22cH14u93JrUc
rkK5m6S2w8IRrxPQs+KjSrQuFN6H8ypbKSZXCxbefNgDCFewq3Y7EzzfPaKFatiCrOIZAYAIbtjB
zmn078WVLpaAAwrLaxnEaXWU2lFCHmhKFHvBh4icNUAhvmIOT3exEOtyk6/xOoyqgZpjc+tay11k
xdO/hZcND7PR995X6f1+rFfTBd3epwcWfrqlRy4ceqJZBej63fHc501swefKNnC2iMyOkKw/gYgN
344gPe0ig+wHNF6/7QzBuoijUcKw42DW0vBHKXFuwcQZqCmc3NfsRTRXMabsaI0FiJfFrvwUZ8an
hmtuWcff/aTziXlqwA6/c+qziNoA3zXo7nES2/l5tj3ZtDSW+PYCWb7kz/WPe93PN4BchnEpzmv3
of5FY9IvHhGhHAA2BMPPE6Lj3QU7N9aP5QPaMQ1ALYMOzIxvMwp1JrkaNTfQtqLtZda0zgRqiZ3S
zD+FTTV5ttKiVXpDskj8lPd1efleS7eugPfxpjKiikJtOqKCeGFNDtcWdfrj4tlSxHPpCC363bHc
YIJzHCTEXC0uhGGNwBWkcWryoPhiDsVJF4c2ar5AJzJXRJwpKS8hS0lbAax3mgWkfL5Wr+cmTb5s
uvj2rPzqY54EAiY84K29DNob6c7gl35KOiWif1+jWg7RcJ1GPOWjp5DNBUK3OCOzwT1UJcJxGgYH
hw3h+/zYVk2p/6suD2uHNOolf1ww/qjwHdakoIGfEGXsU+NBFwkLbSqAGb1rqVVEW74PM3u32h1N
k0ttijoJOUxj5bvwJH2wmaLOUB2ZuIQvmqNDJPpwS8V79l6zJ6VOrvvtlOFi2PlfuKBKUqRcOoDK
Tn//QXZrTMyKazt5w1OUIG0QVq+chrAjqrIUYP75+OyskPYI6b2wi3+KAaDtSUX1IBszRRvU9tNv
yKXPHqDFgTdnVUv8AEryDe1uqVNPO6xHJQ+shvujpS1YAkeIsSdMjh9Q9PTLDyNcwhoF8dHlu5QE
VbQWGQVTfIulb3OXaQhVgblBbOtvKdhTZGzg5uJm/MPMXovHvX09Qkp7R3rzCFHT08FgJklElY/G
6x9HHQKQcOQUoEtBOJhl2+Wax1tEaW0XW6ODFtOQrOCXCc6oPEU3ovndstrMyh3qIg1JyPX4KRc7
Dv4bMEHcRRVb9D7R+xEuSd/x5vT3wmcg+J3SHbEhtI6tGmOF+X5ZV4PZBBTjfFB5Ont9dB+JMHhc
S1c1f8R9njiEy3OApch+f1JOadRCaHDdrEEyZIPM2kNzwwrgLEYFR5ZnWz5w7/Qiw43mv3smIw9C
KyeEFq29tl4qOXhGE7xSdkavZGBD0ufhz2O8cszBs4mXstqTieRgoo7+9ch4ylyc/rFj5p9oRsOu
pjJqsAHBrqg5epVi3P5Jo0hIB7NQOYDq0gfFCxwJ7jgTgakUSIkrVSxV8tLfTciYeJeOux/L2sS2
z34QdcMrVMb0A9U/l1nxRiX5QYji+17yVxsgPH31RU5+uUYlXjgVVMo0iEaKw1efanRCKf3uoVab
OwaNRVl02bGIH76PBAR5yis8Ba5Jv6O2YsDC9XPe3I8mYq/qmOUc49MCRoQHea4jvU0gslcVfAz1
2om756VrFvDn4AVtra9tDEs9getrzS/Ul5DHVhd5QxpUvqxdOx18nsghKstooaBTcSqXT8SvkwSD
D98W9cYXMuFkeQ6jDQtwFrLbrnnfOBCZfiOiU+pMxNJkHmnYW6QBDKSdD8EPBW32OQ+IAy0cXCPf
TkQfCrCOfLF6mAslHeDyGS4nqf5tYRhfglb4mlxLAWgsrVpwCkgOgsdqsfi9lRwsHq5LNVcVSliX
sPDf5ysWnGibO5C/O8EG/NziKp4BSWpn3g2qm4aJfOXl1I96tbtPcLxEUFiRxnR1BN5AXF7QfJkJ
l/eJh7+eiYPHCgZsOEInaOWHH7OFrPzKG9LORu8hYMsRbHFNa9+ZUavBIpcpMQntpqrmSaIwkBV6
LUIpeHZMzrqAjnMt5EkxM2jI2z8iyJiMKdijvU/VbaWOLgEMMt5NQlgs1IBHki37L3rNf13l2ZXp
+OmZqxG/10PDls5zOHQx/QiagJdn7eV3C84WtWsk0+v/RG9J+RX6HFMr/kwSxonwX+x0emho2epC
JbE9YPQXVt48uKi4eFk5mEYUfwzmtVQsOPgBal7KzUWOaVR4AbsI4A7SFDnmqynqW/sA/fKREm4B
iznArRsYBzTS/b8DgEwuh5/QeyGkKGgij9tBuAZbpbwSRGcWoDu67/G0CH66Lz8dFbfPd5JRddDh
SDMrinu4viuPugQOi2s7GxFMnQPEdtOHtEKrm8YcyM89aXh/4dmt31A5OIKIXQvzrNiiW/sMO4oz
b2h3uXyOzUQtrb1L/BBvcdQIMEgC8ENusSeGknANgTsA2BzVy1qlcQ1hslEXDt1VZMSkoLHuprvP
TK8n8tRB5M6+248h6RFJDujpm1xilTjFVq7isDJALc2IJEiu1Lsq1BxhSeFm03EW5//NmuR7Fb1v
kHl6TMo2Ey/mRFu/H98mer87leTPSmsx/j3hj7OVLzm5gkTpJRVGfLYutXK94xynGZq4YZdSXszJ
xw/zB5w6yK1n8O4ppzSssr9bf29nk/oU2q5hpZqUwgY84+Q3f/OP4fWWkg0oizpyf6GCe18alizp
OuNaQgnnHVaJe9tfsvFDBrS0LLanL6WoJm/FxUkixkCdIihZgNGC8xL7lFJEwtU3lu3+79W9YiY3
YZHCRB3AwHxIEu1ioXu81YrR6aEM4XYXr/paJX1LhEArP7Uprg3q3ILehofrgr7A4SxFda4DwV7p
h1qG116DmsXuMluZNt5SZKdsHtEvdNFhtbGKgx6A+uxDZBqkksqG+HGu/BQdWUUGWINnKGY1pZU4
XDyZFXBABnDLsCbcbDO5+YFSiCqAhzZSsDqtAZiTifI2gsdZHK2FHpPx9Xy5FTO7dlbk9gIEyin3
Teg4CchQf9fsZ5Q+ibgEDG0PU8fByOQX4NL/QZEh/OcZTQG7hFyK+xG0TwN9Dz3qNFckjv18nAok
Uu3ZOZQePH/OXk/ypie6+4FK7nBl4vs7/CnQXAxsZHhCkfclo8pnG9Ys0CqfR3rqN59Bqd3v6zRP
ESwCgSgJJPh+cLP24SIcWlMG14RWiax9f5IUHkfr3NOY1Y8PKgbjEg02+SKNiXjCsy61x2A4K5yB
eeDFExIzUb/O72JXm1tKULcNujD4C8gDQPaucWyYI/9vB/jUmYk15G+blouJcDpfXUhtv8SRPlSp
hcsSnKvuqQxEDH1VSy2s8ElzDHcDkAUnltUz5qmccR0Dd0Wq0f/6jyeo1DvX+gSvevvMi001cHGD
r/4kQzA0e1F6EohzcBdCh/aemH0bQxAUpiIuvpG8S6GMh7HqnNUthWp1fLqOd0ieuXLN4ioyekgz
PKisPLIN9iBsvMVxBeoSZLTmJ0JzvxCt/ZL+TTNtXfD6qsIZQG172HJeRenXVCoEQNNOcpIO+p/4
9uqMCRALIIGqCIRk0gzoRIIbxDiD0iACPzhq/1X0vVd3Bx7ajhUJJvuHLregOP29Hrz21KM15k3d
2edECNap/Di2UTU8+vZaOX/cMWf2GeQlJZaSEHI3xEC5b7DsMf7lhdF/5ADy6QGgo4viEUqSpuGp
C9YhNNjlb/AW99Ysi5R/NvGGq71h7Lx9Ew89z4A9wQjt6bCjcRwE8mtXTkgQPA5jS8U5DmI9JAgX
fyklge2rIrtUnKuZcSOM84B1dpq1za0192pf26f/N1G6qFJ4ZlYVd8nFau9EXQ3AbHI5m8GgMYEB
jTXMyyBEb03GpS+dDAWakw2FiExNtscbv9+ra7VWkFx7ZRSpc6XQ42wRar68Xk6H8xgaiCTN/mvQ
hjunjfMbbVG55JYGVWgtP0e5Q+SCIw/LBBvPtLkzMZogs6cUw9+8vmjfKnK9rKWVUolVEDdIBP/o
215lov78I+3e+9AQx2BVxPgsI/VSltMlM6iDExS+zcfsJ/8czBQQd/vS8GrbwiIq3VHaWuXrDmiE
Zn/h+lG7nq1rJ9uNbyEomE6xjUF0D+XRzP3X3YPr30haYb+DWo7VvGWOPcXCDJ9jD19kbB24qO0c
fjIZnycDighNg4rl5hjN7WtkUj5xoYbTvr/XK366hzubSmWBW6HmLYdhy7eq6LNE/9AJc18hR2CM
H5JZb+O5Hf32jojuzp614Ey5EaemWaZjov2rpSArboKgKA8zPQJDr7IQ+cgsjZZIwWysog/98Dgf
RclCUQhP0guDLlzJttMWqtnHLokqT65xObB1JcpMk1O3CJizBw9DbKFHBvHG+KRxlv2LW+Mlx0ii
11BEukbZgCIaJ8xUokznqR2MuSfu6mtdXe632DoI/97kM6+zqzEuzS08b4VkKyarCTu0/G/sOPX1
RXbwlgtrnF4v5mOrisugF8hJOtXLUJL5nHIKw/kQuNh+I/HdORT16GDP98mHky+WqSblWoZfb5sn
iXEmIBJlK7rDQ5ym0Bx3054oxEQlv3gd9b9auvIwLH/SH/TcJJZoyZoTfstX9q+UGbzczZVBYLeL
4xUg3NPIrSpP+WTemNHVwf4ziIo1jAMHwEnc+5IJ16o8EnCXpO+P/P7EsEGxV9URO8zEv8xOrLp9
/vloCrBmLHbdyjjsugvyQcNfyBJncLfxieU+cqQrS73ho6lbOf2d32Qg4Y2r+r3FYZItvIGK2JaE
Bn1MQVpzpPqnoejjyjHdwBrbx63Q8cULcw0i5bM+MmNdPMh9gGWcTOQwoKSfQEvYL0t4oL9Zkrpe
xedBLQqXSOal4tWhvoDrCZBdJrOk8ZZc11+3nNsgjh4zWkklVrw/CD1jUSgiOF0bQRbR4B6CHQyz
aSB21DtgaVLFraNSu6tHVqUNd7dZmN6B0ZZcKU/OA+97gkPohYnMCwpFFaqhSDLqHNOY0E4oKAnk
Uf9naAMPt8w74FWbJE4WE8i4CkWigaNXX7qsmMb5BDhodHcuuv7jRRodqEPSpYdB0ZFlXUidcl3b
UB8Ognjh4+bgORtuzWMeRVTRqgfjJ4odcv4x5culh1YpeeV3veu4qIO5ZLu97hVf327vZVKOBKSF
gr3fTPScH968ymASv8+JXNJgeCdZ5k1Z+jMgwGJdZB6chv/VNF3TgkejiIzBkKoMRM3SO/qqCM/Z
UQhqb+2ES3OMMzwTkMdBzsLSRawvMLxFFfkdu/qhWFPbY+FT4yobpUyYr5Sm7w4KTcwJggYd94pS
Y2QaoM0sqzC42QY4P1Obm8bc7ajB3fIqvdTAsK7CLifN4/rP0pdRJQnMSSurZ67fYCpqj/gm6gdQ
2k1iniy8jhvNldX4I5aWPuaX1b4xqYgFeJLt+0Q7wbS2knJ3BFsAcNivWX97Bq0NQRopfCG0Y3cT
tW9DDypNqTJVqQumEcvssJQtLfrSVIqYxoVisnGqE4A2a1vPeAx3g/xGc929xEa56ADsK44/JRep
JwxaCCfYh1IF0xLyNe1m48RvwMh/lAAy+M5U5PTvQM2t1LquqtXULwDx/MGZ9tixJ+OmKSnP8Z4v
dcv59Wc/vc4IeWy9HGqVGkCCBVCoCySTneUpngli8SoNjFlxklAUdbsd+NrsE1xbS6Bb7dSlBx03
+l1iE6g0lAlX5YQbCPS5GnlhxEa2GfYgM6C9Vb9Y9HxRnoz9YP667JghCcsFci4F1RWX3mN24js7
eA0k9pNHbYLl18VeWhKzdzs38nCe1tOkUaNhdgESUrhTjAoJIZS2NZcZMq3tiUs1NLvmH8phRabB
H8eBPdtD8bYVZ/f359bcyzz/aJpkkra4Ekpvtj+HD6+J1rB3zptfG3oJ9tymAu7B7JCXui7jk6/k
DLS87kqhxK+1mhTiagOAssDrGNXOWpobVMbQfLIvnytAcYasyIKMO2CPbphoTY8FsiSxu5BgUxik
hvYh3h/uNzboSa6XAJ/nsiOGDwTL3M+wB9ygWWJMDdlhFxhZmq48grfB+YVpuXskyHm0KVKb0n8c
MfUCXyxsh+E7Z6YNQ/N33X8O3rk5I9JD+4mHq5lbhpII4bYLiJNd7sQWboiLQgu/z/n0nNx5SPZZ
aZydIou9wZz8DfGsTCkQjQ5JSJi3qmfJDJF+YMOrfhfP+AG/CoE/84HG8f5Q7jKpoMyMYH0ee98l
oaxV4aS3EOfUlK09++MGsv5mgqn4n1hRolNgO0/h9nstFXhgKZpg8vrSWCxpMqfmMoOhz/TlJiXX
blc8r4UBbIcPNAur5WDTX9uZzIG1sC8CjsQ4Hn6IsOS6gKnymXkwppago7hSoDVsyczJ8Nsc9zfX
br4BRBwcnVVOikcM+Yjfbob0ZdLvbvx+WHfQAUDuThkhh7eRUnwUefRDNOopUSdagyVEC+qi8LpW
MA74ZBwqpBIHIQWXQqGRt8oboX9I8XhAK3IY/Nwo1OG7pwjK+4apcEdPteTsVOYy2HbjDLBPWMpy
T1LsWxbh6RNp9jX85KTMCNjMYvN9uyZq91TtKHeKY1SRdCHeWN4NWd4I4ihucC4dE2SgjOWOlg95
pQZTGrOHsknz8BsOFwieHHk6swZPuvbCqPRGuXQkMAaPuASVnwvWVZVcJBMF9JC45FLm/2d50Ac4
CS8yuP9kU2Ln4miP3Cu41miMZF1m//WNAqUoOHpPPnMPzTWESvd9qMh+rYYFP9voDdocechmfeda
Ke4UtjGv+uWf9/V7AUX0tFlPtmrI79S1Ny71VEDAWte/t3STj47bgJQqlOYUq273Hl4ff2AuPBcY
HfiZ4giduKhFEwnL5t2ErJK42Rl6c+YU7//HuFYc7Q+KaTSFciFXAA5jZ0qGYu2Vd02JpMeuv6MM
OJtFN67UMAw8zPod1f9cpaWwlJ/UuTURPkGRZLEnCpOHNr62x7DjtnwifG9PSvcNkt08q0LUJL+Q
tL5ZK5SmAvlFedi6BoaYr6snxtLJet4lEwV7RZWAKwSmEjoKLoMav3S6n11AlHcOGt5kdCJU0OLx
hEjyms0/DRfeIZk4aKHw/F5/YazkKvFhDenNm6aTHOv0h83JMIqr94wEaNxQCgnDnQtri3zVEkf0
peCqNuV2MdYEtEdj3OSDRJF/p5D3O4rqKJNHzszsfVdVFzYJ4pbM2fowoyar6XlI+tO9LUw+Fs57
tqcVOuou4nlMDpYhpDfeSSGwapTfra7Z4GtQgi3TvRrf0szAyUAac5MkKVpydwn3Om5cS68LbbPa
7/iEufquAkVTryr3OnYCyl0+zellsn3bpNDcIwNrnqGiZJIdc8AGb+fC2yH0Ds5XmUtd0RqyxkNC
2vUzz3OwItvh/taWPgTLAVLbd3/IOn56sd3Gi973QBC7w/ebWntsbZmdy7WQSiVtbBIMv7acH05l
uTnUlo7V63oopdkZaW0QorO0e+pL96wLhQFtSJYz5EqwBxipoUgZGSH9xJVgHFTBSejM1PCCra90
WsAkB0wV/lVIxNhbymHn6GuUiCivCIIzQ92axJ/cA29t3c2oJ0DDHhYnmIqZnFDOcD6X5lwz4meb
vgavLABCkF50M8BqlaFm6Q6A9E3yzvIcjfsUZsyqko7iOcdxBWf3MDLWUKBkv7l/gVhr/NYWGSWC
SGMqL4ryB9ZmHpdyg9Gp4x+RqvY5iTAtd2oXcK1Ivqh+Aa++QBVejBNyHvTL3/R2cMZ60X9NBaWF
1sK+jhzxOgqLQ889PiYrBBevWyFL7lIUK1L6ZUAnLx9rq2aYglflz0L803SihiAbFA6aIeWUi1Zg
eEcZJJ6NK84XG93ji6sURag11xZIRDSpdMlbArDXgr5Am8DXzrH6jeh/BLw422i6svbGxOqZ7N7p
IxzAdi8Fvhh4X8QUSSHMz9+TfyYYtxXUWNP+h5eJkiMZcow3dHI5biqbqfJQ82o/eyvXaMjzYUVd
UgabTdTQb0cTG4OaOTfPVXi6GbGZ8q6DMoiP3gCYkVRfSMeOnqFj1KyADhbusjlic/prAL+VV8Gt
mcH4A1w/1AHsl1p8doisZh+W+dy/ija1uw7ldQgfsvRw8KhIYGYZ6ncZbm/lrk9078wGNA197pfF
HhaAo0LUI325kvYQlPT/lhj6PihpHYzjsXlPZehe3xG1EiQuB7N2nraByqda6Xdd+0eatbEC1+Ct
cCnPvKDFcC5JwmeSbIk1trvm+EhpAsbTv/K/wd31lh2oUaV8/faYZ6vHzTk6fYZj2Y0JGgb/suzi
wzv2nrne/upztjfkxOSR6isuufDrGUGDMJ4NogSksS90yysZrmR9mGMltyObK25MdipFsJgMz0N5
vpXaI3ojETd0qxfrQIf8AhIxejbk5dakUN1dEYNe+gV14hfVocjXt/luH1CCesujOfTZ2MZNG/pS
lNdHd8ho794+H7yZDmu9OVZqzj/dOhNPtMudGHUjXQcABQEorhdtA8rsMXOm4Q3QcF+n+Qj+rx/+
v9n4LsBbKc1FwnHfB04DLlvJDO5o8oye3lkM3lYE08pLcmNNi7otpjXUuGGP/TA3E2+lh0G1T9z5
BXQVteE14dszqNXrWvpDuQTNKPXhmU1AJ7jMDNSXq2fARjHIMgjeWbUtL2Ix57fAsy3+KTrdy43t
+MhLtMz+3uWF0rvm4ZtY0rts+LMkWgTY+qjEwtnDjavdv/hy2inZjvBqCn6OXr4OH6NvIi+mQU6S
3YM1R9zWMfsKAUHdbdmklRznRSAtFkf5J3jEjOhsuEJRVKIbxrTLg81eQhgLcjy7njwGsx8nLGeD
b9yl2ZUKBTZh/ApFzDOuRJDkN6VEBJvv9MubEova8paLuPz1Ceum2kMhfUp9e7l4FdqaIefXrkv0
s6fh4vKE2M3y7ar8DjScZu2SCquBJ4iPIzpx4Uhmps3N3Zlcv/3mcoGwER+ESW51okb8Zum/FJiN
cuT/qFjMj4I7qeL/mFTZzjb6YOJYvVWH/cXofH4IlYu/CgkgQp5pVByHhEw0m5QEbJpQqqYEn02V
Z4tgvjGouTqkgNTtuM+Z3kSnlvK1x3oyhgrhUu9C6ZQsVudqxZx6bJy78oA+wdpxku6Q08eTT/eU
SV4qolkCTgJa0LMKiNNKtjbJBJ7BI7rZj/ey4uxAgkMZdlqAQyuEuclYTX5IgyV7y6b9Y0VaYb4D
N9pyxj1mAtBb67yJLUrTCzKEUHadR5M3ofd7hh85JdAcxYc05QC5lnh/3INGdJ3glA/ihXf7lhgj
u7DBdDPB1JhyMfLwUKEZSKll2zTlMTCPG/hOwSfwlh2klqbforgPEoNfjjgozxf+qQPas2L8YXIl
TGERcnUYExCAKJonuBn6Ym1j+n5eSvKlO2VYNmlPkeq8XdDIQgnBB5ue6yHx5jHeZk2NOoFwf5Ie
Pzzmat3HYITzIDHxgkgE+S/fjz877qoftu665b6RaYWymXv6xuS0wI6LiwlrPZDHoqsrkIOdCiUs
myZNW1wRvc2y98HBT1viWRlSomQGIHSBEMD+MQ+X7P2h7gdpTj6l7fjc2xeZgXrC6JNwfhu/LgnK
zUh7jmDvfwoRwOevQMvGESweItd6Gqo0+K69ogsaTAIZ+CMThqU7/ojzvOd1fJvYqYnMYk63TXKo
WLoY/ncG4zmlcjR0qimksM3iQNUOoatbik73HfEKzb94qKsdObMp3Cc43k/sZ1UgF5qRFaZNou8V
Ir8EdwuoGSZxQTEvJKPdV6a0qM3w/Wdj8/KdIw3vkdtPOnJZwyaLrpI1mEt37TYhrPSa88WxUntf
xGFygkvpOSS6wUfOVTGpn0sMyfNMECTXMhWKileuc5cQcoWFRl3xbOpFtI8T/uADOdhHrXpJVAtu
t+agSlYT8+OCAVA5YD3RsSHTAqhyhS4AAvmlrTbHRlru6ocbZdo8qE+/w3UXKAGMGCfzhbwiA7/e
t95VQaD22TN2qpMrqh+/C6qyENB/m8LHchC2kUMqeluiBVCz+xrWwRvpyKg3tjOnwa+3Zh9SyqCL
/qVU4x8nDhNbc+LH201m7NNvB44YcZIpx9HQB99PAh0XYTEO0azRDnEETt3lbSmp+cRkRGV64rsd
MQ+oIe+1kA++FkgeW5DilKysMOF2cIehs+Z9WdFMQ8/2L4VrvcboLqkI1quEJQNUTVXt9WHGTE8i
69+7JNM+r18JXgO65cSfGywPr5tVhegGGuLqrSa8RTthzE6lSoRNH4htodWTI07g0Fhyu7crKljr
GMbctIsdZI7YYl/OZ1nfl85PKxyvP5CoWCmc+RNov53ABEykt8rK5ldjaXcz8Q336ABBLOtgft9x
8TUUNsEqjqIXGaOyV+P4zW9UCX8g3IXhc09scZ3qk4ZhWbnH8Ka1XejEk+1cxAEXT4ensCPfDAH5
SOa+QqbvjqQBIOPi3fLwQK26eB6e2bkf7kvZawK0jAWe435ZUCv15nRZ6q3CV/m+gNkwu4gOW3GX
yLXVBf0AZijxf9qPUFBRHXcJ/bH6f+HefnY/K211CNg7TZTszZ9C3zmjfhDBgDCmhQMky4WZutxw
xwsmNd34CDiznLnpWzK2gkEfJ51D6+7X+o8exqYeZ0oM5jhBAp0ODSdeIcgmvaVCnAM5oJ7m+qrH
yPhK/Ht+TTCHXVB7PtHZfn5NxlRmJHjWS4lY3yf4qdtrUWTPqorvlF2Gu+QNctqZviwH5RFeXUgY
nqh3A4Ln8bzItGBMMCuU188dnH4TmhUrPyeCQO/M9ahY8hkqDMwRA/LUITnj354Gqsls9FAOpVrS
par4xNYGHN4sbm2oNSdRIeP5j7xe381Wdlc44s6+dRBriF5II7/hDjxQpDc1NxGpvrr2AW0iX7sB
+Qho0x4jWjd7rg2NAUWbc0MYzEIZJqZJe2VHtNctEKa6DEe8/Osfty8lLqgRM2Au5ZLLOFra2BLw
a34fGLkHMx80wK3VYvncBjsXWfgeEdar5bSW4ox5FA8KjwFJsNeP2+oVWw8QIbtgi9bN7Qvwa8Fh
eZgyKBvfSKGBhdyH91C+bEi15+qg7KZQ4KxOcoDPlXcMCODcFvyoJs5FMc3XsKqnqyhvj4c9/jOd
uotyju0xyueo+qKPfZ+O05gGBzAEBw4mWKM2tt+clLKKKYGLyO36cUEC0HHl1QBUi6hghIj+JJ7B
2e985FbIwSAlBXR3ZOouiuRCOwMmpeSD9GD6Nee/qSI0fJv6q0wLHVVZH6Qftt2JJevCX0KlJKH2
wLl55w3/NjcDbCtlRL5hZbiFyRqsT1F7Gmz2irazvcpb19LBBUuFcc7Uy4SWpTQ4ihGM7AUiyfwb
mFTMRyouYeJ7rrOptNtXuf1CGYy9OoZ0mnlpLkj4P/eH7d2PuEkzfLaql73ccRXzL3cXaK4aCQ2F
WqGSUb3qJ52Kw09U8FWEwmd29fkaSvLnm7bfxP4PSIAuSSkcTl9igQGvXXGL2B8LwYd3425HrqS8
V7vi4iQMtalMIBRZhJbQcKsTsO3LoIJeK686nYnEezilDE0xSy0/Sol+ObNETYlv5HBuq61e+t9u
yAhswjL1leT58kdr8uE/RpQg6QRascubNjz5Vtb0BBgWDiqo8xjSLoQVuWp64n+pTtw3WtmQLNLA
GKWbyTKOM+/ZX+JCLBQrtcACg9uFHcQe1WbUhON6r0neSLaYL86PRLFU1Dr8w1laY139CcQTb3/t
uEB9QMOpa+IoJ8YSbnDJZtYS/x0D2ieNyonEdild53oE/WGRstCpQCRMvAvjX7bgTQe5DOqXyUfC
G+W2q87TDpAKkYkX2KPS0vTCxdBTCAnegoiQc4tRiGkal6k9dwFNRZeRq0gqIAidkpi6AfmCx7JQ
CTC2Ge9itf+5O8gALEM0ICs2G9hmaJqPIhxSM0lev567y2nMR8fSO5oxQAa+GAh+bnglDQLexAvx
B5BqDJPYUUPP5Yrd4SV25IEnxTsyyj6qdIvHdxgbHDVKxm+g/TnnHksi/wdPswsf6lYuqwHGd0fs
iFi+q20HaFiUKQPTJB4oov5i8MssLn7SAD9ILqm8MLX65wjp2DwLIrCZ5I/07qmxekvlSKUVVNZN
XyUSj0pZXb5R14qVJ/U7zBe/zQGz8eVwOh4v7IWx7m5X+laJcAbmPBUebyYJkcWuTjzd737nmhvI
Q4nhTN6/zmn8oWB+Jdpt/ERvuiHIvJX2CTPQjp179WYsXV4uEEqB6vjN+S/i5ErSnsm4DADpGv1+
N1rCZBb9u6rracGZUeKr17T0DInhSw6XfkZgTk2+4RKGyAgQDD8QCsOLVRdnYbYQ+iCC2B6pe5XO
HiHQKxM0DRkoAMjJ8VhRA3rJMhIxNy8xSgE3ZHMArjFiJ2eRN1PaPZnO7Q/Pdf+F9D70Vuoeu65j
XBneZxfHU1Hkm24IOkacbVQsvIvrwvMyq/w1mrwr3UNdZQDSSe3Ebf1BmcvLfPB2pLqZmLBN9hOG
vNCBTwhUWIlrhRfzRqq/rxFlfySFO6ZRLUYEwQDXc/jjiLqER/eFyB8VDzNQOgPbPjzIpMEsdZPk
Pn6x63IGr5YpZ7xx+6KZxyMUGf3Y9jVWyCC5JtWYlJxMige/1jMdNZ8m3tueue/GkgpybsTDHQeP
gkaWAnmHvRU4tDUdDxzuV71h44X9iC8WFTA1W6k6/pkMAnhU01XkOBOvsDfrqg1w0F7ZXImXQAuK
K7dhdnzWEckB0cU4Tqj8MLmHCUlZEhyNCOtjuX3vdQT63By9rhb0cvTQ5XTI15M0SYJb1XCuXAuX
NmTC5wbMPQi4Ek6CC0v0fwE3byAGo7HwkdEaYQv4KS4jHZ+dOdmJQc2DGEej2a1a8MGO3lMJ9J5M
yUwkxabKTbXe2tEg8hugaqqmzwRhhoS87JRBuDZPVa62oKYZiNdrkVTa8ee3WstFl1waXhRm4Cmd
Xpyeb9cS8BKxIazCyPVPuhgjz2flHTIN2e/qD0+9DjHwRfmbuN99JjR6CGUt3WVQcY+92Fg4weYC
91HGIK+zwSTd/mKty9w6Ptds/l1P5sxEATddhLlFThif/RWNEaKXUsY9ZTzxbWTsxtFUtYuyJz+f
VQiTL0HU8cWmoNKi3ZvkFuTdQsXDr2mZq8Fig/1Ue4JwVw7RjuTPRIRKFMvKiAdA7o2W0fTcKJuJ
zHav49AdADbSUWRyv9oJYeonnOfYV52dOUkyfIuBQ47ax1ryG5U0R+Lgw2OaXS60ZhgIYlBubssg
VWVudWnqoMdt90u+6/seFXM04G8kgUpxP3IsZ2G2/aHUwFHAgnBDKYshUQGI5Jm1wvOnLD8w1V3o
7M2nb1+y3/Vg8UPdXibtTrE+91n/IDHmTj8+6GoJx2npq8+YoPvovKRKqhqWRVsJg37rKb0sp0kE
kfUK11PiG59LPr399w3KzldSaOHWqPEg4THYkNxKFeLc+Y0NADMahfwv+lZx9r6RS/YxihSlDuMk
QK7Mr59RQEG1Hy8GigiTf/2Oo+INNY1EFAUL2ybhJ88GsIUkP3cNH5NjRAEWAJgOeb8qPxbgaoOp
Pt+oLKHuoQpQOgQ1o/NFc7lPrVMVdlniaF927kNtKwRlW/08G+LMDfSL6XGRWS5jZFKYNGE2Zadx
s3KtLmdqmpVvQghGjLEfLnaXpT9/EQjbhYQRgJYwnboU0oC8C3z31HJbqlD5fmVEeHIrQCk5mgFA
0XjlPWVfyOxvXi+w9gn9J01djrbp4yboUE1oM5ZPzst6+0PmSFT2TuDWFN9xhjTW7FS2pwvsNWxD
7Pk1D6NJfsyKMQ2ZMVDdRpccRJqijhX3ZlFLLw74GCx0dHkzttUtkFBLGOv6h4e7K2qDmxZmqufY
lQOhManYtrHtn563DFu6xrKv3AS4CRAqPFS+9fVGVI4XWxaUgA1nVkzBctIv36ioo+VHNiTXHK+F
bAs6PLVyGUR10YlRwhnAjnwxE4WbmlQDbByRAKTYOTRArpfwZVEDArmb11cBU1zamLsM6dSemZCJ
FJMTh8NylRc6HB5SHGLiz9EHiq58HQP9m8piBv/w+YcDlJYv97ssrtCkzXT41GnfWKg11ts3TJ+w
6PPaB/HSuMns7AOM2JM0R9/y2OLvqjFMfRoXx0N4vOA/4ulcGQlIt1u63YCk25VAWerQOAFhpSdF
TBGB+sdi53s/zQpBBgXrnv5tQcanIGDm2eHNskATIP0nj9Br9KAROZFI2cklfGgySJPX08ZlGo+a
YoBAVQHerYt/lQPIlspoPB3Ev2rYrRqhyxcU7uiyyx17no4hDHgeRX6WnBQH/An3a1whE/JnZJhg
7Z/pikBfoQUwBm0IP/lS0aY0bk7k3eW44paz9AadOCqmNjqx67IMb7W3GuBfDlQNjFg808cEoIZo
Cjqm55heKDUsslj5avt74YwPjUB4NNC8ZoxoRfq5Gv/PH9+rDVMd14/DbqYcO5c+9u9J2OqjUqs0
EFgmJ+Pz1xISLb7H6fNe84R/j13m0s1g9OQ4EKA30yBrPlVyJtJ9PjlCUi6tnbTy3Q3zMIJ+MKah
y5eCjKvvkqdJSdJYVQrndAswtXX/xf+LA4ROkApXB2bRjHsbS5FrqogcDAGjTCHOLxwzOMJZIwA0
up7mIoRjCb21Ld5YpYx8mZhlGuWbLSXkdiMMcrbovOgg1rtU8Xj7EQbYGZQYWFDDv+k53Lzw+aUi
6o9BVbZyWMEa3LIpLg0WBDBEmYGMbBSVVnMkRHUFYkruvxFH1aNIDqQR1Pfj6WSux9KTskCi3uBY
3dHT1GXFOAqWRbfKURctw1lSt+9rEQ/1Z+k4t91pzKAfVIjGzlG91fUUcygNOrLCc+4J/cGpVLii
b/Dg3Ux0cI9rpErPOi887ztPT2XUf0ggXeeUE2eZYi1siYPCEY+WmtP433p5ed1lLbWOfgBZyJ3n
uxBITiKtX72Ya0okh1hUPiJpuEocJas/d20cF3xktFYkt8gPNwdGXNixh1/xxC+iIlaqtMrUy8DB
HL8qe6F98uTElDSEboOHdSY7Lx0hDMW+y4py5UlV77c5yZgoM5Z0pv8ev+9wXLmQD0KmII8Ls61U
qiVtjcZR2zVlOiHnPdXEj2n8RqCtvEY/Y9BpDaFlIu8eZTSV22DIvpYjY8RA7+dCVkopDjpQCZwF
MbLHHLdHowsTHHe+gRTV+W2YzOSHXDYoUOtFzgSAdEfvA7/PBZUYoflBZeNwPsTqTUyA2lHXhB9v
wKnQsjyD1N1SqX8xojaYVcESniOiPeBV9xp5BAVGOxvKdWB+6s54cY8Y3z7Vm/XOHOC64ZEDRc6X
pO4yB2yWnQ/djlzb4NzS0/Ml6tbcHp5GZ9FSMxl4E5V7PbhDJvQ7RgEk5QUQgYYU+NV/HNL2uXKQ
+rma9p43of6vUSpZFWCjmw+TmBd/iV6D8AqLos2i0ISyayhrjPvv7oKgmVSiGZcxaj267wodVh1C
GZ6K6UFuxIH+ylEGH/od98efRZZXBuLlPYbQShWvUMa+n/ptu6qaaSi143fluVSgQsHiEkNWNc5R
dXJfsQVtFZlfmkBw0wFgCLMP0EW4vsgEPE7E/Fk2k4vrwqMqH63Uonc7GOL2MxUMfI/gX1lJWJ8m
CcDr9IAuMN5ws1a1ob9yCcBKA+X2mz1221AAk0pyITA++SMo29C3cQmHushCRp/4mq5ySDLK9K7r
2F2UuAF3rFFQuW4HBcTCmCavXqCXCXKw/2e+Cg145ekMAHVSt8WSsbCt5NduMwTa4NMhpsoAGsqP
ZypPBhDwr6K27NTlvMep2ImadEKyt5urVutD3ZthfZUHhPEcCSIl3zn63sC6X19zNKN+RN3f3CBe
6G8zHaOOmQCoSwwwlaJ6c/HV9wM0b4hIh+9YpfLUyG5a1+/u+wHhpF8G0RpUcwpgp3pcWZlBTeBM
DH7LtFF79L+w49/UlDerb09vnHjuu19nfn4c1oXBKGMhOOT7UkTdahU4cZgq0OutkNodFKH7Caui
tLHVIS45AD+0m+dPu5PimG9+jio4W1QfBnnioOhonRSl+FJz6eaZSRM3WboMiS6j/DwdWnIrzSs7
fx+tioUMvhXqMx2AkppX3ThMhkn1TlwEAaazo6P63OkmuCEAo3JwUDH41+V0y6HHD2nB4j5JvD1T
WWMmzogG2PkzvT/S4SEFyaTQVb9BxCoI6c3+2sU4xocW7THaRCXOZMvxI3YH8GKOPNS4VT1Od+Hj
BvIgAOQogCkwtNf0ucKWf0mb1jr9Ea6qUNgruNJoSAkeRC8PY3+sxC5ekCASHoY+1CvDXUY7X+o1
ogddvHYV018g7yOlqeywlGpNU463YHt+qUDFQlQQCwcHDG6rzgk05OkkRE7qcmh7a9VcpLQiBgl+
a3BpQ3ISL8NxDsPf52ByTEtdGkVEozbJt5K0+z3sdXUjcU362FZQQxXlEAQDxvxtBRHvcSN0VDWQ
JPiR56ldJSOlLlmYngIOBfZg9FBvVVvJM83Aa5nw0DZCH1GSpqHMOjF5hCf55uUIfKITqwKzFz4e
iDftL3I+3DDYeNgxLpabZgRisxpY2dTCe+WGIMCAiSYbcE26gnvDK0X6WweoLfso4IxeId+5dEW/
cnibtyKRY8smaJHiHIAzZhWUo/PqjPMBb1DkpEp7BNEgn0Zl2p0q8cFnaa5Yhwg74Iv25ld0Y1Sp
sveFoHRJ7XdCzwr5mIcUwZ7156UCX5ZWHn3r2bM/FjxLLLexDbhl0zQDRqm+iPPmYLCx4J0AS7H/
K6RRlyfG18JwPLQhrbI1A1kPNSWo6v9yRu+pCk4EW5uMnroE32E5J8boLA1vgZ8cvmbSypl1nCNQ
etrSblBfER0etvYUkjPGQJXrzU9cVutVBkOGXPfCE5+OWwG/8aq6a+ISm30tIl0Gn/xHqSayyRSO
l461UbhqUSZJLaVctgMf4CQbA6WErH+wWL2LsPE6ZbvmC9nfNYO5FVTQ2YSGi8uqSDlWQE2+cDse
Bv04woeqXMfuv3B8z0Z1KcmAC+aJkRSMhwpBd25LJt09VD798dJFzXJCdFU7wtXFEzlgWB2I1L31
Fm/fkQgtnDns6w2EpwjaXkMsLUaLQMmCN4SA43O6x7gUZkRzcE5ByV4zE4MpB7OFmlBzewFMfbqT
8YBM2EN9dv7LCHRjDv+FDDy2v7Vk/z/NUKQf2F7GptcnkyJF+tUu/ouowtHLRGTpME9FXLOwUioa
2pJSAcBZZgWjgraZ+uj84X3pvSEwoYmzPQ51TYghJW1izhevaVrptnk6j+cM3rlr4wmnX/YmBdUz
95zijTgOctTnTo46vseVND5s9s9K3UfOf6DqbBIPF2EA1ZCuIeHmuqCmDrGujRDfP3EEFXJtVgR9
FhA2U7u1267ZRcxDaIDXJPPGiMwXrtgDfpcmmyHcd3G6D42bqVpM+XD3BZdKHmzfYFn4uN6Hk4BC
HX3yc9rSjqSunsKc0HsN3x4/M1CfviyTIgWuobRTdXFX5yXyVTEgJ2KOgRdQ6JIUwrx5FLJyb6n1
osiwSthDZuAiUHZPkwYKL0Q7HFDN4fObumUhjweETzKjI4T291w1aKqzemaq78poHTge730JSdgC
PSq5VEaRjoo4ZHh6NeWEcnJF5qm/hRhVoI05ZFSbfOGLnrEeyKKsKus62/zrL+wQxmrZ9i0hBIbm
qaZ6Y4fcyo54gpkcy3XhFSdDWr4EhQ/gsvYE+aJMAXyo4/FCb39lyIUmiqDhIeyIKAmql6db4Gnv
wXj0/UpJojGgghiyPvhmXzp1G16WfovWD1MhDlOFLCi1idIQIzaV82B+WzzJ4lZhXd0J4yd0GD90
YSvp+6RAR8eYEx/UiR5xCKPAK44XDzVVFsp1V7MW0IE+Py0UAEmpoYzaDwVRNW4Pd0TyGhthhr2d
pA809dmdJdghjwdG/65kOv2zicTT/6aTS/lV1mW3W/uDaA7/LgPtK2Yq5R+Zw4A1zYfylHAJRQvL
JFg460AtiUDDe1xn0PIPF/+YMegziekt8DFWPKmVs4vwCglDdnbPKYpXp5ObbguPpMBdMcVVaqH7
qHZS1c7x0WkaD0t78biRNHuRcooQKLMx+D/jZ2ltD7qRE62jmwI+qNUxSZKTkf3j0Kz4LmkoKbky
kmPLwk1vyvwRE3hUDNo7eUjLLHY960kG9pUfVMWAZPFMHYWTnmGvGz71StSSnrvq61bgp9yBw79B
GhAyMlAKvE4bxgUEur2BC7FvlJHtc5CI3nDm7K2m8xYqg/GUo2kMl1xkVDXW2khL2jIs2v4t0mXa
uf5snEjVDPci+GtsDBzVIKWxCCNJudfAbpQx1udiOwdRQID2qO97RMFESpVAVemXuwUH1JT0Zgdt
dqvoWBDA5HffR1KTfNT4TMcu4tU7yfCXtXK3EUAp1hYNJfyqHyUEfM+TCxBzTMFEbus/d3PL7mT6
/afLVrxNH8b85DI8DhZwJci0K0ny699uoqYdCdcgTZk+jRMPIEAhUWiY8a8II5dVdOh70JdNuakd
F5OzwMGIYeG7hKgNI0OkwRzpIuElg0xQzGLMzNgHBFyo1Kuk12V6Myyq2M6l7L/Fk2VEy8IXs1Y4
Y0TngbAAbZZfFCOkm92r4QNgNdyVYp2Z/T/pqwGh7qhtY2siBUP25kwsn2xVbpPxhh8ixXXIMhzj
CsLeZXaDs7k/47R/8zeMTzoy8OHOFNhJJhgo4NUrO/VO4JV5zKPEe1G5QSoxKAhKeJzxt1+dlHF4
paOhzciSkY3EZqQNErWWV37VWzPmyN1/UHnV6HvrXleUNPymWCycb0ht+Sj5SZAklj7+M+0Qv4OA
pq1qBsMoV3RxeT5ZZCSM9nBuskcOK0yMLJUbY+hvgKT2xn8SE/hd3e/CLpTLHw4/73YBOuXTpQus
6Np+wY2tS/qSqi/ADtd1OFefX9tprXHk/Fx+wl0iK2Cex8JA5S4gapIrZ7T8A1BUm0jP9kdGmlRy
YPDMEhpRZt1G9fWH5mcmJhRpas8MsGznBU5izSveIO5sHceH6HRaw4QQW1PWIEqjypN+T6yMPrEB
gmqw9LT+1cQFNTQVUbg5AtPu7Vg2h5jge01lGvi+4xWe9kVRj5GvzPDzXg2QK1yK0xtpTS24fvIU
tmu6KHxVw/bqihGG7nyYU96HTqNoHuIuuFm3H5W3QxxXETi8dMQ0sJbowm3gmRt+cMPDrH10FbM9
Oc36b+wbUAg/AiVTuJjlb0wcUs5nq5y4ljPiPBEd4dC29VBfmDYND9mDxDLwZU36Uzaut778M5er
KSHRdNiN2beOe/uvOMMgO6xN124J3S6MlAUoOE/d6HJ+4fiLh3bXGtcc4+vwvhEfL4nNBmbgpGcY
DA8QhUD7+t862fX3RZAzcRgANi872r1kOSm4ko+l5CB1Jye4PWHishGCLnvs+8UiBW5bU4EQK4yV
P/bHNBA+EbOSBZJLgB2wj0gJ9Xxjm7yxqnFmxmInzpllDuO3l8LsxcAEtboyqDegOyct/S1JVpTb
i9y5szX9zVW48pX/UIA8TIszhBs/W4EXibhALdK2utEOnOc/lG//tIbDlVztCJIxFQG4gExyKoGn
2FB9kgZ0LJ6DyT/U1nzesFum43mY1O626vfcBmLqN4YJ1P7fMkbELE6ClRvYmrf+xIvzEX6uoLlG
OUviSYja8jRoMyYtr4ET70VV858gD9hpBBzGpTSWVHnzb7u0tbwUGes5B7lNGQkq+MWqp38MzWQ9
ykADH1PoDGlu8AL0TsT3Tf8chmJA3QeV7wyK+nKhsxgK0oGJUPpg28IQ+8ACy+pS3/MSXBQdAfkR
gG6WytgNsgabRM0Zrq/iVhA7n/KzSOFPkrwml0CVlAMPOAqDmfOQOeMQAvd8XiCqXw0fvBKhDVb2
3P3zcSfe2SW5o+iBI7HT1jQ3MxwrxHM3iOrpQmZYY567htIggvdRyfCZhW2d837nhPKtyBc7Ujho
Qk6IM3szzlUIafOWckAkXSnjAqhumiV7SOslfAmtiMuM6Bzvnq+Woz2QQAlZfNu8pPgpgKsvwXLJ
Rrjiz0MFhvv6rjwnsTZleFUYY/1AnCS0bSEKcvvonvOKlz9mLkQvIr8rRz/2v7GrZcRI8OmyMwv3
1waE4raV1wmgZeOrv/Fl6lsGNViz0MzTzAdYzfY9gAyYOYy2gzxmOgXRcSlOf2Dg5lcEOvNUaeOo
smba4UkB2qfmWvxzsL9gFGMOJalQkSuJTpv5oYwhc2583t0PcXESBJSkuzQNbbI3A1YXd3J5gh/F
FC5V8NRG53X6JzF3n8IcBA8GyYrUb6lP7rGPTq9VypN1z6ubdaZaTS9nSIiC96HToOCRdbmu3M6Q
aI6f5H7/URuUctMi67ZRJJfiySHs2qBME2JQKZO35bcil24/vt40oflEMTNbROdtrJc8R4ORMFh3
gqBAIObm9ExXSn1RKmY3MOqYdpBxV/P+yfO+YGuOp/JGpk2kQhZyAJS56nInJ95ZI/p3iMzMV5yS
pxD+Mq5e7Vr23VWeiV9nqF1WubtMCYPYNZYUICpO0Y7SSj3EiI/HhSRikdmjXBFXrLNiIXPb51Kb
6NIYAvBUid27HjBs91XjdJh9+J+DDr/z31dZqcPbH9ejKVYlmghaL3zlL/0G3L4pdWCMhUSaKPT8
I9IdpiAB1eHu4KNbccyT/KRddcnXouTOTx2Of33CMfFMuXqdRDMSqaMu399VJcfgsbRM24cidnCN
7ZOhTqT9Jo1y3qKKW76eJLU4znnWevVmkRy0phuqiZPTBf80S/s40ehrlpWo3nEs3An463DS8Q8k
gl4quM97hQV/1VYHuwrE/8Mtn4x4lmo7n7D2jHHWWoR7CY4XiBcdEAjXB+YXQ9RhLHql6OTgscLb
fG3LyHwRNHQnb2g4SNWGEILDrgcP+Y/B96NEMVGL+q9jCWyldIGhtqsGzh3hXV58eeoPMrbIuA30
ltWlPoWnyRTa0coci7//W6VWLaLZzDfoGJfzHx6KkdQbqRjJ3hi1ZuPKrgSQpMJ/wAPBVzewXzb3
EXvUpvyXyPU0fQyERGQiVrSWxVwL8z+e623NgIwsGII2f2qx65M74RXmm9K7FRjNT0bQMemUfB4l
Haax+uz0CxYLVShADMhT/NHMX7mfk/UZyj1HO0MrZ8OMSfMHqKJswc+Mo3ICOSGSCcMBZDGe2slk
9P0LzO2HQzt4MUydQr8bhlZK5bH7yyR5cllV41axm7FsSwj4o/or0Ket2M4PDiBo6UU4LQGL2mv3
X6NZHGWJLRoxiPoRPEU9Q3s3rcvgaig6Ym+gGpEb5gkyPtejF4Jhamjs8xS9TXsVpeNFtEhM4+7b
6bkUuX0ZZ9xJL+Rj1Fa2lrqeuFE1lMpqMcsiSnX9VR2aoi9uXcczC8OZhqt2vGSKGH73Ggh2amqe
e7crq9FsRMlCPgVkVyTjCF88RgWiWJUQ4e7kAoTBCGPj8wDy4g+R9vIndVNt8ZsawfdzWaUOiaL1
x08OwKStWWvU5dFl3VuLKrXUVv0x7N8eF9zKlqXMCNq1Dzx0/q5GkjkYpr0o9kNb2+4ouiuaE+rD
IbfyA5sPrCucu3Kqr1E/Z92XMw5DYyTR9qQLhKa9533R2IpOcIplZfVmpwzf8M9gopJlFgFU/pRA
IHk6Srvb/U9aY1ETKO+JcdKtydndsvBBSIgi70c5k+MskoEMALXaAz79Cl9zpwnkAZKyId1NnWxR
9Yev/h80K/2YAV+Oi5H8WSWS8wScVSgAdCkYJjWMK+DGE6MBwYxFVGPeew48gE0/FxTjifWFo84S
MbDpbpg7ddGqSFDGKz/U2GOObQt3vG2dMeYiZ3JAXse5YuCQArUy1b0dbx+aCm4Y6/B8oPVTY3Hp
uN4P7q5laweK/HVX0do03y4Ap4TQWiuUqczOM9nRvrKbrpeZ8dZW+RXM8t2zYAa0yR4g73Bwudxm
6ikTkGyz59wXnTd6BfFsgcSnf2fkwfs//gPP9WlJI/wn3RkJir3nzpeSTCMs69dz2jKigpIBXaj5
in1FAvG7gU62ur8EA7fZ2w2n5SySd4sHaWJiyDYBBT0MiS5h+IaLtfNQWqmg17dfwLHjt7BrsOtn
BPaJ1h2Jh5+fheQ7MayQcQw+YzS066+FDkEs7EhcKt++IjXQ6I4IE0W7e7dpTFp9PAMn5NcsCXE0
iInipdJbjMTy42NTBeh8KadZXITOYGldoMla3Va7eUynlW3X6v9EuraRg4ECwjIQQQ9rKscJx/xo
R5ymbml3j2Q1wUKdCDQYga1XoTYFDaFhojlMHnhgK5aWfnws6E7KwKeyJU/iP2CjHneK0dUIiGRm
1QMHYaERzaRpvjNPjiuTi0fdoZ54KMcsbHKgPU7jQxN9zXaoiLJ8rMkczWwLgPTN/TC97bzO/s9M
2JL16gNVa/1/naOgbuuFOgIIYJE1OWfRQCGA6CmqiM+ch+NtKoIserD+y7t/n8lqBLFZ1uEoxGMw
SM7pyLMJL7TvlFHQirRXuKNJw13zU90pSgMpKQDkDvbf54slJnTmvmEUPLS6J2oufhGugSJIqZDm
H1llVA6dZm3Pfw/wHQ3mBfqc5B7ci18bgh/uIjpqPJg0liwj9/v6MXtURts+dYx/D6uAn7iyWbIA
cnEd6iIkUYeXcIc9tIJCTZ7Vyqs5B92Z7+jkNJCAZUcMACSP9fHtZcdlrDvKLpUHDFC0yNY6ZzDC
sdHkaCLBWHMVFmd3UlcZDPhCz63G33AzKJPJeCZg3GuZvnq+IhmpJUDaiOz8kwmK+2tToK0gziU6
PArb1ahX8PN9uY7sKRFFx7Zf4C1iryL3NQtVGt4MdTtlDoDEvalh5Y3gUIosoLBFTGNYIxoVgEjt
mPUzzBdYNXEq3vUKsLkVNaaQMOtSjCY8IJ/0NRdAqdZu7qJXD7FLxX01SuDR8cwuLZvG+Hnt3vem
QdGj3sFX23xv3zbLq+U+qtH3DbkD6P5vYICiO0jT6wEf+BKjMrGnI/APrA9vXWMe/rqUl5DTLfLO
TeugsHBnr3tZUk/3Y4Vo4HFLWQ91bmYKx1urkTB/nVQPFAiz/VOAWY8Yxq8xMaXfILioGuOdI1zB
5HESHClzC0fVyX17wlF/p8ljyUfdTGVNoFidvJVj3/8ms7aCI4JAXr2pl1JqolVlEamk3S4Kw9jj
pZqlKgj3xWTA2+hGhUzHd++Q40M/K0H3gCET1Mmw847yfTMEtZCLsuSXRptY02VP2ldNj7RB60Zs
v9hnYMMc1tuGJGRdjpjZA2IVIuvGmBr8Z5u7/GIAvHusY5oyE/9aOQGppvz6cZQlk6tM2t4fjIAK
Pc1xESU4r0fuL43NgpEg7rC0+5P2lUKj4+uk+o3damleyHl8yfyA1ufrAtQTcZRSqtpstmtEF2IW
FAsdop5tkXHqumIy6hgkziD3u67dr0w/yoUMdetxJd87tWuVBy0CcaF1WbtuDs/6I8WdNhLjLsvt
RhBq2232yAgZJuV4NzH+hg2WE2aRHFIOTUg16plGIIeJAo6SPzZcnarpqu4CBHLs//Ln3wbrxzh5
x87mgoGM0TJZ4Rhl64CzBN6OmMFRwBkYViw3N+ukyLzr3hHVK2h2lNGPBA/tagA3PPUXXfNYKKEk
Vui+5r5hgK3PmxCy1ArH2IcVApwgBgPBWMhfwphVXLzQtO9BIvo9+ZfsvWSFViXC6GdxYn3Nhq24
nQu5T14XY/Aq9DcJbYASvfcD3GV2OAv3ko4RCdfJK0bAo17AVEJ6XdDdjbhd9DAauIeyiL15wJMT
+/RLQ1D5+51si1d0sJf6vV/gLre/Afre8Hlllfpk8Nm2+TqnGRI4wmlz6swfs7UOZZFYAvMXlP+E
NMmkgM5gKzC2yccFc5dBD4qruo8SXx0emQ1R2kHfvoMxY40is4PydO1GvVJVnWoeiWK7RX8mbG3V
2D/1fr6p6npI7IYJLXAe1kEjoJIbNDY39hByY+x+LOLp/Cy2+7OwYUPXovx3Nj/7s9RYg1vW3/96
5DQ+RYUmBhEOdS7yanoZ2ioqTiVO1iRYh3tT9NwYlOoaUWaDP8fpJoNs9jNdIaZ8bCBfz767a9RH
TUpWSNnkIVs+6lUU2u4U8aptyuulL/3yzfs5K2SN4yJ1lWYUeK8YaSrkfOQT0D2Vlv5VPNPEeQto
6lVSJDQsR58fMo3iTcOiEFbmB3/KerPUriMwxZc44SXjS9LsKZ4G8/c9d6We9j0hMqGZf8Ss3lqs
VM4CopK0TmZL315t53JWPvdRBk1L0nTdmK8A++scnQ0GyJtAy1ofYkispTFCZocjtJj3rZPRq1rO
G4EUXWk/yTnpq690EXfAYfVGj5BU95FjNaX4b/1PrYyd5/LyCyqg8TDq4lJfdklveqDYiPcmpN1j
PdP2kQXpNAr9IKYvnzIODoUl4HOjPfJfByuwOBPSJ9fCHK536WnKfG3JmlvdOpSHWTMI07uk0KZa
13q5+Vj+E3DCc5560FIkZZ7PmBK3S0/vUehF4rvspYiRsuqrdaIyoSRr+m4EPBV7DHyZWAuKXdlR
nzk02fGQ3DeD84coxWJCwJ/WAWJN/e5EJ94ZIrJYKQ/JYl7HS8UEgF78SR2PIUxfwy08EBijBX1z
B2e8lnwLxteuvebwQIlyecAx6l3h0gw+x4jjiF35S0KKERzC3JraIBFU/AiIL//RDXriqxWhorZa
Yhg/ChSIcLrEH0a1xULTXD3TRgNyKPwqzjvRtQUeN8RfI2VLfb0gUswt4PFOqZHVoDjrGIpcblEW
tE19UOPuBoWH6evIiscP3GRBFeJzh+BnBZBAg81uMY6VcLhpky8in1JpkcBlFuauU/Fy2cCN1x4/
lqe7ABTvTgekSMg7MXRM8m1tx3Ubl51CP6b7+EFMT0qfZqEG6szWI2Z4qI+vkrEEle0cxwfKXxXm
dV1CHJQKOSP87oU7I4CRhmw+6xD4dQ8qaE+LmTFfaOua6XwVjwPfpEz2aHUi6AoJ4wstRxIMdkV4
UP7RIcZcPdP4xXjPovbv4nVcybppm4t6qfFil4a+PCEwWzesUgNzBJWmycyhEE9AML3POkLDoIkr
Le0wBvdauzR8LOGnQ8IsUkQ/ReLEADXCxy+Eu6dFHtiO6bObP/QCQT7fWkM8kR5u7RsekW1S0sW1
2qEFgexD68jORhduGWdTQv8P4iSRqQJalKlEhlA+mj1c/96apIhRCuHcOQrV/53Yj9la/jItSv9j
QBuF9odUC/+E8hbR2/vi//TibgIfyXj3yPlpKELxBMAU8dFjamdg7mCXApZ8LmDkgI5BdUzHZEdo
JUEApNk2PEteDEJFLVeS6IBikNn4CNbxHriWzy7vWcwBo0I7ENskqfsTRsyNacEw/UjSrHfW2hua
UouQyWaZn6ACAxiJg5BFx6fJPDfIoDM4CwdBijNJrZ+jLW1fHmw0Hai+3/vGchk8UuaoeSIEyYCr
hqJqqQPFvDi6LYxPJkXUV9EIvk5Hu0AA14MCE2FTkAUO63V45p2g/L9isocggTvELVIvdrLlfYsO
NuLov/KaZnAeiOj3bJ+gnbC3Up3WSlFz7eWf5aAdSjCBoCSj3GqfwbjYZA3w1uYx1/tcWLyTIQkm
xBd2av8X+TP2rTw0zU9Krq2tFGP1mmwdVCMY5JcaiG+/yhQR0fYViWt0DwdC2bsTO8w3+k6P7Tan
RLDS7ImvxR9oXlLkZl/qJqCcZJOc3SPrkVXpE0bkkav8NTHzmuEbsEQEAerfBpDwhAQI7IG1jDBj
HKvG/ZrNxUnbK9waWei02daIHCaoueDSHNWPW44Yt13InQUdBGvYMYqtBc+OB7Mc8pm2WVYwRnbk
guBCvFP+rZWx7ExBg1qRAzBxPwps1ceyRbg3xYE+gEZclEhod42J26snN6MDRq0ktrd1aiYCuNs5
yUONqyikl8P9ZDz7XCq03uXw8r4aKj1XkALR9xaDPwE4rSvb7OQt15QwvRFgCp2Mv55AHKzjlH7P
nx8Fm9nCxN4/cM9WMHWYBopPCzeuw8hA6hzy48hAVDrp3ceWRQ+gPT+bQE43gNNs0Q6kegyu2Wcg
esY/gI0WyW5XmxdXGIljaIP+med12k6zQaR+Pq8VxEpp4yGKyqKIKkFz4t4axUGFYHIusBV02Rwa
I+yIi6px9uy0SB5cSnm1anAz7iw0wXxZ/9wqjek0U9s6PkjPT7v/uy7WK7j3wEwA5XbU+1+c+vCE
S+rD8yXnI6eQ6BKR/BZ+zQt2ay3xn9a25UkAhKynXo+1ZJ6ZdGeaFqCubGuc1wFWUSPa1IKbt53T
y5AcqAqmrByHQ8r4BswfBNwEvu6Tu/5n6/OcjRcKafD+e9Ll2js5D0X8s43MOfInxIaXCmapQJa1
mKMQWKba99R0avYn7NTAsjEDy0wrZXoQ1EVH19lfhrIBuHwTFXWKMY1vbt1or8zq8HAnAb6bIw32
UMM8x1aV5ozd1fD0jxQk5Z1m7fn1n85yzZGV3XU8ktIs4I/PwPjlZxaM0u/3sDvjEyMglRl6Nen5
umOsidEPab766cHK9vN067sOWBNN1aOnRChaxsvWqxk6UQ2M1Lh7b1e0nrmEZrMa1B3GK7d+sDjq
tZg5PaTH35yGVQqWErLj0eLPj23bnPS1C2rRrDPlvPpq7pI3qO1Vfadl9Dff64H5H2L2I4YxWUZU
VeL5AavjkSC7E/O4oRHVG/S+qWfOWwTpaSg5nGDJsDNdWbDIfUocWosfPDhUzmwRLzsbueeLpAdE
/mdQNh9Oy81eJKBORrK/9NZQs2XHe9NcTCEoQkNf2Qi6QdEYIC81xCuyaRZTrbLlCkVWqKsnaYRg
Qco8XdHrOJw6l1IjyjmddIKIkhPmtNR4wR7b1AyWmyT67v5QbnqPxg9GR2eQ65EnC6ksGPni4fez
avybYSf3tLu0ntOwwuVeOLgsy1nxBFhCXfjRR4gpFy12UFXmkqBl3dfBxeNBSomrNAHatDj/RfT6
vxjyORbLrwUURV3xea7mptrDvQZ4pu+qCIxV57K4RO7dpXfXR09ZskafnfEvwlETJGuf+fSWHqrw
BKOvFI7DMU1rQMgPP3P41wzRH0daUWDPCCU/SNIL5Qu3FrSnmvdqTFkrRAvpoetUNlxaF3qUsZ+7
45482kIm8Wn2SZKdi5H5Wpvts5aqQgIxqghGuUCxlk8r7U+A7axg9IpQUOoMZcCKFwZCrotiZ047
zTNPwpXxEmkvirQxj1Kd11sBDEWJUe+zvDV0rnhs3ponFr7ZBRpJOPNLkXzMOiPUDGywl8L1nuJ/
yFSm2uHrGHc8XrzVt+V+sHv+Fy54eq3C4X4zgyuLiF9bjosob2/4rdmKEh7O4iY5WCQcUBTOvEHj
l/DrAbKm3IcTBBLI5Ha1JygexBFEo0dn576EizolGP5UFypK0TVzyDQiBmTVYNbI/5eHrIskKhKH
6vHxwUSin8QHMBkihXsFlKOpMtwciWIVV8INZLNAQ2CafBTuT2WJqSdyHm5qouG9SJj1FwE1G+m0
li01mp5shLXRQMRYlOllNfY39NBr1FvPqpLwQGc3QmA/gWONIeagQsBe8riEb4JZL40Yi7pGclIL
sHN6IlfWhipTutonLQuPfc7GSIZGwwJABtejyv+DugD4ZXnBXQ6L0RA6EF41JNHKP3oMPnjNCo0B
3Utww4/Ko1Sts+aW8P7mN/CgYakFzytvlVnI09u49gtuD1EvTEC2+R/+esRsZW7ikQxISmuTxgcG
huupzt1Zh3k9jED78OsCsjKRGDksdSUR62J5+WXrAOY9igC0KwSmsNE+qJ0zqplduHH6aiZRqVME
mp/R0OtbY9H6vWE3qHQqHVj84HdMpOjysNcxZfQpsccODBWuO6aY22KNCwzthH9UjsrwlIw/awUO
UtkHZLSOBAt7AOQYjLza8GAC44bvU7cu7YcZ6jlLP+kVXLrqJVpo96NLGP3XKQBD6t4Gpdmenhww
1VDWnqOgL4ya/Ui1/OzE4Po6U4dav4CvDdLqcYvrdIfDrkENbFpr0IoIs65/TOrr2U3SF2oU/hKn
ioZF5hBggNM5Nv6l6Slvu85vEmgMXu1Anyd2NtD0hQVbAxxltEHs7IbSm78wnaV3MqaZAX4xwm6u
7ggyjzLgvTh5j+5t9E4snizrMlbQr9iWyqEEAaElNuMmnGccuF7QaGceGvR2h6DxjNwVr41AUXbe
UL59rUo/8M79qwcndCb6FsD3KlV0hPkMavkMtX5dW3+YWQTJpc9Ekily96TTxrcbMFpvm4kp9wrD
tnc/K+vhV6/qJhYjzWRLNeAJqeHjY9jRXn1SyecDuYDWLe+pkGyZO/q5N3CirK/ZSl2b6Ch548TR
s+dtZxrLSLcYYXNIK3Yx10o9qH78wAgBo9HyN4UzDQsrRdFkJR1vVU+2aoMZcSCPuWMB0l1L/15n
iHhI0Jp69wfgF5aPASskQk3jOAwdENJadGnjJGC0mYMtOxefXqVNtG0QS5Xug+KJzjlYRljEtWZR
adV3G9WLYsDUzGthh1PeZ37tjpt+f+w+BjntoTFSjxSCnuQSuw4l8e2OkxmoqrlVn8oS1zABa84h
sIKhfHi81TcmyM9H0rZAUGRxaw4TrRbI75gugCJSXYjb0MBNiyiLzLov7U7bzS0D0DsDinvesrvD
Iga+zsfh/sCyjY2mQ02xEeDp4f3YAcIG+SaE5M0Viv7Be736jsj1Be2VWuaDXfQafSuKbKBHfBEa
0oI76Jy7XH65bJbFl1QGqLu/WWvFY40lEs9nx9oQi0HxP3lC6yTqyMtNcetNeXLEDL2oyBV9nLqz
y5hWhdoJQjTCH/BCjsPfZH6iiBN8rpEa89bNxrYLSTeFWP1aJQrg6wBr/GNU2n6/XMsgy2MAIb+y
mNHpyRvj/Zh7B8KTYGQKqmSOeVo8vVAxKwGIR/HD2v4Cmi632C8+O9CapChQyyguQd05qe2iutks
7+caF7pBj7tLMbEqSfVwmj+JT/wOS1NnGlGeeSnUz5jJBOLinGjrVhG2YsEiPeW1OOgxdrbWZ3tA
A+1ZT3I1pHHJxuaH5a20uw2uT4h4uMfu8578YC1A3rvRflhYjHACASpVME1zAJcfpJYUepz2EnS8
qtmWipEtcy7LDmZCg/8Ze2rk66hOV/Wts7qE4zciXY5Bt8zxLOlj+99IZb9PhvhO5f+mbFOS/nRW
ewP3cADaUIJQENdKgotY1A4kJwwDkLg/OEaeGt7hqCHzGvhR1YmzUNZelsTmCcrrJ+zbQd04LIxA
8YZP6nCinZb3jnNnG/3zu4G6p7940aK34gYipv06vJhv3X1IgrcpzWCFXPHuUAwhEgHq0PxgIO+2
9PE1yrEmaTuUuVDxu4sJkRyrT28zYzs/l1tLnDvP6ykH/4LmgYTzNWYekPv7CrlMdubDFoHP1gRu
ftdLeu38rXXVqw1JlNNfR2gu1yyXfBR0bsl6KhHeNc4vc1O+jSAFTK9ACliPOIx/R0uQ3UKE7J/X
X0aTgLWQ5MUWZURZ7hnwB+q9f33KvAb9xwGAjJxTQH2lK4NQR9Vb/DyjAGKgOVGyoC2KHEi22yEX
j+7prOCGKW1KGBI5TOcYPpRwm9vP7Y0VCtrSPKr75wj3k8QduXr2k+ke3eb62CDGmO3cc1fZHG1V
r2GCnMPEJaJh9lgCFCIZKQtvAQy7RykDdFdIjk3MSX/dbemOyfOlj36UTdjRdU9/T7BV7HFyxoe+
XnqK0hnV9tLDQqb762RnJk8izbfH0orq9gSRsoeIc15ozZIK/gC709RZxdgoTLBiJb0A2BW6lDB7
yh/k4idRktY7eCS7zMUvoPhRmEFRi0viZu1cGcIsqGUUUzi8yNo+KKvuY+pjiu4XLBqKZyPBaNwG
jl0Uj8yZsv+yQNGL6tFOdGPPZxIzj9cnj98RasnPNDJrrZjumIF/u2ZeNStBj0pqMLxUXOSS45LT
VT+njXcS8L7zRZY8fLLU7V568I/yS/UjtORTO7qb2B12CX1L3UrBZVEq4xcvK2MvHOp2rTQENAoI
CZBqZrm9emt5e7sqNy/v7nWqzJfs6F6Gmmb0OQmPvBNugl11FcDyZlbiuqZRP+Gte1cxxGQhqpFX
u/ksbp1Up45bFCHLVqkN5+ipYwORd3I+ZiEySD21Y+e42Z6yjTMlBP5WUI6P4ITFKSkBtXfW0xW5
vd8LLZ9B1b8w41bvg411vZWTtyW3GUyswapHnakJhWDmqep18/zSs4Ip66SETPoQYOlKe4WdojuH
LsC+SPwLXA+tRwiI4Qk0Ygs/iE3CDalKxXuEQ6/kRVhMzYwSTJPGoyvh6+IOYZVR6oE/MVgH3927
QdplVF/sP23DaffF4UvGDoSkONZfVFRRM06j6Be1jjEdnXUEPPws1PlHT3swIZ9QDcG6X7jegRai
v/LFyP/1M4ubrfEwflQ7+hVrWvHSKXRGpS+s1fdWqX28pfhj1zas0z+sZZmUJON9WEqhWh/6vvWN
T6OpB/XVYGA/UkadPc0dQ8GTUovKTzB7eQ49Tae2VDSGElK5Q7Iwvyv928QfgcB2YXpmrHLJ2XdU
Gmxfh9VFeWmPpbqvX+ebBQVjC+qlaW9SNIKxOY2hT7d4tLx+5j4vyMAIpS2zAXj7jaFhFDpoU4FW
JmKq2sgsoiTyssAeY/UvSGWcXoLT+Yg+V4yF0f3Wc71kFh98UUDzJ5O3IPZmjsiWhNqPvpr/tvor
Stm5QvfOUmXoRpCrSwMlaZtSG7v+L57M4c6VuwUZKdZnadT0r2crK4E4hbFZMRwuzB4pQsxY6990
SC8GAz9VtG9AtGUhsgZtkgeHEuHw+1uLQ0yPlaUqJ3vgkyxvqweWXbPad2pJToU4tY37pM+Yj0AL
9VA21FlOQki9+vofj/WO9bMTvUQrYlXmizoA/ljDGuYwcnUHhZLRGN3C5iTwmRuyLW2PidlEMTpv
VMWTyxKsQBJLFHv+JZfWgT1y+AF5hlcjVP9EweKTJJAmC43OPk2yK/HXABkBcIMObiJjPH9oT/PG
J6hKdZU8ODtHA3//1XGsg1PPjhuEJnL3IIMGvgbB99f86982Dk0+t6HNUUrKx8ICGVBSGhEteneE
VLIE9olOUlXRp1+0mqwB7kPDcKfXYqt4M7ABwfRcdnbWKae9nMKoqno2eUX6YfHWpEG24mx4ILel
UwU2tofZGnzZr0hXEQc7xMpnaBmszRPdkDEkZ/XqTHtFTv2lsKEMeJKg/+s+Bmj2zSXQ9OaYIwDA
S0AhCVW9LFMipH15gnSzihD8a0eGAWokIF7RUB2HNODJpqGqgbWzzRv0662I8yZWNN4sDaCso6lN
Q7KkUOSJeQhNp8xYsunsOtJQF1dFgscnKPDm3Nui11r7RQR5Qb9RTN8hXXeaBAevJ1Z2Zttr9wfj
BdHfby1d26Ns+U/+dfBB8gB89U7dzqfCn33woCL/CC6yq8El/rXohkKrst1fVwyADeOM9zOvivhj
UDU9pW80g29jlSVewO1k4mInuctSKzAeFDzbjrxHExidFJRiCEiH2yLVetdCq5Cuid3Wd3krIVml
BvK37BnY7ZTkjGR4Wl5cDbd2B7zD6kSGmSBGuCBTkQ7rJUbfOBbxbbXBjcK/+7Xs/XJbwBv8nrdh
UCBeDaF5laSgazkRPjnjd/8QNopJCOSr7Bnz6MLOrX3+OjKUzMeR1wqr4nVmz2iiVV1YU0rt/7Ip
DJHS4Bi7X65XZrny5OZPGKoQP8OvOHBA+L4nMMO3D6mtj536fePX3+FnmwzYk/5YQQl/fFwBFt1i
R6pjZGTdT+m9t27xo8HOKm7/sA8m+rnsvYaAKA4Thu/frbopelBbiq7QNhrvoE5WFuWRu4sLkneW
HoWl19tTSC0gHST90XXCYhxUeIaHWtkGT7Qr0U3TQsObSPkk9mRjOkTrel38GTeSd8Fsyis6vV2k
BDymSvO+jZ5H3geUkQGPwoc6oBJ7P/d4l7E0UBLFWvXym71uRO/K7XU2Laa0aW/V0rkD3qvxmdu8
G3rDjdZ5j1W2hOnt/vMY+8XiovcI8a5n+KTvtjU/5j9VC9DOYPYwjLe9rEOlaXvAUp6UUQvCm2Gg
h8cz0/uggT/bK1986+T4HhPKYhxkqNj/RM2+TmqNj1jq7IMfXySVUL6JaVTaNXb/YToswMZllWZr
SuSXtKZgUqddCi9BKrYarJbO30+OEmZU4ywnlCXyoYu3CNdntwaDsYyQ2qLXQyzeUF7yEWIGJjSi
wgs00rYyxk/pzfhVj3oEw+jNSHkbo61O8CoZH4pURlMiFIBbJCEK2bkiRSu0dVwjCtpPg1KQuOMa
ZZkx3zCO8JQlqGjIhOtPnWf/fmKJijbaGP3A0ZXgAyWgf9YbEptHXQ8BRBtaIIlOmUnT6OekQkrF
GdULcur8a+dGnqkq6VFHR5dr8VRP2kATdl0M4h4VrY6R7iphPa50dyenxPGRSup4/wBJZ9GMoTcf
QHvQSxGQ5MTuTooTuw7D3s47Hwuo52F9GRezfGxSCWV2zd9KlRtN2MXaOajNfZraCKlB2eKzXR+Q
romZCnJPpsKGAEUpA9YHB3lINEJSKsH4/blRtg+sYbL7jFpbicxv9ivIklvW5svBa6Z8EHGRKqqJ
u3gOWwaPw+a3w0cRzkFXrsSDjygZ7Q9avtGOnt6Apa09HaEuBIlM3LxZVfHnFSviHfHs9vnL89Nk
jZNXR7KF0ogVJXt7GVh/3j+x5vsoWDqqHcyZXZuCBjhmxAagc6aWJifb6H0bzH+C83THskaFyO4Z
uZNsVfqjYJv8FG3KCJthkITLNddnBh3qDCB/OeaCUwUtBfuZCbXeO2KZrZV289UzDQySiui6KcZJ
+yZWGxef1FMCXhJtUD1UllifsFVTTNolpbNzTaxo7zqJlKygGMFjnRz/LN/uvuILyIdXlJ/6woJ1
DM9IgfhcK4qab9WVxyfAWmlGaBObNUwL56QeqR2zadp5oEtnRYYUyK+NOFvQeKOVRZJMziwJVWLl
bhAPjPac1r/Cl0QnDVKzAeYMrYOS2O+TRqXUhehtvpNScClOllC5jH2T11pnzw4TEKeOijHy8Nge
dJdHOVzcNu4DM6dtq2QZFR97fbwudwV0GcSrBRUWhyhcC8AzCtTEYBnOXmuoxnR+yN9BDpWwKoMi
GDZiRAPScOm9U2lOwDQSqZ3fV1a2TqJYPCILkFXWmmc0D+0jWq0x8OaKr2C8xXHS72mxCdZATour
0yvv4OOsUoOcoOgf1maSk8ALaIURr7eK0Fo6rZ23ie3xwvn1fE01oXlUTHVH98JT83BlWDa+TXZn
q9z5AsHJNRFzzl/k2mUw7t217dxnNy2FiVEkLR0iWlZ4AQC9IEcCx6RsxknQaITXh0iXCXY8xv38
A2Om+ylQn6VZQJnsvq3uhTS5ZDRMUXSmfvCdI79y1ZcEM20vjRqEIXQMUWZX//VijyLUUm+RTu7v
M0xnsupzzOdKb0twuVeS+segvw5eIHWUEh0LsNwxdtwzQEf7ZDuQlFGXpnJrDTHayl/YZLeIXHww
EgcKlVbBxKofsJy2qpS9+kQ0GrFuEksZYqJwPJcJ7I0I19axICKpogfb806CCgBgZyBpbNQVfNdx
mNKqx7xbVk5m98VMqKCJ8vvB958CJ5ixy/s3dzOSSl45QBf65D5KBelPCKcvvjxAEBUCy24H+Hyh
CJcWdJKKuBI7Etxo151PNzsyyWZz8ELM7qN8BudSktFNl03YVYmSG6SGPCAtMFIOwBwCN36/rFL5
6jJm7rk6qCFVoAi3Y2N+9oc1CFhGgcn7NzjRHSk74b6IhN3KP02QPWnDWjmWsXUzOBmP217FeWMN
it0rdrVo+5UehkleTxuEGRz1JihJpFx4IhlnADs13xmdIGns7HcHIWBQCThuTXEXgJ3KeJDlfhbL
NV0u2BkaYwCKRAuDLvE3A+yf5+s0gPiy2DEa8PpjhgCYIfBOuG+rJo/CEwaPH70GDdVHJ01bgie6
7WYF8UETEV7xtKRRvnhffSrkjkrOGM4luo4WNXy/dBCU4MAJ9/fyeiqNn9C+bzKdoQUif2ynOLHQ
zEnXhNwHBNujmDCK6CXVRaYww+XvyQKEc5fbp9zcBdLuGSyBibju2pruYKqbDX7lCrFeTxUZsGEA
WK3bvNOGl0sc5RY7POUXJmoxki6ytj477mj5TM9pGCbYDnhUaC2cVAYoDSUK9IXOtCD/EM0xbpxd
FrErQ2SUHh7UHtIKy99J769tH5GakouZZt/VRt3jKQvFs02StHMaXiDwQPAw5zAoLGhUBdycAdeH
2zK5Blt3mrqnMQ3BdzcvMyk1vxnTYE/muW7ot0otaI5V2EzfLHU9vpQbNh3w1a5NFOWd8a6Zu9/7
MsjIxA+VnnJ49Hum9cO5wRMaYG1wpijjOOAcFBGhcPkIt9ekvz658vGWOaBzNNVorKpJZjBYCrI2
YHsdhkX3piCt+fzGl3EsyGmMf9RrK50AWF5idLWk2aTNwS/MpJxyOJKMXXEAV5Gv/Z8ZJS0wqUxu
5RkOwMF6XRJdvLcxO7XCbfgrzeASgpmXFU9uVJrWN4j2msGmOi5idXMIZE+r4koXepqK4Mh7as1R
Iw30nHCZWq5IX17+VSQ5L89RgCLNaNIeg5StqgvWU2N44ZEE0QZ9MlD50XXy6yHd7Eg5JNRm0YVI
7ZuEh2axfvGVsHlZH8lr6/wGtevfqJChh06BtzI7VmQ9aukLbAxBoBeFXel+5miAtqm5sBO3GTcP
1FUfKGoHQdOUUyio8PJ+TLm5NunCt/Ps0Wx9Lw2ud4CWN2Yn0J5CK1xJlTq4ppdiS1OsVxkZ/IUa
v20eVeVGYEZpv4nkQdMPnY98jNBt2IdPLO1xoNuwPfsWOWt9161vwYpMlsiJVQyGg73cxMdN4LPN
CfjCJy42d1ILaosiV2PvziN1gdLIOAH4bApimBoCNbOk9SA78ibkESuXiCWyLrXCfV4OiVsWvtdH
d2V8Bzu0UpVxH4f2hKQ/n8l/Q72QbYVZpl5fnVkOQ1+1BUSzRxppVTwYZJE2oJQy6Y3gmmul/tBF
iCNeOgjlk6sGAIFSkt9/ZXKmByGj5rqYEAU4fkBu8UE2mtrzirEgd6/GyLO6tQcf4MeVlj3ixx2i
ASLgKciNbpgN+DNb0v3JeIairz227FtskaaAfBpksn5soe3+xiitkOaimagJlZvwU9xQ4INQ9/Ke
Fg1TIFRxadJf+7mvzrIhehoTCgl77mxUVxQg6bjceLLgPqvhnTbmE67Jnvqv4LQ/znaK+u/Mfi+F
+KBYco6I5gQuYSD768oDlPkiL6aQ6iIidZ+IZLctYAAjOIq31JqrG7MI4ncOCBFVcDHqUKv80Rfc
XUJbgHkJT4BYQWvuX8veZI/fI8U4UMQv4HUpH8MJo1V+qLYQDAqmspj7t3LKEk3xb24l8TwrfRZA
QeK2jBONAAyn6sllQsAlAZOdDkmm8kabNFqi0dr7dviZrmwqcJElnKP3lity2YpT28ttclSqdfTK
y0IiBS2DRfrelak7R8L0ZQRm7wV4StKefPHuRMpyDK/h0+UMMQo37iiFtwkwhT1Nm76R7Cf6pqbs
c86XbQtL8KRYTW9HcPIioMwUUPmDD7NCa8r3wJi+879oqmY9IX6p/uLDMiwGWrK8sQNnI5EjfqLL
CPjK+SGb89BjuoO/wfiBKa3x2DvvJRwH91ZhgiOBVcoYWJJla04ecRDbIYSGV2DHCTSHt6GGVrPm
/dByfuBM6mWUmlX2x5NKVfRG2VMIJklbf/FAFx39uKKLG5mOAwJ1Mbx0hFsVCQ9KgGU2i3z7gq9S
sLBsgDFRnK/41Ku21lBWNj0e/pulc8fiFjxCKkcVSpz4GTQc62+LVTXNXXz/mz7oO7fi6PsmurrG
4gDvEAicxf2ZGdnM22dH/8r8VJ2vJswqjq7iur97xZdIfWw1yZRPLjBKLb5+qidddHuSPRo7XWmU
Xnc1tMAFqmHyeOfv53vPbPm2el9MZUMmolXvJuS215O9uap0rYBGz5NAwQqKLWAayVZaVs30yyZi
KxWfAlEQFS8pl7cMQ0HaLOESr7T3uAkwCoUW6pl4wSzIeoMaxqrip4EzRHvJ7lcxY6+ynubyf0NV
rPwq7h+E8acg9X9Me6ca2JI+rUGsor7UDeUSSx3fPPgTbqlip3OB8cQw3fE/QqlDWDezjeRWRVUo
9mrTmssvZQjPCBhKDjgkKZuWd2hvjwSCqQ/HFO/qiWLwujDMXJWAAoDjoMjrDIS3ZmfUVHJK2hP2
wPuPfkC6bP3ov7XorQfgd1vYVGduDyXg9rYjPdgqBFSkzfOu+hNNu7tB1Io72TOQ3TVAluSQ4DcT
472WJRheFuzBx+iP1WleGRubbr3604AuWEupiz0Ekyz1oLCTR3KkDEWPwlN19pnJFk1nIegpwE5f
XI8VF6OhVE+FsJnd85pvAyHHysVr9pKAnMZ6F+AxzvmGVPGoXLFCTYAzBkUcxIslT53Koo1vBm6v
lpNmIuELhch8Z97dZwhPb5sxRkqBsz/tDkkus8O7+D+hZRGy8phUfbAA3V+LKnnBGpmjvPrBMbDM
vYbUWjZ8oLDrRgnsl8dnbvR1R8VKTP4QuQi9aGh3otPY7jGMtT7SLxvGxGFQ63uztmMHE/EqJeyo
Ko5QpDxmn7IijYO4sgf3EdHMXEFL5ur07vJGTxuURzr5aQ14kKZHmjL5oaZnjJs+o1JrM4idUJSF
VShH5Qn2dF3JvUqxAnc0/SOt9BgrEnnjnvWh3ZiHyroB/XDxrAKUcLFjrTtG9wfB4roE0pJySSIr
Nlz19hRVkpmd3d8V9/GOqmULJ5zdRtT/csFavyDwj0bJoIIeH11XOsj3RMOq5+IKvkqvfDzarR7A
CMxNfZH3zpmZftk48lSMqN6qHbFUmpeWR5EW7ULR2r0I/EQ8kf14KRwqYLGBP4R3sH74nYRJ2yyF
60XoNjuhKYj+4+09LfCmxcAS5J2ucR6j5NFRzqmIAD3eJd9/4xkjczI75R9M7n+nsz8IDAmBs0c5
JRa5WgUnk1LlTfzPwwfU1/gUy6AT6SCEG6dd3CdS5fNQvw24N3iePANy6sXYoa2g4BnDTbwhv15a
ECscVPlES5QRLa56WVyhc0rggE2zgm1vzU77INRHqISpjZsCaF0WmnM7V0ZCuGsWUv7h8LX7zkke
LQysQSf4bo2tsc5//67ZWQ3PCYfwlP2mIDEi4g7ONEqIXPU/+FcCmmIgwVTEAXyqt6ftAFqM7HFZ
la9BiQT91PImMMaWN4GoSb+g00AP43J4WwqVznyZb3E0MHQP4awykVsxRzdfpIbbvd9l0ssFQC2A
0OCYIl+MYW4h+mkTdR+Oq1Rkwj56KXKFCR+4SkHMR6ik0KZyfTvNwjfkh4JEm87oHBkaxvzrBLFR
CD4JUnLxMsTqUZg9awlpO5EJ7jmMoxLVD1iNVGSnL6SMpGM8F6EnjRnPD4ZB1T1FDfd/HG75Tz5Y
LPdh338ozZD++G21DZoGrf7wKS53U91JVm52fKt+bpYWVQ0O+grDEerMU3fu8X9hZ/57hf6YwXLo
ZOPHauTky9v5Bocmo0HzQDoZvqAj4chhIuivqh1c5eAgvVTDaCnwaVw3y5YA9Z8pBKtHH6v47OHR
SmWb0xEVofUmTHJct6+vzRo1sFpdxoyQ5aKSaem6CuXc2VtBHeohVyBI9YCmq+h8kxy0IAjhl0Ne
sToHfO4+fJkuyHbUp5UZslgKn9YfWVoJL5QH2XircqiOYWQFVvppzv2b+2L6ifhN+Zpoqea4B+Bm
af0cVOmip7XowU2um3KfblHWegxFU+txFBeX9j6TebAajdxSqPsbOIM+l2DR7LuUhy7ZSRr+AAzb
LrYwFtbnAAxriw5hG0/41DrZdeaFk1NirUg7EoeIZUimJR3HOYexe02YAm+5lAMnALH8DGGc0Hbr
BQD4pNrTk6qnIGUwg8o9dH6kii/yQFWZL4w3eS3uagXJAYiiVdzRRf3zPet1pxA4wBtLR3JdL3rU
JLbnmlqKxb0AL4xMNsZrrZMq+ftMI+RqAhcHcqlmByDlYLhCTHZ/5MHKZ2GWIwdPCzKN4xjk9RTR
XUNqsFRq120197lwp1c1uPpcdOzGlKisCPq37fqsYJ+axUQKp0ptYWrXv+5Z2jS9uBISx7iyqUnS
O/dJdce4mGluxc0g8ZzOp4Mlbb1O9/kZIgA8y42E8PBCXVKUoJBl09C7UY5FJDbUSjnOd1cxr7Md
lc9wiuiRwIJwibKsspan4DY0FB2UojfuU4IsVhmYBMLJ2d6MMblJmIO7QO6Mf3tRb0KiKEEUOGAr
314Hp+jtlRym6VJixKkKy10cjryh2DXfWv3w20RyZiM2phtnAMRbIIl2dNpA4ce0dtdqSKyX9DYg
ai6Qh1cnKVh0vl+10J9bccA32lqbavAYL5oSYqF4w282x8HkMfdSlfV5ulVEQRWdkdZR3e7QHJ4/
0YzbTUq0Ht+HEGMk4e1ekElVUOouAl5xQ+UlHB3XrTw0juVMLOhfeS197oYcm6vtNK0eL9a9INxB
eVNTDYwQspjurQ1mwBLMx4v6pcEdbXuZYry4sUHZMTzLAe881D4UXir1ZB/bE8StuBka3wugrOiw
FzEGKuHeepIJ/c+cbtnTXkrufENUAhkjcy3X7u/h3j3FAsDl9EnJHKDeiWgqpirTqgQ/AZjXnz6/
SO8BLrAokkok3B7X2cITdp/Rd2u7dRoFywoCgmXSHSE0vvdqqXZ75IwzAF7+8zxexmrd8EmvbxYy
N+e9zp3d/LdJ/VJFSrxZ6cNp9Ip0O92ixjqg739q8VjZQsK8HaT9yiE9DxonSuvHtFeKMmsFuPkP
AscVERVD3jAvGHEd3wDO1meQxUBjUzjj/8cGSFqEemt3hzj/gpjjHJv6/kUlOsYKD2m5OWbmmRQ6
+E+FEMqZtk4lOzQ0LRCNtep988F/gMyZIpcnTqBlmdsKa/+bPFnNFY70VvZjqouNjiMoCnzBVIbe
tI/rRKnx3ZNzgF2YoANZdrRPnmmhwxu9tAIR22wX8OpKPCdRZuvzvE8qkEQJd+cQksCNm4rG6UjD
B/JmdR5MVrYokhrNXogY0Tiu1Kwm7JHidF91N8Fi+tDcCXpJaloSRAHx8dtnqVXJEOzlf9uunnmY
FYHsgCPNgpLWNeA1d2NGg5EtuWlAKM74HJ8zWD6jfbPGKD4iVpPnElJGyFMke26s65lDluhyhfFQ
faOaS+4sUxzQHHJXL6Efq6RMRMwnGw7JBgSOeWPzPwpwG3QUUloYJuYG0gx+86fT8lMH+paiCKBO
aLGP4e/stK8S2chYijc1d4TfwgW4aj4ZYFxlzY8h0EBKiB7U2YsV1gU40/fmNU7Ug5QkRGSIzIIf
s/Tn/eiOkzb/eqACNz2imkel7ib/tLnVat88u1L8e2yc0Rl1RTNNaxVXGaZNJ/Y0DylqjEzyZ6Ze
cbqM911Pxz7whicrV9FVKHKoi3Cui57TcJLKG9vNAYmgu6kKcFROX96zXlegLSo7PKIcjDPzx6Ue
dCFAoft+LS40i7HnTUHRilXpA67qlX6BMGkUvXVl21nXSoukXYu1HN6hcp6qemQlSM90dDYXpnsI
teXgBwwEvI9zGzrH65uCcl/hHGL5yIJWz8LEUMsYg1unFej4zAF6YM2CTs8zSjD7tvMDdEainstq
Oi7cRETE78xcXoy/tB1a4NQdCOHloErfbw6sKcT1SJtrosCMbGhGhFCxwGxHtAc3Y+HEnGKiUyYx
dRsMTClaeeKAbXHOAGVzi4HiONscSbvB2vow9P5ovDmUJi3YE5sPQPt37bmBbASzdectYTNYeFhh
Yqf5vdBsT4o+3NJHYVr4Nl5INGJihzDpHVBLz8kZa1v1lPt9W02JhTo+NV98j5JWAS2kKZoIrx0T
tSp0kmRgCUuINlYMiv/Qqu30YwJIqvGa+sTIaCGb1GegplCBQIbTiEKNSqcTikMXmx+J6+ZscCBT
5HGDJxsuAur/AqpOM/pQ/0rkEzn+rXLc7zWN/qUbuVMhziShtsITNV4u/tWsqsC+Y+5vGvkEiZHY
ZTfPe19tWKbgFadVJlIx8CwCUMnoUdoxAw1aRyV4HHqaACnoDFLwMWTJgWSTY7m8/WRLRzZ3QUU0
op2okTKyuktnMuOzri4mcSnnjC2QRve4U7Noa6ttEAkDx//IivHg4tStTEegzw3cXl0FKgXCAG2O
iFj2pONMBSLsV+vJeLfAwZuQz/k5LccEFs0YdOyV10+qC57SSTAyyuC0Ulx+u/5sHaZsodV1ltA7
1BeAiIyFVjKydbeR3ZEyXEZ91Upr+xvstSluwwNKeFIOqwYo8b/Na8J6sgkJFVAvGDgl6RSKHfMy
apR6x/rKiRIY3Z9I2xpRXJjSzw9embi6M+4b27u65WJRo19cceb7TE6lfxwHfBKbOFqr0++cssmv
TFxwhDDe5zeJg2YICRGr4KKhZPguh5iMd8TJ9hUS5mtrSKke5DnJardT3BNJx1tn53CdZRhN81k1
UWiU0jWDSXhGSbmGr6PL3Mn5H/I0bi+9rjp734l0s9aoHazshwahcLO0eP7RI4puv8CLesDUJWTY
PrAb7Vbs1E0ZWEb0NHsfo2Bfjw5WzxkuFRxtJa6+O6oZHHvTp2atSLvHu7to4nF0JS4tlkDXG/79
+vpJSbTNSiHkTemlVbnxvjxjmYbzaLS2X6UIW6pn+yo7CrU1qyH94BZyIxIgQHk404OmvDZ0QrSJ
jMjvcY+17W80CzrVT3IxCtcGAivtyLa46JVgJJ42Mcfgqb5NEAIeJhvIKeSyLQvjRfP64XX/m2V6
gdxToRwVrX4KnbzE9aCCzusVmXWfXmaOlArqvXxH5N5sGyzXDE3PkB5oIIaPDSdbVTbY7ZD42jHt
rosJ180AmsuiRov2uHATnfV90+MWnxSXmLkaHBrohFcl/RkLIlEfqsN9N0ohvCNx9gwSVpXpVJLS
V50+tghYhY+cCJ8fXXon6pGADa8sILo9uPzCjTs28Hjsmrr/4hKKaec/zUWYm0HiYasO7Bla8qch
OH9SDXMeOsXT6fw3OP2Qc0jYio9nAenXv3LCRC/BCW1cmb3uKnz0cLBMlM/93cTbBrR6NEdJJAjJ
bcnMjbrseljcOQeAaV175vIT9+kbdeN7gPncHczKxuuLWieI59oves0Sfoifrl4ztSnEeZheax+4
cEuGVPXktg8F6OOOwBcCFphpWauId+v/OiRLknO9cB+NThNU6jbBqLCBCnwCBlAe5R9WsiM7NX8c
8W0NvHY1TKGy/QejBuK97CTME+BrOi2Ul5HhRG3nVEs8+6whUp/itiejWIsAFDS+9lksKt2KkQMZ
bofSRum5YsfEQbuEs6CNWgIes5Nj8APzvOzjBfPqwbrCmnLYN9MPQKNDPK5HFP6VGwN5oENdWYd7
88Fe2TghCW+seCsAl4gLPrQfzfFXNVfgo3Of/YVGLwncM6pqo8iJ52SOPpCMUfXbsq5EJ691S5Eb
CjOdWtH2y5uYYYKy2pFZcPHwtXEBQbzI0j6CjIOaArezwxmpWK4huXJReX1+BzCDHBr+sxkOxTlz
TeLEv4XzHAhI/kAYpbuY6Bf9GyrJrZMIqHE2hxl+fb4SbZFPrg65IW2LATor6rS6wNW9kYgwZGAN
24TEHhEd2vFI+c3TeLHY41KIcghZypA2GHHawz+eG4mKzJvWXMOKtC/wME89WC5LOKPguiHCbr5K
3aNVpyiTZf0QnmscctVgOqJHDq5OeDQg1CJJKdIT/Ne029kZRbHBGwMMgyQywB/dHs9HQgXcdFQW
j+R2FBR+HOzOikihSfSxlWcUvG5+zwYaywKtuxIEQC2QLdx8bAN84QlGNNg+WZr1/PTl+2gLMyqS
slvXGvJ8abTHdxzVYPg3KufmTfyx8dknWRhGTOHQFfu+S+ohmhWsrdez3hpKbv6+5sdWn11fPEnp
JOTb35sTEciFH2drI+9w4NpXQv4wVNk4FW8EFDQJ39pNN1NdoHnhj3xi7vS8oU7+ApE7GFcwBN2l
OQ5X+XhT60h58IUiGvkWUgosgpTDuBLjoZ1+Yv89g78cBv0e8NB0eoGPmXynKw/UU4+PFH10b0fT
ub1Z9iCygUnTpRrKg71l8+J05jPscQ1+r9IZyj4WReI92aIJlf1fIpvX+gu/3wVSvV5qQXS/aoio
my/q5F3swC+QDP66x3JcaT9TLJFoHfGPi6fdTj0RXuWi4yav0tWfZmg95lz/87g8PCmwO3R5bYW3
76qRnXBMBACkbeotfe+wR/QPVut8vyGelUdq38gU+mkyXn6vWD6A9DB7Xr3IwnbwG+dEQuf/u8Lj
lrqwMEv2Pb3CpVZkgpTGpYznE5CLwYKDCvzVJS1ApRBfWuTzUs4iL9ZvOiLUGh9TVtHsFu3oOFiU
icQnlZ77yYMJy6GYBPxibZJpyVKnuQILsccO1M5WkgLPQCRi1eNQxpTD1XrsHTnsY1R9arGmWQoN
2ogDPKB5z+Y1ufucyfNjHNV2JAZcs8VLGYhBww6pP8b/Cungo5+DCIMpOHXiH0kD9E3ShiWLTv5c
A3vE4WywXPMmdSqfs1jdhWRW6u+/wSrQ8aa9FAkjjF/WrAnrv6jVZqxu7gQN2EOHpsCgvGYx0+Qu
OhiO7khODeZOKcpaCFmwnytB101U6BVPFctEsrz9DUIfAfA1KzW6I+0dPj/fx9TxobiwGSIa2AhN
Y/eBlXPM37cLZTzIRty3sSI3lReY79AdOTg+S6rVhtg5/K/izZKPoIetpkybCe/hlBK2NrzAtgLl
RJcIH+Jx4UhYiYNuuf0tw214APeTac3QeaE/wXZTv5FEqL/namiPRX7s+KpC9RYJARLOTjpiRMaK
BeBTbXwF9naeAyO1rBPfSRO3intOhKua3nktCNCmg+v02ATnxjfxgZfyzmdKAWOar1b3JzOtoBnq
puhu0D2+4kTjQIeFQiwZ6k5687iJ7CQ7Go2EV9qN78VYdp3mfMdWDDaj+lx/HrEOTWxL0rov0Jp7
gF/sW/6T23rRhfxaGvBAJTkBrcw8jQkT2OLI/VewoerScpdo8MOjHh08u2lSgOEUvS3M/8Hl+1gn
R4y+aGmyRryBqPDFHfdaFz1ChOFBS55AIpnSqQnkTHBr4oXJiuQbEUo9nUfFMNS5SMxWYCZv2yWh
wEtTxdEL7eZe0VnJA6scs3o2MF7DLzGdSWISwfnohI3JMlCOZyndxUabTFpfbixN8TQNox3tQAPn
oEglwU2ayT9TaLXNjjAteotZNYroD8e4lE/9cbf3TGDfhuOWnSUzN9ok+MXHlRSONvSWu2g2efiv
YbWvna27UqwscUw8f3WYStEuQJnHasDATrDtvOOyUfaAa7Mfj7mZaKmeXFn30ZyxvBGUswCmEmwA
kFuGTrhAbRrfZMs+e1bygJI9yvjhgaGgjLlmFSuZjx+f5BUMxeDyztZAP6Z0mGn41ELT1UjKCZ2l
Ej+SFADAod7qQWOZxn/fxYcp8CMVaHZdcFcoAFIMMWA4dENIq6RbhRnU0Xb7PWh2kPMlY4eaTFfp
vUSSqqf2hdtSouLaO/1B1ryvHRCzrEXjQl2lmUe90ctkz2rehXTmOWGVIlr+1/6WNR4nlf8gL+sa
CjzFrYTd9FfWse8JsJr/zka0YMq4X0j7zf7bTPt3dLqK3z+Xw2xp6amnNVBQBeWVkxqpflsM6hBh
StTL9jftjTNE/KrlXPgChqZd4OJzEdKTj51hADIkYpu2VDGV4FO3DYZ1BgUJBZypa0+HWLaOc+q8
+gg4yS1hMlntCR/1jdUnr63WxYm3Ilm3eyopZ9NS86JEBQYoA+10DtOm5Jsya+DGdi8goDl6hPAr
u8ENU9YydCeHK5B3nTGS1SJAUSHOBEKryOnGRpf6DG94jxkADCAXu74uDKOxe0s5lbupuuovPACW
irnp1Wg1TktiPQtv42Qck3DrxIrlbuhfqydzQ6WYcHO/FZCkE3GjjCWzoQ4pyfm+AK59tjH3bwzl
GDsGFhXt0SNkgdJxSa4iXVKB+I1YE1wdNukpe6PEohhRjK0jd8BvlJcogr9CJzYYmweySUBn5Nkk
nCvsITHtTJ9uYG9Mui1hiXPC+kojmR5DXXBFxBpxfasQv/hZEAUGTUtFACFDFZJlHvLZvEZVcP7r
zzvbg/saVvAE2KfR9iXWEFrNXjqOiSBZlhG85q/ml16MPd/sNRwSFhIKVanNhtdeIkVVf6gOH4cU
sV9cDS2WUMIDTrEm0aZidAaayZ5zTQyox7sV7/4KgPzPs/1Xq7Qh55QnmnFuGTPiTdpvBkNig4fA
uD4jysdigzYmUSD3wZpobx1c9EqQwQl0Rq9PpTydSoOHwn03MhPObpoV8OIlFKfnuBDFmfEYFYC8
wsJf2BTTPc5V7bXMpiE4WKug0l1YwzgZDsRfiQG1WWSq05jDkI1zXWOr8Bu8dgbKLKOSstI0IUtO
f6Qi6tMTSp2pdtfFnEJ1uNRGyEQgCu6o/AFTJvjz5rAPu1KMB7V9T+4qWLT0Lml8HCMWRhesNzyL
t45jDNyWAMjYuC3Z0wIpsjFzClvWkxMBFu2wVdHdaexRrhMa8PbLMOooRRdC1RWeMttd3M4fHDfp
l4rGsNCNslfkp2OEOo8sjVmaBqSHtzyDf1gEa6Nwdh9+lUDDSfBRQm9o1HMjCeNd2GmmZ8qzOh8H
EgfQ5BWMInM92s333UGitjg/dnj6UyYb35akoEYKUtwiauz1BpNOyBfBZPsP9fe4g6NiLdhO0tzw
UF2mAIUEyX8UZbCpNZM92qACOfBvXF+KDSHXA0zPR39r9U7A4alcNc9kR5iX5/1buNQ10fV1jgnK
w7pbXFDTRzNGw9iCM1Wima9ZiR65xpKXlUXfe6KvrrhE7U6iVgYaO89qCVmYwhX7dmF010XmCGyX
LICIU5H274NQgtCHApmzcjhWed6Mht9RuKC4SI3CGCGJkX556JGQ4c50rykNcFWd7fDZG1WRAD+f
GQhPaCNEAY0FJqhrrHGkbwmwA4xOcKL9E0KT4r1IudeoRrPgdpR0lV+8JA729+vSnf9I/NOZspw8
SQQxRg2KjhI93K9I5PMsP9fxuZ45ahae/RoouF4cMiWuG7M9pvOMbdXKMzqFDEjINDUpC8jFhAfg
KPPqbEQVuQkzd0MnyW6qEmql4Dqjluz1py5h109Mx9H9+/Nljlmn/Uv3jKTBt4K3ZRRLFCw3oMna
E/L2s5k7OvS3Mft/8r7YBjci4DgSSoQnFGbIKLzcp8x3YISSqWyFBtJgdEj04rMPJc51+R4w453j
SzeO9J9eZdpDiE9DCcaeebdRf9CEtGUsXPzQGC4abP8t6gbQ6JOfcJYMXcQbUZHo3if9DFHh3eC9
MQSXvdChaEkXZ6Fu9UfX0OexKMeAWXuyyigDlB8eghQx0Bqazia4HCc+a7FEpG9jkp37jDhrunYo
hCoWB8JUPmolt4MisR/erzmK1/XD834nGBKA0Az9xUvtI8Wz05+oMxXmBkXtaxxF43H78EfHpr6f
2A1+KKCeR+Qv8QGqbMm8MxkgXsd63D0jpJeLYo2SVVL8Kgt1u/KAS8dFL7tiXAs40VwUOOXDq9L/
WW8T6uz7nG5vJISMA6pCLvIM72RplXNQIEyM6xMKOwB9+v503tPPqCRGKGgzj5ESJKvnnqX6J5aN
SE4qZjEcC0mDV1nKboe0M4ah0O933pReTJ00cxL7T8jHdPKwWkqa6yRncC1bFXtHddgQCIWWW1qj
+BlZcN+uJLUCyJlNe09Pv818eOxC8FK14t0wdZy3FN9PQPrYnNBxsQxjh0pNUvrpdPxfHa0jeHZ1
n5zzbFqmLXudjpKLe1KqnAzRORtV3JC3fTNieGUjH19svBXWqdUmEzwhSvLvUrbZXlGrjhDpGjg+
sD0gUuJF7IDjxmdNVFEI7VasVyTR4NXmzAZDgFPKmTF/3aMetiz9ct5R1tyWlAoG8xsO+em1Wscj
Sa6gh6arbVMe8S9CnQfchWcH9a8BjRwR67IiJwYWBS2nXfBa5ype0gVJM5tlaCIEji2IrVAwiJNF
6+emWrI8ndmqtFSXs+7jjb0j1lTmojl78P4mU3MBnWJxlSu4W7MgSrD099JeHSZxPrG24djibl0h
M81YuLE1sXwDP+ewHCTuca9AsJV5N2psR1D1gkY4qt1HubvNpxH09bKW3Wl3CElMscEdiOT/FtZP
rWl/9W3dLxCE/bUdmjHWNkqAnkxRMIELjpIWlXFM+KBkQafjCaq3AnFIU8eVfgkTy1xsqP85KAV1
JnKsRmxN32OkupmlEE6bH2ZTm6y8DqKG/2fgsUhbrafgW8cU7Oo12WyJ7AS1qOPqdAjTUlZoQU6m
SkYv8vuCYgHQs1n1t3A+z10zc6Oa/J7tWHJ8NgDeOCkluz5mKLantJSJR3WfMbmvHs6SYO+kQk9I
IBMkGEH72+Km0EiZW+k+jwkws01K+yqDSsXQSKQSjWpBvCTuNVCe0rieUX3cYMq4mDDsLvJV+iGM
VjwAFyerm2uV5NccEDwdvAUor45Gu7Vexj7CWNzYWwKAqTSOxoWU23VfGbNaHmJxktdBGQDfG7Zj
pPD/PYZpeQC1GP+riosoPNYYRl4K+CWZYTtTH5IS72tG2ua9xWR5mwaxRsanYvoXrd5RZERiA1j7
6VZQ8Z/zRGa2n3BewlEqTksnbGm8jf1sCZXOJGkuJOS4rMrzh4VsUS2UrVWajHJY4WFMrs+O0X2E
VX07SKgKzGk/Kvf6+xthhQqaYm9f4Gg+vycV9R1rr5lbIMduIJ1GD2X1VWc6T0xaEtd0BOHUqFg4
/sMM2tbtOxk7lf8lQu2cxpG0NzKE95wZo2wRjKwRcIDivVCmP89TaS6eZenI7vtO+vpQWfsInn3B
L6iE61/Xa26o4f5ZR3MjrelRdfHfqheDxzNnVd9iabSmhARk9Nm8svTj05jJAZwNJiAuz7bC/xhd
gs2iT9FCeeZ8LLxGK95HjAmQDS4FMIDcY/lt2+RNQZ7u68LbB4dymXR/vW3wbMMXs6z08yFw74PH
L1b8h6TM94Fllk81tbX7JtjtuXXfrYR7Ilzw5lJ7VVhkTIsf02UxR8Zr2IAtnct+OVFteFRlVFdP
iQAybCD+oRggIPlmHIncZqpEDqqRAs6jPcpZF4gMtT+ePgXSsTpoRhDeNczZhakRfeIQ9CD82H7A
jmhrwEoBuO8jBygmO9Gz66hvJFSEDroJO4Rd6PkLRrrz1YhM7IWTf6+xbOnJcdcopwNievo6EyA5
M5e6quRvp9kXE7LTw4EPQ4UC+2K0SRc6P2GYcWk+PpRELUXBuZaTx9BQkyh0i1A4W9Kj6S+DjyOO
ZFA3wY1o7kpJVloc2H4LSfwr+Plv55xf5BSLFJnDHgYOG3nFBM0rLgaU44M/IsO3YiUVy8LUB5Qb
mJ7LeCa/pSfXGFYVTeqjNN7hh/VwvcztmPR4mignM4FPsiarFK0uka1kAZbsIi+CDBDD6xN7d19k
RV0blrM0O3lusHbfOeVHWd7Q1sWSYra8hFYGvLppW1dZA0ZzIL1ZxRgCGAsecaAcfWsKoocsV7mA
4Us+OdBQcWGKcLe7ZSNMwDOAPrww6NAU8qbLHc+eoO1cABwHpsMva9sQK+gDoiyy7Ds939YYCY8U
O1Pv59H3XwhR7ulHYB2FIoQ6nRkPT5Ic5NQ3pxkGsAbgyoBtnGu0z5b0qSN6pCMV30j6TzG/X9kQ
OcMY2tuRhrCKV469TRYgojf5H+g22XZiPzqfmD8qJf+rLXjcSRT3dHLRU7LqYdL07JS1kTyvuEbe
8rgq3uYQdqSTJs0tQh4eUaM3pl4Too9Dw6PaTO2MI31zHVv+mOBoxMp5gZruFqSKPB5UBJCV5Jj6
YeOJBKpNxthqOdkPQThxVuZ3Aw8+oeDla+dxxO5I7haSXoPGrG8oo29JSW9mopofUBSWa+IaLag1
7r+Qa3csbDYgZoyURrsGzmjUGBBTMbga6RdVepH93gF3P+VAQ+T0b1a5/z+k/nqTrzx8haGMPluM
jKD2v/DsAKoKRNIY3C0n66/V8OIPz/hN1lUEOswV7AbB0M7FZwcHwv1XfBRgHyfMrElpr2W7bogV
t8ijM+Ek7AQaSj4cAjA9KMxR43Xvt5Tc0oHkbfdvCc7HMDALLzykCvIcCtPcnfdSWsJUk3zaboLa
8FsWKZNHibjoEk9GcJZZmOy7rA67eZZ7Gwn52cGymLiIQhlnmP1Hi4tqjkau/DuyyHBy6u34CYtN
eBoTJHReqOFcqdNZWAkUwFZXfLrexKvOQVdQnpzr3OirZ/8unkjPxImRu2bZRYwbYZk5NUsE5xMd
RUnJEW27xM4LEiCMvMRIZJd/JgUXZqttU6YVD17WWj/Zrw1C6lNTfzJcfteOpbK0fzclnsRWkUro
Ak8wOh0YbCAnncyzvuQKPsGlgF+7C1JyyQHZnl8zJdKyIwpnAR97V9uFl3vrOab0+yF3R/jpVRBh
MN+9urJLZwwnDFFVakz21VHNvgpJmy0k5AWvffrklRU6v6gk/pwa9c9a+pjTkpQp+Zb+RDJa+TeD
fENiThzDcuxj2A3ogPKRPwOSjwCnZr46AKDq88u9yIGE8KQJ4z6EJpgZf3ehn8GxzvHza36Pv9pp
UF9KjkTVh41qHQJeJo2JN9uc4e4/q582tu22qsTTc6g3H5blOywhSorVH1+O+q5HRsqTIS7Sn3dY
f+rKQUJGHc79SXoRXw2hpBwUU1RO+zfdaB/4cCDgTuBJ3LRwQJfUJDb81JqAkpH68cvXYaDyFAOG
5MENqZyEoBY4wU3bhX91YimIYKQvyCpNoatpBf5VsKnckhz1VBjkPTPbnxjMmPuUDmZ75QkzhZxu
eHMbJGbP1bmKmg77qcVhoFG3NbHn8UswPZF+ZEPePCXGPyX1e24rxBqP5tNOKdey69TBu+/75fcy
QZNoov0rCLGXDvRGwJGjCQdDfkUlHK3ITG/8yaFlWEOCq2Ynsw1rpEl+XtrBKsFSoAj5UWrXjqac
B7zOlgUjHFcliUxNXePC121qgJxcpyBN8NKVfSXqfj+DZexaH0Cmu3HzQdAYcdI81LYa8SgZp7Tf
kCrOgFo2g6cr2Pix5EK7XQzjV+8sexE1NAkvt7mLummsOVm1RpgehIH8MtFXPvNTOaoDzzqzbMKJ
ivEzEG/jSzkHCDDGg3mA10zRUrBF32pCmjQzO2iNm3z3SOmruouMHnq806REMXIiARod+oUFTVPG
NCX0oY3/kp5GZo3k7GpqL4YiPYBI4iYHiF8grYuHN+V5dkc4ZKifxbhxa5Ysk0PWBveOrpMFgD+K
lLyWJcovHu8ekl08ztFkcLp3rQjj2Hh5bRdvAr15c0HFyd6RY1+2iBTBnDASyUpcIbahAaZSoELP
c3eM2AWwlpdnjC6wraGhuLHe5jd8eHlr2UpUTYPwcmM1+lphEv12eW/lBp3qZmsmph5utSvxosD3
zYSyNWy0axPBxygKZGhnk8sAagUIM2SB28t32vTkFR9H9Gl3BpG2sjV96Ottze/opiZFkukw4hr7
jSXZKjSPHnxdA8cIf9rj2SkSu+FcKh25adyGCSRqwZIRA31pRs3VECQrIgNWw/Ntq3zDrCsXo410
NYabFgxj6H/EXQMgn2UzkPShuSdg6jS18S96xy7zxhq2RYvVj536DtsPMLi78+70U9UhsaVr22jN
qoDrxGd7uXFjO823nc4JpapCy9nafmh1ZVZymcIFuy6Gf6hDnFzp/KYecYaFa3BqOkPuRnvAhNNG
4FJbjPUtY4C+M2w58hBs3rbT6RfpK2qECuszcdjKbS0frRi/nOcG+BInzEfsMGyhTk+CuQ1zpsZx
oA93E2hYtdSBy0ORy9vnO8yRoYyxMGjLyMvwTQw7ewbICZ+o5G84Ua/03SjjFDSZgXM7ycyFeHws
rUK8OUg/23/yUQU1qNgXGNC/6jGdXYZpkSjf/rX8n1gWLpiB2ETI+kPizthSqduy7Hs+nPtpxEFh
azIPNBBmYTuu9iWO4p3FuT8ipf91WXiQG58r33QeZFNsUv20Ujt3Qi4f3/8DUYkByj27kYrbTe/z
16rLvxygc9lXyy8OC4WMD5C9S6s0aSAQ6Lf8aMuH9N/K1/EUl9dSpAxPCKBf/ubfrxiLLMSc5yU3
tCGzWzbTL4BCOxfqF7iqP9l3wOWwxDQfMuuxzyW/YvGLmAFGPBpSoophfKDlUZybWGJ0vb2dhvye
aewPquNZAnaWg4zyRV47/wEoYdnrfcvVqc9wfAchyeJceYEJRlwBAb/vLzYzbmOy07LpVvANSRWR
qMoIALu1YnuE2NYV3m+f73rPY+smswSQ7JB/F+r6DotgjYSm6ki6rARbU9AZuQ1mmMPajOiAu1OR
UJouB9B9Iyr3hYG5AdAD2ir9KtpgkLCikV/a1RGlqDM7boD9pXyzKe0agv08c0syD+hHmIGpljdp
Wk92Ht8hjHpFSMJWv8YFinVfRQks6Qi0JMv3GEFw8AQD07QX51Z73qornaO2bZLKQ3uXr8MZshxY
EAyUvDQk6/BFd0z4sknewnL8wrXKjdjcdPVH/oMbWUjYtP+sBAnkwgdEtKs+/g2xSy7TMqOwNC/t
HwEWR+F6zCia7Y0rzowb4eRX1UjfES3VQfAA3CIQQJDku1VwQf7Sh8prupE+ClbW+D2jJmEvyvsf
CJwTZJs7I7BJ51oWhZxg459BA1AtALltHhrj7k2gdaxOTlY74xVvp9w4IfEUaBzLvhHaG/NY1a48
KU1hdmuqSUVueiQJc035s2AzMMmlMDdrYIbmjLPL95xjkQzGWF3Vf/ltPqTrzfPWW5kWDe8Q6pHm
a2HqRyp5s48GG263nqhrrnwzdZf2LiMLMwtqxv3pbhewB1V4umTorJWqxsiZRSAcMyXFXQ1ZXNsf
mVvkMPNi26i4BDArMcl66cEv4bm9c7P4ysqvrBtv5P4yapqyQVQQci/lKWzUis4G1kM3HWxdcaCG
hSAVLaXGbyutt1Enp2Po1OnC/7m/7esnjgp0/GfPBOxU7p9Pzjgg031FKePAssBW6O7h2CtEFYb4
+eqXoNx5gCMGaPnJ5K7m0KYbFu+3DpFTq2C2WtifareOXYvCiP+sZ83MkvtNGGcJ0JWNXGpLWGon
zC1OMhl5Fi5MBRsyS3BCrmvAxO7h6WpFqoTfFdECaUIp1ZctnP/rp6GT0TqPhf8AdUhipc7rkzha
dwVEoyFiGT3IPpHUqHlv42IOugornv0BOBH6sLC4mkPCFxRzf4O8KBTjtkD2z7AM16v0/T5D8HIH
3JFzvPQE+Gk0vjkvFN7f5oPVR1xoBDbfKhqe+NMbhEj4N8FfoGE0O8T50/ItFdKbLBaxCOJ3uFW3
RDIYXyVo2kG4JOPCTbdjyYsHijZ/GpIgi3I4zAHTiep5jKaxuwD9H0aFsDD4lUGwjkjQPSsSlUnX
mZBsR0jDq/rzIEZgr3B8CdAstU9Y+LUlrT5O8/4+86oB2HT1J76rN1GI9mCr4DoLorShx1a5dEA/
YSlClOfRKix3OgcAkWlRj6j5tQPhmm0g/zcVomrQI8p3au7ogSAWfF3YxNmLcWVS2UElIJiM2imD
fY7ZusnjGkHpFasSSvjBu4b+HWAGDaegAOSD7CM4iWxxd+uBgzi5wafuHTh8s9a7ILpOVC/tJkZ3
J9uVzgWpdOuhfs6oMumg1BPpbqBKAbODW2XEHywdkOp2P+I+9jRn9RkRgBWJwkp5JZgThES2d0ZD
0QiAsq+MVE3VzgS8wmEfnQtuu6Jct6efsIOjygyyZ7ZEBJ6hvsOYKeFJGjn4POe0LXbMnqJNlHnI
Gzxk71X6ZvqkJTfwz3V/C+fD6qIX/7VAb0tXF4yYiRrXS7o+GydZVJw9s5cSCxVB3HRswseVI/GH
tuHh+CwAbeWu8kMH9zH6OEgF559HnH6FzAD07QaBeSFioGpZtWSbnAdSoqpbQT2XrgRZnVHRfvyi
AMUwxz8GU133wPYmw6vbAwz5Z77lRh2AYtfd5mf55XJj+gXNAd8hNARQmZOKaOUwUjuPXkZzssXp
XcP9KpedRIVT/QBtZdfM/5oFy7MeIh5YSDxU8bWxNdtjAdcl5rxHGK+R0S9MQsy5IsG1cdLQPNb+
u/nDHzFvPuTp3B+4QXkIkqM/bRKwZBIvULH3HMazHphRTHSNIezqep6CKWKL+ulo1eQZc+FFV/du
8ExMwBRbSNlbvKoc4ZgqKzrxIQSKPaM0Bx9GBQVKlBMm7id2WyaYR7eeYy4d5p8LdSFDIEoc1d5R
x8wK/nStu639VjZPkMMxdFGeRPc55wzLLnecE8GG4l9Pj7RxudQFb9qw7FvHqVhESLV/lW5Q+bVx
d6CeqL3cCyaI7ObM64wG1YnDlcEJ2fgZMMRlEad5Yk5Q2ST4bcZZlcdey1XP5KH+MsnDkULQT1EP
mmos5sHiJBvA7HOb8PZ50euS3Ca7sQaEbWJjzxcgPmHwo181gDHCWmbGNIBoxHq9fsskBW3c0T6C
FFBa04L9GpRci52Gg6NjYTe5P7YZtJODFVc2bQGc/8sGvFhwXl2PCqLpGtja1FguJ8vyuGRZUgqy
7G38yPFf9MSYDa3/qWgPEeYPhzjtzoo2CvpuOzQLsH4Z7dNcW/fkjcE4Bt13qINAQcVt2ojxX/0G
i1JpgXUYw8pedhCv02/8mkCASDkqKPZ7nDPOjJ2TmOB9rayKPCCbqreT2GulJgiuwVJd3EtEbtj2
KS7wXQoCJ+MeCiiCbktN5Qw2Rl/kduR9nWo4KCGaMj0yATHcrXr5qIWLcXcd/xWYEK7jhynBdSwS
wsZpVXrLUEiGFsK3nWqUW2M9EoeXkeiBeLqZVqRyAzkGpxgl/1hn9x76h0m+SwRkbTXiCPaaJvfs
hS1DusmN+pk+H1j2uhbgOgiSDPHN21s1e+SyeplWoVg86Gz/qvUsxjNfvjpo5OSrdgF4Jl3GGFaP
xxJfd11IDrcPtbjD4WSA0smeZeCdkomOPcLuEMd6wQtEnbHb/omSBdZsUJbmDcKiAcYd35daxhhx
oBq1l1UCLmMHybE0b7HiIW4M0THXPyWGbQjhbGeo285KMO2KvVOvYpVn5/MEB/me1yCMvszBvx/s
ISjgs7H6JktbTbKZb4+iRjVnBBQAn6fTiB+NipsgLby1Xz4V5NK2sBXHNvHe+74ZAjvzvAA6zW7M
l2SpjFALE8CqMHQrwOjXgRqDb5951A8uHeZlW2J3IwK4XsO6MWRm8rekbICuIQRZmlWfspf0ttQ3
sjlDLpK6eCfgufAPQvfPSY8dpTcz4ECTrQzRVwEiYP7cmEyJj75L4r9dLqSc4XtfqNcGrHwrvSR5
uAOFNnvcJ0f44Kfk5fAGd1KC/0Mz4gZLzvvC5CMw3ryfpTKK6QlDmG+nZ26I8rXGKPwYF0nDiHCk
jH9QyCcvPjz8Nb2iPM4ABV/4vArO86t6gjqyemxSoOSvo101OiJI3JGfAjNhCKjDntCGF/rydWRj
Yuti0AHvcqsxxc+petniaFiYfxnG9rot77ieOAYPhpT1jqKATmVJMy5T9hTFyxKXJfjDiP9fbzzd
N2PY2FxVjeTLurQVdsU64n872ycH5ewQGnUm+18tDZb6rSMmk1fq9z3+6HiExU4oI6Vo3Wm27c6e
gWg2b4QbB1ztiRxNUmQ3+j0Agj06QBU6n1d2sivycS83CRtTZmqcXozdejtfVY2+nFr9P+Lkph7q
2ziEfgTM1BuHzzG9ljKijhGywjE9VpDYtpHe4hnAHK6zEKTXUdUJXdQyObGknAczO9yMlc5OmZ0V
DLSeHaidg/h7uQEUKXVruhY2lfLPq8HXV6dbTnAGtarH2QMbmMQprvnaymOtrW068NjvndASvfeX
eUKoebdLKyWQfSVTgVwCdWDHjQZHWvRNpbhcb6Ei34hKUOp3+NrYUVIepqzwIGgLtBCSmHBMVIv3
MHU08/sIxwm/quNekt+IzIoz4TBnkoG+c9cn7Fwe0MIjFlXi/0z0BcFWrqDEiID8EIhFXn7yQMRo
Q0hNm2lgj54m2hOFDKH8Vyxl9UJrW4oHm6avtlz2NDjU97dZ3ASd09xMWDN+xeYOoTuVfiLz1Zev
XGyOjK0QxKFkmcStRHzLTurtqWjJqRVDpkUeFDsetm/N8P4U8VtUQvRxDthPlNzFodG56QVRoiCE
53OutWB482utn2WocK9+IQ7Nnxiqm0EY9fsXQZ+tMa0W/GlAE6pDM4m/haqphDV0MpX/sMBAmZeO
xHlzFJb40W1scg5AywSBbqPluhrRsLy7tJrdY0D/9KbKdQ9gyoMJclnGYGrXMavKs1hOX7bRAiha
kgkwq7iF+3D4jBVRPcZzmUskBdcx9PfnQAnWcldAfzinC+tAN1TXPYWYo9wRYLumvW8scIZHKjki
VMhyM3fd5pX1IaRUtdbGGhkOX0zmIUy8Q8yOFc7YllnV5NMC2mRdD7WMuK9ay+5/FDUkO4oVUi0g
qms9dqCDDReXE2YOKZpKusuEE1oeh+Q7+lVvHhZi247NiCyVdodIUqAihqnJ9wyM1nyu+8trnUuA
Z8q/OQNsRRkmrrW68AxIfwmUl7NkTo3C2RVedzSYztfEzSTOCdd7v5BrDbZ0kpqbcNHmlVlYvFFZ
4s4XNIu72lEPpG98/2FTNHxeZRScaD2jjbp01p52G3gTAbw0lnwoEKswXlre7rtfqXG+am/1ESqm
5ePE8L1lghlqkwPIZvzjXddwac26OzEyUgR2FDoEGbv0XBIAzUm1VZB5nSMCAmPBQzUAeqeYn8CG
yAXubkfha0z88sR2+Ay3YeQgz2NYzSa9uymbwhO4RGxfyVMpZeuZglZOPGlbOJfdxYNqWEajSt8Y
vl6SRcfnVklGS6b0WZ5e7GodLbD8f2kxXxoszOTE9cw1MwpKv8kQ9LRTQNYCDhUAfwaZ+gwYwFqP
+gScYdC94C3aHpbQnm/qYWXO/qgSga0ff5AEZRjD9iRflGjdofOt/iEL0SH83jQ1Ue1CKPJFRvyY
ACwMgbnxHsGG8P2sXH7DOWFkXXt5/J4C+bHZ/CAFVNoX4+g0xKDNNUFZewCgMRp7Gx7TLvdbk8Xg
rcNVpGagA82nqbm5zgoeTmrDIrQIkXiNkHWdECpdgQHLVHi82oJOlpaVz+r8P3XuKAk9pWUgRTTA
F5hW2DtyNkjmrQdFin9sF5iG0Blq12CO11F8xnjLd+Ha5fWMOFwvWssgiW9HIv5LxDxX6oE98FOJ
LU5rXHWNzoHwcsbg7Q+ihtvDb1TR5Tm3SEVpJoWoaa2lF0Eu6BcWTEjgOWYWKWPhTITvTTMrgZJY
wA58l577ev0B6y92KmiPgUncgNR60Cha6OUv1oU+MHOffaVAX8A+LXIojdDiqSD45c4nW+rXolRS
fOIaZKrwx+HVv5nPBfQ20gQXJpKsI1Omglb3HQmh7N2bUe+RNVZA0/zznzrVIxWyJxx3tDfEsqot
/MCeKIMSndAdP3le51waZ5KngL7fqNFMAXfA0pgGSX50LYVC+Z1iznPiFvPegU1qAhkzgBONXGZO
6IUlKCpUFzaueHMhTQjWHYF4snYxa6uqcxpNeWaxSXeD4h9uQrZWTB4r3N5bU9rk8+OKweXlzSu0
b2dwhQh2oTZ8XfKXMChGk9Q7MyYJirOCmFOpks8ud+9Bl8MgpdQ5rY4O/x5YB0P4aOCeiAfUgfSb
zEijOFFZpe7jExUA7XeL4eWvwT3vt8kZN8orORTtlIzN0eORCGy1JtOkjOY7Rb9CGifWiT50uC90
YRST4BdsU393K+qF61knHS0yCd6lgxRC2yD3d3SAYUe0eXqS9xLQUnb5U/9tg2xfNxTPJqAV/neb
5B7nw0oOpMKhhjhmyn0uaM7hncdhY1oiMG8vex7ia/a4mw3RsuZujuYrRUeMu2/s2/9Qud2zMoRh
2PkaF4CKKoZ4rBHUAP5O1ClXyikHLddziYOWu9lDpPha1+faluKFpwrrhZU6RTnQgyKNXGxfYz0A
gB1S+xCZ41XUr4vG+2W4ij0T0mq9zB+oiM1YL4QdEQY4J2mDKgkAGnKaT1+pzAyeeaOXe8R77kNZ
5B/6WtkxslCOo5P8nVo4j3FMfVRCFdk8dilQpbsD7nXVNWpEUymfSyHE+2/J5/RpUzbNmv1n+xV5
1qjmEH7H0zdsAiNsWqOcQGpK/l/9YxchuIRxlxHyCCqyXhd1NLVP8QLcFVlxvyCxPvZhR/YMrk2/
Oy3fWSfyTiFsLkYjVaBE7zgCiIOOHYbLuLQxJADblS+d8VT/9tMlTHCllPcnYMlr8NGHHhglN5dR
XYxb9I2jWvz6a+D3pvUCVYzxY1rZsbT69ndn3Y5yCnHk7sw3bZVoJKpyNlgXQGhFpnPXC1i2k63w
nzb49bobirI69TBHbwpaI7c03fSeJxvhuZ4C79FGevQ5lAcAQ+iIYWGZ73N0elxaWJmkr7xb1Ryw
JA4BupsurPI3nVkhjskTKO7TC+Ks/k/y1PAYBe7NtvXGzONsxtpkWX6cckEaDNxei6kFYbPcz8D/
WCw2h6abGvWXwTg0jEG/puqJjAwonjcDu9lmZSv1pMri2XKO+4Q/1XEMO0w66freTNT76Bry0nqD
uLgTyYEZ0IjqLTK7H7b2NznPprIUWzc78czeW9PgRSJ43xm41E7/1VQw8wR4bVVK5ZVA8sYTrHVk
RcjTHxr//LsxmxqORw5S75NEzBUebxJq3EtJHUwpO3DoSDMKas/Vps6jx7GsQpuH1QQXXXzLbwYV
EDhTuNRDHJd7nabNJHhBvHSelBp04htvl74S1W5NCma+8iaC6S6pf979gMyy7iQIP3Z3qemTYSSJ
RiMrcTYp0T5NO/8KR+w9NN/kktefN0lBpAs7vbSfNz2DWFaOmTSz0tgvVvb8eJxSAaV1ZLMcSyks
+q7gXZAe5hHweQLveFcS6UvZ9QhhMZKew4HlGYqR77lC3ScX1yPT23IJq5qhroAKdjgXyzXc+mli
RIpN4EoKihMdbjBP36BX/TH81KY9i5JZ8KFuNGSTZH9rNf8v1bSde1tISFxiQhpLNok89T7+rT1C
ikClt4ETMCNsyOuMuMNfQfjGcrFNZAjJM28Xn5oZT1rA1q0FFkKtJPC1PWncFcfpKItS3e5bKRnz
U5urKbb21k+OkiVYjcLD2/s/+Gpa9G31+OOugmCoRTMC2pM62Z4cyli22KAjZeNnkZ1lCEBTCS8J
7W5nKO8BCOxu/AvHHDFPysKSLSTx6h/16PL4qxGL62XOzIFdAJzokLGWq/rvDD5yp5WkOKV1yEsP
2pUfmLBXdHo0++4EE2UR6IrJ3MOr4CY7cZVxE4ftlmjhsR7HPZcte1zAUn7m/81hUt11rVUzstv2
+MiEpG36f6gyGTHfqZdtYDLI0dP6XqdtOwtCHuUnjjaiL9ca+V2ShGt1MHPIVWc6zQ66IcnzvwQG
PHW7pcZb9L/KoMo+8Wqa/8OCch6lEMGTWzhunVivOb7v3EN4j0lHCJlXVHeGT2IJJlc/apDcQPes
7aUazuQ6BI+sHeGlrtNmjFLSCwe1FyYh8Hxz5py+YHw4fPvo09n+i9u107UIGHC9wQgGb79kZJzy
hdCjMk3OrFoeBobfjtdBuqaK3pPY/MVF9i6IaEWFSf4KqneOMgfvp+ia6h8Y3RMbCzaHh1uCPtbn
06Cxa0fCTcIQKAo7zqk0u1jBYuvojmDi7PvfSW3uIAufRbM+XYMw7sHiTr5H8o7ua4D3FXBHB0Ji
jtcYzZD4ZVg+Rq8hBObY1qlEjmj7c5/Jl1/fuHJ9ZuNCpEt7AFsw2jR3Ot7aTZDWFGDLXbD3JGcm
PrPRrg+TJZrWkAFsFlL5kNoyXXXrnChUw9TETQfa6fKD5obVIrwj4rVaj1JnWI2bhY2BA6v7gRXh
k5J819hIwr5riedDLH+IaH5uLoDzZC0mxgWdwwSoMlBbJt7EcpUNJDB9PCHW3xb3awV8kNIl2Ri5
u4a/xOpdN4IC8zBsBgmM7HeDcq62gUSQrIig1hjncyPPzmCKyQBxLLH37QbqMf8HMKR1KIs1p95e
2uE7sEcUpC23cLtcn0Kx2OedfznQtyaRLmZkHVmaK+YMu4NzLiCopmzWUhQ11CxHNSyetQ2CqW2W
G0B/iMpDCyKl6GAE6GFu/xTHFki9y7X1clLCCfD9aXo+d1MJhPgeFSHT01k1Tndi0XgU4wPnlzzp
5QoDoPJKiBDoGWZf5Lq0Phd6XMxguRi+tvMppSK7x9mQnW7Bx+pcugqYwjQvTGGwucuQVRWQ0198
gOw0fS3ln6Cw77a0AhSzoBH2nv5b1FyBtyVmhjReIXj7Ml3HEV/pZq7HxewuYhEjs/LmORZbiNmY
LobyuiOB6XAMSonkLZ31eOXfWcaypn/+Ou2xXV3moTBzuI5ppZCdElVO6vbsEAGIXloqtzEB1Jrl
FJjPdRfGHsrPsVV8P1sfp9YR4tBpskZ+4R0kHUj34wsNc0R8hVVwDT0RujYa1Si2FKIYGyXxg2qN
HqryObxvNpjnwEB4oXGhC0gH1+jh+ACoQR504EUasfzUX60kopZczWvhAe0mMooUAHPBMxeYZ8Ua
sRK/+B9fEF7+xexXYnfka8ErJRmfP6D5WxhucXkqiF20+dJ8+bjUtDC3k/muFopNLeHc+kv5QbRG
i3qqjYEsF/JNdL1fInh44aWWRreP6JD6/MePQXwQrPxQWE+unqcNdzrUnioFipqzm9K27IolmEx9
2O3q6fYtI0GlW8mtdnCsRcuXKuqTz54i2ltzbQClE6IveXDU+wp7WMEe8llSEFwg/KIOIShX4vs0
lmtuwrV6HE6cNk1rBL5mfuO43jj3K+9j2Qi0E6fMUuJuBSHpSST0gPXAdoc9GOLFvdHqgUW/r6HW
oG0AFbgDEw3ms5h0xDG2+M8MqNpXQrf4Y2jkDmst2D/JzxyDVSTEWpLTBWpAsyalQSWALBZQmmD8
egfTgMo23zSzjkKGO26nAM+Hpmk3IBawRkNdlxu2MKi4PtKKqA3szS1CPx8hRK+bbbBA5hazVG3/
iilqWE8pU19SuHRGPapxm1fv6Q11sCFcKE+h0YDyE0sdGxLgMX3ig8+48xsjG9pJeMQFXA3OEBI8
dxippa+YBws7Z/5GciyzAkVOlWrWTggGba/WhA8TDIgfnGRtChZjAbt8GHefDNLGI3AQauk5H9r2
P7jurBu1jy/zxt+ykouJqcj45GlXp19OoiZXmD11BdoV5xo+yGOJLKVFmFz2dJ6TVUhfSRYhqktK
Xx5Rne9PFHnj6LDdI4AYizHuNyfDDcRNUjjta/JH+kAcP5Rmm1jht45nuycKQwH6jeiOVQmTvdPi
G8Bi1B8rY7CJxtU+OsiyarHF00rwMY8ctirkZAvq8A0RwDN24R2pQNHpXzrn+/SvHFooVeH+DNuf
cusv2oet022mL+2YRaC+ua9/E/I7AbC2JC1wiiZ2euoYkOZqqklrPCElP6WQOLV47DopG5eLegMC
xCmtb1eTF8Ju+ODjgfUzPEaTs8Uj6cTxOEHecpNhLgwfre8HlG2YApiuWoNg61gC1LSLoX1Z7bkU
bCOyGPvLqjBA6+MxmZB1Fbo44FbJEdCLfCUvR8E1z1ZMkcYqOXA83PnwYO2aoXxLGZZMAbeEZSLC
6IoCiMIpBqC9V/29GbKqmgj2O8/sh/VQ+SUJ4968PbWB0fJI6JqFlrn9zHvMPCFbIjQrhQ5QuFFe
GGwnnnUceALdYzka6UUVyC+h+uNcTcbhpxhbqgI4CAeWJKAff3wlXecyoAzY0oTvVbut4U6lYZ7l
6JZoQEfNLuws42Pw62aPcYlVgWJHN8FWmI5dsWBu477CNI1zp27L2mRJXRNPmciJj6Trq4BVJK2B
zagZyOazVoLXXEH0j/A9xw36wMjAU4P0TX8g5MWUeqAhxVFTSQOTOMOW6EHbDtaVTI3KjQS7tbZ7
lkBFZlPCanK5/w84wAcsGoxhdO24Bla+0w5Oo/9DjSr9Pk/xQhjfpvkOaQzU9RsKLZypEqZLLRV4
MF8x/nUqEk44sS75t36TDZPplkfxTGuUptf98eKvinEAQCnq7zu7jQ68r1Dq9Lz71YjHciv4eU9z
vR2HMeZIid2XPB1W2hXXdMuU/gLSEwmHWLbCn3Srdxl6ZhSNP91zMcBqG2D44htSfBm1vNyxYVmh
EzdBofWHAnaHGi9OmvoSn5xbgNvMDX+iYvYtCHZRgq7xZXVu2a1lKQGc4rfl6w8YQ+QUCRW/vZKP
2aeo/PEKwQYzTWuEkC7fHZB/OfVX8qX2tEZCeqHNmcVdPkHHTKZQzSeoxag4emb9Lmqv4UDmMff7
mil1zW+FPnEkQXCt4VP7EDY1JLckCG/IGGSb/GyjpUrBI8YAIqy/MHQ0V7N4SHZM6xy0LK39tlwx
RQc7apv3tDdBgYfvPC1sa98S2ZvCARGQINEoo1tqyHXjQWRUWiDTcnmPL1p3EgtMYKLKk3cThWKn
+F+22v6s6J6Yg3h1639NHfZq0zF6y3MbIZvXgTBGovJ/XdK9sosx/VqQXGVe5aP2PpMc3wbL/Q01
tNpqcOoNdwyziGQibbBg8IcpwvNDjZpmsH24e7oWx9IepJ7E+dMlq58EvCjSo0C+5wOPvxY9D2jR
p/TuSpW4jkdD81bPe+XQqX5+0xSyZshXto4PAx6ylncFpRX+dkqkWjWy8linmc9nDWuUySOyKHFR
XZNTgdr+wsvJpzL5wcrgl1wTmzqZTyJDkVasFJb/FtQGi1q9kwYKoM4xAitrterBXNqjtoDu1njo
YVm9eZDJfOflHdtquiOjGQYpTtApxb1aFo/OjpOwHiOxFTyEPKFAJKXLdaMVnino5aTLo329SGzz
QV8JDDq/5u/z+DHDdt7k3WWGqoaSMfG2c8iLabvT8pfqc5YUiMb9GqfWUz8T7gDKgErB+7VTlvaK
dWUBvFYuNd6izb+vy5laXS+RJyQJB1oeNWqdbpyHem8mDIFcycDQ5AaKEcNFBWlO0wRqWmYs6o3e
jcDmvFpppN72z711z+s+bWpeuUoP2O0SgOchesaTsa91ewsnxBkf2z/fydiURs9Ot5PvFtYsE7kg
hHtq70UhgpNF0OA9PGOTvh9ZPnUMP8s+fvmaEYOBsoZoDFUYxxRTBMuGHpF7eGEuwHlb4kSL2dou
KE1A7ee2UZrm11370ECxp78qxnjtFCxw8EcsZxIX/AMkQpgW+7LDbnTz18ANCrq3sG4zg6Ae7xo8
KADtCaPfhCfhyyZXg1quG/UQj1UuMYizTI+RB+L8GppK3wvfVLQ/B3mSwemuWHndBXHdyzRKP2Jk
zpAxcJYacaMUAkozY10lsmd5sskSBuBoV2U9Nb1BNXyBuW4q8qxe2Ql/nYjlEJ2/1s3/d/PJP03y
vn9q0HJA1PUmbZCE6tE5R3yZMzH47w9Bl/v10V52XLfV7CiRfcVGE37/uIbgXWJ91xbPNKeJRHeJ
KjnGTkNDeFCbcMbGw5xL+/aSDYoJaN8sPNlzppvWN8ioU58PleugbZ//RxhnfrLCLRbkl33SAgXX
ksxF5a4+EgubiT+5XgcZmqqE3DnHJCZGmmI2jqJXnbhGOOA/rHxqztnScGEJSO8JydrxnHgnrS2a
t8dzj5/cuOphzNPiEpnMPfayBnbWoKjKjX8s++vetUhDHN0LV41Kz0lwDVkBznOyFUr2SlT8ATzu
ls+2XuO8crpE7rTQSpii0sdX7sGbplyV9yLOVLlgtToEtBraRduS+lRHY6PLYdLBJ/hIDQcKsPQJ
vq5xx5eBJQlSfrLlV13+4aGPwqPpK9D74LC829wo/7S34gONbA5PahLtbGyV3EIUXirCBZaYQhb3
S9mp4zVH5Zo+a5YnBoHyA5TL2HDXMDwWQYj8cz9YOcckjjtIprMZPSweGfDZuFCASrFzB0PW5kIe
m7DkAiq7GBWt6d7+3PKKPOhJFZRFVbLO8KWZ514j1lKOB+7iycmcDtr9mMkNw5rgmcJEXyDtwQXP
n2Q3saF+TrXWTBt22KOEKsLeyqEJi/dyWepd5bWCFXcpFBSWk9R38YpbASLjWoWaFuKcod3O+hQQ
iiSy0+kmEw8PhQpXykLl7iShlv6QDUsxTxDosCCmtAEjqdJ1GdJiyh0o38Eb6z3ossvUt+D6iGnK
Kk8jRAX8yL03MEheYkwX3/KWkuZoj+IimfHn2MpRR+O4230fNUvA6QgfTGrWIudVKeltCSG7ty+5
2q0SSLkhSqDAFrlYam6Yu939S1LmFOm2wAMnmXvhFfIai/lpFfWa2L79UNp3fL9fSJLtQOkkDQyq
i8oY7ipmGVaFT9r4VQYfiCOAk7cfxJI4Hg+RbvPsESlxBwxQ7t5YJbGU7OH9LybtXnryYANP1EIk
R3vHVL6wC0fVtX3oCp50BGHcXAmoN39c9ki9X3WBNTBrhc9fWIViZcbCrqVxoJpr6fAxGCRMRYKG
m3KFhmqruAqZP3louYF9GsmuOBHaFrFyzDqMtWfVuF+d2aqFJ0tcVuWIrzeShkwjbHqvgXRx/11Z
+c7jrQM58r1XkDNvUth75T8U6kkAeZFh12Pxly+xNzAmcbgyjd6bs2USMhtwxOK0TwAcsOXEIQq1
Fw2kVsm5obqAYmWfFDmSBFBZNV/Ll+FhA/29LMMdu0A23uXqRr9fq+Ga/fEdRqWPK/SlR0xPvVtx
XN0I8aFAricJ/vgb3W/5KltdUN8EhXlldEzd+Kbhf14ti2lOGKxu94YvpKFr0uDmZe0TDdB+TzK5
tJalKsLh86U5pPqIGJPO/GeDgqGQ7qBnkeAW0ciQZnlGDBu+KI4pSjGHwpsAODe540W59H4MG7g7
UY3/Zu1NaiAyG1cmYZKeMp7wyuV4sGII141Jw7tRX2U7pYYEs5tGHKfeue5QF+Y6v9stNAq/7WLP
kWu2ZhIs8TDHyDTbTCDcKLezoaE9RCsRJKySq8v+oaeRaxJuQPlgiBNB27SaUfxURhXILot9PCQM
PWjKLkuN1Qv1PWWrHaJrWgKncLOJ3ksGVikkHt/9YZOfPlU81+Dka58L7t3WIeLvGadVRwYrniTt
zH2r8CNEcfJ5QgKJ98D+rsafFHuEhvXmAM76XLfoQmrSnGp2hBytVw9GVL6m/KPVIAthiKZ2mgZJ
72X0Tnek8Xphs8CefQji70Rbz+MHYUV93izRUoKiLrj6JOjGIwc0PRifaBLYmiBxDFekbo3EjFUh
LlbtkwhgTpHKsrrsokNDI/Iy5VDG9Z04JomoTkCR+XEuCDXHmcRAXCf19xcS9FZGt0d9wLPMv181
LS4sOiuH1+Rz1q6UnlR5WWrl3DVsmu3Xs7xUckystlvZJ7f48AI7VvLS9eauvY5SmVV3p3z7Sr/4
em0mHVlxaPEqFQ/b2MIiYYuvt/KSD6hwiz8Kwdzu7wd1DwZhMTB4CtW2DEjxOVQGcxsu+PC3z9YR
cuT+AemxvcC+571Zhk9dg9Gr+Omo721ZHPLNXYyGrpgKnzQsTN4yWvXKzY2RCzRTsUmiHpJp4z5A
7c4cFi1pmIEOsaxr6G4BQIp6SP+M48NIsybdFWh5AdLPKVSwVdaoyvejUx8B0q327B6Z97RFvKoR
AhG693l1grQ4cYfn1CGaCclIgXEC11FMWSDhA5IzoYcBu2MKsHUswWeUoiZedwWKS8mNDmOqnlPb
WYfiY4NaWpZXZ9dSHMYHpFTdE2SuFdP+Jt1glFrSf0vSxGl8D/CqhRh8GdugOIQ9kuSh6Hsp4wPN
xyGC0pVqPBw9DBnjHfwlQseyQ5DQiIMNTPVeJ7Y6P+xg4Ltuh619OzyyCFBko7voWuBQ4Wwyk2yd
DcrGivuWKAQUpDLeANmHBuEyruSJKj4oLVuvVNHXugzB5Ykagz2xsfl9WDerOXETFh3rZ8sLcUD8
psog3FTU3qt4usYZKEEPdI++x1q/RHn28fr/HuKrlLOePeWuRktlZekp21W8spqwlvchTCxdZpyH
RjJKyUxtDDH1ZY+LBVOdSKFuklwY2rCtHw/JeVglLO4ANgf+1Cgp2q/mOKj1T/NXqBSxpfGWmMrh
nTgAr7x30bW0Io8dZ5jWIUKVQUc8q0kKjEuhspBmMSAZSZ4KTwc+zIdB73zzu20qfbS8lG7HoZ9j
y7QE9vUK5RhNR3CzKaQPKlcJMRmmuEr+X5u3eT+EFzsSs6zEbfgKxgdt+grqAvvjvsBKfmZZVGuQ
MZOjT3X8B944fr2xepijlhUYbNAVTYBKjCREIq4AfPpP9TvXk2rtzeTmlRwzW+WHWYDw19r0i2sa
EJanDS3CwnyBaYVzJtzoG6N4BTgUy5LIz906Rzx+w/NSrBDgDuDN4lSEQGnHNN2WNYkZ7XOXNTjI
YyZoVsZLvepH0dHNtP2Sv6O3LHlIdv/R9uTyNjmYN3UHxQKjs48ip7zzyEWeju3Bhxz352iPnCq3
BIWmzMJe/izH3tPQx+x6MaRrSXwqQX9vrY1UNicJMvYgvbFpsQem1wXGdvZ4Qrmps2T4QrKkQwt6
3F1IuEbXG+XhKMZhRVD1zYV8DqjKGlXLyXPsLJumrhcCO+VQnIJw5E4ig6srLVy7H368xf/MTCcC
oZy3fzCR5WoRqNSfo/gdMqdds9ylj2h4R7mgQZeEGvmxfiTx+TQFNEDUIOXiKL1aHT8SWYr6PawN
wLRLaFsoyWKLkZXSTZuS/kj+/2Fo8LhgFAoHla4HG0IPHC1O1vDJKmadGnyv8xn3oF+MmVPS806g
HAY/494EE6lWOUbBaPOzqsvvVNTR3trjLK+kCR5SOS8ZZkXM+lEg09mBioJDO2ezO54aAdSyhAvh
u17SirMTL98r2X72lCAKr6Ysn40AwM0tivHWWa8E3N4zkoF1LXzEr49qrhTUKLexapcuNsEdkvzP
9Uf07AvJfWb8sZBJi0oYAZLwUUg3nDqIKs252+TTT7i7Bq6EkGu6hKebpre578rRmRAlccffk9xm
WHbqguJwH6s/rwKjYlKinasqlTWjEb0P5xM4Y6u22AMThtH+513yCOfQWD3qCwq+D29PySIvo/jx
UOOtN2meyNeYKqNZOz3DHKL20plnOu1B4rfQCIcZOjXZz6dgt3wHsWBEbVN/5dDsdeiHLiwq1RK3
XroOBzyxXtUcxSPoPZmrCFwgQFhG53kExFsjXJI2CR9bPPe/NUxW5v+yEIszLoUJMWH5ZeWuzFZr
Nlkb7lumNwwNq8jEJxHCbI0OrzADMw6pNfd2G68vXeEZmTqtanBVJ7YGIRddLl5rFwwfh9B56O7J
vUfyl/m1IO81H1kSPUXTg/kzAkYp+jBnAQjd+IR9j/U/qi0BCyRBFva071pgjKXSFyeimH1ojj0h
TYxq8QoR6HJdwIJLOUkWUYq5Zxs4jpXcsy47l7ufWO1uBTXO0GifnX7Lf/vrEnyMX+N7PzAAl88k
5EhEYO0zLR1G8AA7orVYLNrS2zeIIggWuJjri2KBFUeiFoF1OYYhid75tv1jOZ5WruSg7NmR4TBH
sQMjkz6tBV4ixz8qTNJMdWseF3KEMekRL7AO9I/6T0iNwI8T4eX60BO+16uxAqvMoBcOUpPZyZAM
mzu5b69AQYkW4FxY1Ur20S5L7nqVLEiGjmd//ouj1O+vh/DA6yKo2e4K6IKroiTVUOBdHsGE4Zp/
c5p92QtQwt02oB7B6vAFNJkEFY+D9Mlq3kV3q/6qUTCPv6gtTn8tt/yONpkE5TuU3/Ux0vyjY0nW
IL9sso9qv4tqMv0uSEBLBXQdJEJXtxfAkzSKn31vi8Yr3ldzlpCUEfOjpZF975Z67U085TRkP5ua
qFG6P8013+z8e4gSlx/F22zeXCvwHWJE5rIWf+cQGzJ+Q67bHoyR3a4Htoasby67QZXsFxtOHw9x
WrIu7B1Y+pEXFzD1DxticwmGrBuD2GDwDGGYcm84dqNSjvITUPqw6zTpU9LrgVe+oKy4keJn5C9x
WqJAaJvpn8oR29y89j/VX+LutSGd65LabRQodNl4OGdTOAj2Oo4oQ8Oy0oDVp0RnbDZ5xc2riWD7
AJ3NQJ/supQwIGoeAOOfwTi0YCn/IOOALHxNsr5g9aNQ5rLiejFqnEfm+FNZWBZI52sdXz8dLNuK
FRod1Gr60UeEX2dM/8oprE8WAP51B/HHPk17GPks6fwatHkbymZz9d2k9lLGmvjk3ftl3E1mg9PI
Yr9k5ob/94e3vlWWFn3cS0t1pO1wTseF0YybKEfRR3avfe68U+KGoJuNNTH1Rh9svgVTevw2G2O8
F6PIf/iO2zyjf7ulw6qh7G9DDLkUgomTm1qPdsGD+09q3voI7Sf0lY6nd58QXbYwtl6WoO75DL7i
s/oNjz8eVNxqRf5UqvZeLYiwS5QZunC4jqohUE/w452HErjv+lQ7ttZf3jAMykOdns+y7xsi7cU1
xwmrA0eJuygzy5+hhaXdT/GawDVKTmnbH+6LlPtu2jZgf7ZwB6JcoPfgLiHZvLsEREvi6SDtuqLF
FyktaDqzX4qyqBo92vtWsjxxDRrNB5XFhpv9mGgnAyGxZxPjHkJxOPQyVXMd1oJlO/K3WgMFEp6q
8ueX2wD7Dk7vb5cz9u2EIVsNnhGBOboQiQxSz0yzc9E988/4OZVzrAoRKBBYsA1ysjztCOz/WkK8
7IoAceY+7oD5byf2dZTFG6vXKjPmwaVwpDth0P85mF2krG5ACoqHtaA0HT+qiUEXur92pgu/fNJc
jBirf2OPqolJ8PZgq9EIfnueQX+pbyOlwFWtoNkNx2jvSAj7ihrAJ0hvNYo1VglTu5NWf/cXkNAR
kRuF7yEV4GAgiEi7Ni0SQMzqOfgWeWeP2Ui4fEg1pUjIeLdJqLEbLEl3V+hOPPsMVLl4VGHB+P0j
DFMFD0xJ0G2mjIATMsXglWsD7BK8jEhym7GxYVqnWvswQVc625LPO5WZHbjLhwK7X3ZLS296Bau4
xMBTHEnGtu4TCH5LLu/hq8S1eeu+SyILau2xxybYwM8lgc6eV0IobrwbsEvJzrzXRXoFIj14ghO9
rj2Olfdwbo8bFQRjaG/Cqa7h+DsUOzScvLvArJ3fTAuNXl8xS1hoLhpCCiRV96FvxqUJIIkMJC3g
XhG2/KqOES5rXsb1ATPavYIBNBTP9C9apjHhvc+r11B1kkNhbuMy6uwgcMGp81yi1V5Fzc/SwxXx
nVzBBFe28nAsT4HBQFSnwt2ykJOt3IZyE+s4CsJAEs0UtGhH7Ow5OVmCnz9k5hofsfuAowInvnKG
TdetUSHToeZIZ3OC0NJVkXUgLWugvWwB+rsrmzsOgDpzlAzqeFJnEZei69ovuvx5q0PnHQiL7dc5
sTANliAlTDwir9ukF9rCfI0XyyH80rQHTJfvQUDAWSRYepj+zrMoXUHY8XSvR0RJajN2V1rkad+T
DG49KXgnfPF83rIuu1nAQhZ208lsyl1GAoyMUZtHv+66B61h6V9JaMfLuRaSXlqk1ojwH15EzT+r
OafacTOT8lUW7/3crhcK47QMvaniQ7uOC5gVKdV6s4XQSQfBV0hg2TtR4HMg9hlwCAxU19cSmjxV
YLOTz0cGBTY1sgG1ysPEdaTHZeQQnu6Kz56aRgyM8nSOFOvsNkRWt2kAGTwtwRlP+rGpTnXmWlTS
//8NHvdGvMrEbgqJvhxBmQ+SNNykCfA72exoR6BvwyvJ6+jwwimN3Gw13tg1QLtMpXpfZiP8ddSp
azCe6ZllkZLd6CYwdTypzl4mjEZRkEZAvCpkRB2PQvnqEOHfLhJJz3YIOuJqLoGqW8cR2eF9dfPE
FqQLngd9axjlWCMtkXdsgcHiLrjNFpFyx5KVqXUI0k4n+Nl8+X2bH1FWEHHiyoKkClV9gv2RtLBr
e+uTPkBREaFBquomcNqEUVJOmkhzfy87JtO+lYmKE3W+C96SoBxYV8lKfuowUZk6vXqYACf792Sk
itShxD53+RTfSUc9MVAnIl6FKiWLA+1ALsOn4Ju3c1J3b/KbXnkTygrxG0vlnZrBaTmaf3hpkKmn
B/4/5AaS+jrYvXEQ+zUvSt/aapHHRIB3gVySb4IZM5QKzaZQogXcnP89yjo6/PNWgwM0r6Hd2BzJ
OKm+mKAYyguCNl3rlNhkxiuSG+T4zLfSZ7a2Itt8LUtn/3fIfJx3YjOaFqP94uATykf7AQqBtStK
VpUFnmKdLwbPFHx+9PYIaO+umoIfXL0Z6frdQg1I60JVlC7KKJH+i5n7nEd9pgxNm2R03ZCIhZ4i
NF1WjfobAhqtz4w/2S18DRoVaidD8udeus+1l89/7LXDEPR+Qp9YTxlZDE56ajB4IJLM62LgOrhi
2JtGDsuHX8kG/BQBiH844L7oBO4f2lJOQtjR5Wyb74CScNoTDCC4EeIclvsQrH0OCyIPDRIDTIbD
ctW7qXqyx4IR59zMYWhXLJMzBFktoFJsslW309kiSdGCp4y5g3T9SUAafOgeT2/dI0d93gF1kwtp
OuKvKCpi9QQnqhkrib3haMou1fPrXB9zoJoQHU3aYFnFgIOp0J0x/v/35MT2J6LqUc2BMv5ZtNpn
rrCjrDAxKuXxJNTJdrRFm+B4MFRZefqngssNeaExKrHqEdYGyRin7qGbA10COeZEAc46VIhmYL8P
xtp87uIU8nbYeRZV8IeR0b/hnOsFv71SVtyzY3V3eZPMEqEt7MwBaCxt5Y3GCpU/3YbJyasZ3fwJ
XaGsxRoKCOvVTQXTtIR83MWvxupkOwMHHHRky8N3U64hkreIgFQermcfM+wDSekEZYgSRYVrlGfg
XL6fboLuYE6Ivq1Lc+YaQVvE/n28NxLSb8MRzrjF+BgUsJUL77DvH6iaAmIj3zhCXFy3+lgLoNf6
umAXmsBszvEMms7sO9eF8Yayijo4E9IV7k5vdAMvj5iTRwMrzVZSNVbAtgs1Zk7VIDWJLJypP5WE
r+FE9rYggxVeUYNnmw/Iu6QD7PbPfSY2skZOuwTCF7Dkh9ExrdS/QMcc4Rs9cTLi1uiZaR3FQE+U
n4DdsHLcJzcTa8EMRoPjiQO2K/40TJJricVMb8RKuILnHj8O+oD3CoPDAMyZ2gUtH7duUKL0UMmg
190JG7QwSKt4nxfdiDX8fiFihrdc5dqkIimGSLhPfELleNwemSn/97T4qkNtWXEnJY6LwZBZRYQQ
e7UfQPro9MQvsgZwsWXRknTLWXOn+hojIZmxxlz0RR6As/WMqqdHAek6Q5Iy3vXLexatU8bV7JGM
W/fCSoGck5YcUIDggA9EwJ4iLeIaHE7ZGoPSAXBI9joiycnys1bdFa/qL2doB0gWnChFniadRszP
84QB7azz92vOrPBydzJBV5RNjZiEGGt0Jg2BabcjuwG/tpoQL0Zg/ik1AfGndHvsI6DbocgWK0CM
FAc5GBRBJk1fwJ7hBXx+CKHQcdJ2TWjROU/brzbMRqLltk2yd1J2d9fbhwqQ/MQqTBVphppFWKmJ
eXfoyRLCbSOCHlNXIPhsAq77sFW1N1IAnkYlzBH+3mExT3t3CXSxcfwPFRKz/dr9KCNJMQTCvHHE
Q6uXI/JUEwC1H54SCXHiLl1ZKKPZQNMhzvp5c6RSXeCriyUE1NAPbxoA+n60RVtH4OuBPwl+SnEa
KUJqHPNsTCOYQ5jCNRf5JyOeH1G7pjKOUzS5AIGCSwq34rmEYzzqA78RDxldQQZKtsvbo2kA/n3e
NzjFY1hH2a86XO0mClAReyY+i2fi5136kQyAI5gz8oD9XXhClpvJXoHliCFclDgxKSgGsbeaxFVN
xt7Ium48eW2kbwQdG48TuVJNQTFoS4QgcZkMWUK9BJ4+XBRW3sMSunLmi3hbEWdgWvLaomLczUVZ
JtdQfhmx6gM6I1nHz0whtdMtSVeWHpl+UNjfU9PGfP5rovOgimt3wKYDH7iiXeYQ9aob6Gydc/BK
9R8LnJ4MOOH0CUufChPUbxkxbL1Pu7Q8AXvIUgdLp3+VR2U+dMfo21GEG8AFJzpJz2YeE7IBtQWp
WY+MwK0RROSAkiwnZLTfqJ30Vzego2r1AHbc9Lyd1AuFUv/DSJildNM7fcqtxGfYlkaVFDKleFlW
6jqELgTdiexZ00CaCKjOHe27W9sNyJuEBCaYs5qmbpqxorq0rAPRjV+kTNxkkb9iFsoeRESdCHPx
bSca+2lTbSrF8vuZy9Rk7C7rw/3pt8FZHBiGzwzdll2aukHiQFZnALVU5TI2OHogPjZKeEncP8hK
Q1OiHoZnBfnt8EyU/DFfc5oGuPiUqrVGronjybfJbqjihvzvsaFOgy8WOs31zA2FbQ6CimG87975
mXTB/hxxWnllUymnubiER4dLz+AX/3f6J/LnZndT702+HFf3DnQeW4btkB4JHZNFtZtXAdHkyheJ
aahGCz9Pl0ZzX8NXVuFQE71idqhSOGtfoOqge5KQ9BMuxP4OpH8nC/Mo37C5fJQvs75lQev4Wpd2
uvcKzkzx7rOqzTTC4p/WsTV5GJBtTd87zJjXqvpb0udldS6C/WDpuglDsw1EmR6vC62/64Col5Mh
1cZVQMe6hbcK2V8u+k94jKQ9mfdpTb2WlIeL8e1CEUMrmfa8+wB3wszBHxiu5flXP5xl9XkvGd8G
F9d1AmsJUW2uLkIMaNVPKGD8B3LSjBQqZuEP/YnvTWN1mT7a87FW+ARLfJg5gRKUI0QQqbFgWGL9
p6Z+3qrP27lBY4vpUcN0XvPP1AZZxtKkXaj9G3FKhs0DIBNVoMLZlrN119yaptUJbs53Gr7+pFWe
OOgUqsQ0rHSAjSa4U3xN0H3G0vMsDCaQovfc5949CJfFr8rrzI4/k+Rwtp3EVq3QlvtSlp0Ls51r
6ESwBspbFxekZL4We70cVDp1bFcBCHw9PbbNSquQA9ZFA7UNO0grS6nbch/EM38JMadXVNqX0iqI
VJfNFuXbfe9MZhIJtNz1jubafzBAZg/c1VqTomu+2mU2+nzvtwNxnV0RMnW6Q/K2LaYB/C+YsLPN
R4FVGcca8VkABI/sK1LtdPgP0lq02SdzH9+H/eubBKqIuvcZAccSi18e1XerSdAQySxGtVN2RdWW
ZbRFWr0SD69MtYZM1s8b3Zi+1Dz+qJbhkZO80Ek25lGKH7qnu1Jd4MEBQAd2c3+tm0ybiT3N3Rc0
Bpb/vPdf6gZuGglZnJ9DiZPLeNd+ho5K+nT6PNbDXj6VbQO0P1hMCICnXERNkoYX5XArSxv7//yx
pJH7NOpNw6akDCOdCIkmrioZ5INR0dcWLF/Uty8X9k4bh8WLiRMzmTDEEDjNv3KgKcsHc3YWxMbU
dCeHpf7MtJbE7eSsxW/ikQGlJ3Bmx8t7YTVKuEc4XqGDTcv9oanPOJLU1btxE0jnPvvSFGkt189d
5iKJFuyupNBtECIg9lY1Vz6ou6kE6/oFnu1RAjF8cG2/SaEnwNmxkWaW2rjYr9Zg0bvw2pxb4mUE
0ozzL1noxfjrKG169RUZ9D4jHDTOGofOhRU4NTVB6R8Tl7bjOnLln1LPIQeqePL6SU6Pwn3bAmDT
FBxXZKfGjJlAbYKrfXWsQfk994Qp8qKeTKpM+wZ03BpGf3fZBtwaKnhLzqRl/3XwxS57v/L92Zho
mj0uIgVRCFcIUwJpCn5kLs1cBPCNHIr+OYlLA3ahPiQ0X8d5lMIMISOQ5TWvq2w6abcxWROTHR5h
BWU8j6hQ8GM1OUKjnVbrGLgNWCyfHge6EuUX6Z2UyA0yOvV+MhIWKdVesKUQZ+gjDZyewT3snSGO
pDyik5mwj6/Gq08cR0nmMD770UUXW7w0H/aSCUHUfbiVfn4VF30bOa1YV924IoafX6nirilGUPtP
QJx/72UbT02ndnhVsND+CotG/I6qX9aDedsMyW6jEhmvEM7td3oD6QG6DWdB1n+J/yUKddZ/zmsv
cqZkbeFkRw1d/8AsNWiHKXpfoIVuXf2sCUr8si4nwbFt8YIUBTIbmAirW11ObRI9FIg9x9T4LivK
W5ddK51OenyGkn2Qw49Fefht4BmPB+DEZ6tkC2zHnwnzwihkUDzzrGvEvAyNklKHE4vW3MXbD/qP
JdWR1ASIx4d0if1zFfCJ+3GnEFZ/c6u8HkMhYMk68j14qotZZA/2nrzkrosy3MfSChq5bdmXB51F
D4eY5tMQqQkpHhAUeYqpgKHnnBozFhHoLiUBNgmn+ZnpgBxYuIqcW9pxFbFG7jUEN+kUbpbH0PyR
Yu1Px3x0lhhfbF8TU7xPYqpqaipNqj/u158UQWY5xWjmKqBgyO7EoZD/PFDJK75LitPhsGCo/bl/
canrgOf062o3Mio9+G3/YfLOyURUyCBZ7FHBPYOa9fWrOAkYN6bIR8Aucl9lteyr2omIpKUVHOmN
+LpmBQkIOC9xxTVSO/mg1+tKvqK84guUD5Sz9Bo0Rm9GUB7y5LSnsWqE0sC+7aYHaLW/uPKsBkCf
KOvTVYr6Pr9cPhVjuRysNJ20nvb6OiMErBfGYzV+LVFeQGpAVOTCV29MhRAuTXpHjlKpu3h/PW5K
nuW+EnGRxSh8lRsmkm6k3e6YPiSI/4nFJPgF4jZ2pdo9DhEqGudcXcB8Q1LG6Eghodpp4A5LtuP1
BX0I//R6WGEm1KWnNFikChxpYQRO/NjTKZY3yfhE31RwA7KOyvDHp0pAL58Lks9S9H7pC8g+FPHq
e7e/mEGnKrPXCn+O1EcqEVkK6M391juSfQe22H7MEZdb/uU3qHzAQidtUCBT2sVfUzYDLkkk8I/R
zfnpZu1FRPvcvuq7yBGS93IHhFbpDT9rNmtUafOFz47IEWjXlykpd2qQ0xgGTUa+YLW8VpBOmr8T
7l6qPEyKHINfjHMhqe6fdwb3LaO45UqX8whFOwqcPSmHQGt2I/nXX5OJjtJBjSJ/uC9XG//0Wc/t
CyR3SnguyTjM9dZQ6eaHdn5Y7gjGUdZkSqpvVurODLgTRs6wqGvZEFFwXgwjn+C9kX+mkWxwMCef
Z0KFFJZIJMixQEuU9MwbXWAEo9iWARi6mnKZR+Ewhglll9lCBN44fuTLtjDs0cVikRVudnu0lHsd
PoquWyUfs2K6oZPkP49lm06rov7pgXdZiuYegJxYvTJSVwUxHrsxx97dr+/v/4MZkk4HcqYjT7fJ
cnDZrodPcjCLHV6G3Ms7C8Q+lTD3d7jDgxGzDxIY2UAhGjzFOPhF4BdtHR4LNoEOslfsQ/XpTHo4
8jMCPVIpQnylp/d8VchWBvRdTMG6R2xjB5qO1CdHBFQrOiC80hAQs1Gs9MFCKiGTwGQDnQgHmTsE
2hBthzxM/yKlv4N++RG6kEu4UlcaYi5OycK/0VG8Jw+KlDImwhj+JwsXeRn7EEe8St6D98f1LdQG
bPESxlncTihUU63Ci+Yz4Ozt/36qrlgRwPEld4FwADdzLmeUoJ2tA4aOaLYm0DBUT6ieBlEazwIe
jRIkFDgS2k2cw2+aDWfKxldoPBtmjTCSibxL1d0ZIrylQpUkP2Kbulkmuzi1ZNsWQ0bqe8+Ehbit
Q1ZkEtku2pMPAh5tnCBKrLfQDFz8oPJG+Z2v95bimuG3HGAJupV9GLMZqqmH8ZxD5at1Wd9Jn6d4
H3I+2mAHbyXDPMFRnYCIM504Au3ta0QAON++Ug+PNnEgCyrM2mRkPqBgZlVI5WIgMyZoF2dYk3tT
BaPzpDaYXYzlL1rfdFs/6yPoUeueDW5Vbz5ib5N/xHaBjK8YMsSz4ikA2N3ICQQnRo/35KZyKekA
L4vu42Ud+LasYW+BQnMeOe9KotfO2tl+rSusj2vK+AEJ8cnB9ru0o5eeoTMbxzmhZe+5pPU2EyuC
kaFeoSUBBDrP4t4ja0mWOz0o8R9Uhg6BkEhPY6HOt/P7qYIgACC/g/amkQNL71S9yARYr1Tjrip8
z5ngGBzNAvuF7LXeKrYe5WNxE6l5aHOa9a3zPhX9Pv2MF1IRP5aL6Qxh4d7F5HCdVRp4mD4f8rkb
m70tqGu/9J7XcQJ2ZcDVii8vMqgeA8X8Bi3arMKXoOBh2dTYNshEyOGaO4HQxRIyQcULzRA0ASGy
G6UZKlzgf77kCLTUXXrbSaJva//yE+6sad3/dsVpWrosPl2dFZh70etnjpckEPAxMt+GYxiwZAfo
UOwygO4FNv2UWGM6AoB8v648JIRChPs6sg+JAtiwOv4WFxhOXJWfRSttVCfQfGXktT46EVIpZsnl
yi/WEoWBBDeg31XGfshGv6MI0fpVdgWM1Fvz7Wvo/j0BO7VLnLe69x8Qd5z+um34r2QdQDwwwp5C
7AWRA2t34Z2FguD4mr34r0aDUxh44RxryMkFN0OG64a2r7zgMiog9aCTLRH3hrjGZ0is8Suxk6AF
zqeErD1rbNcgAo6qzlnr6rOsyDDKe916RxUCKk0n3yZ0MiEYtnEoYI2+hCtx0HnuPHJpgoPEpCtj
/C6Re5Zo9EYtjXYrVUW5sMfiyf1bdegsEITJ266DgdKN/oUX6iHdN+WWl/nvcjPNv/bKnRfQx2+T
SAaIa/wk052DTiOJsKL0oZN8Z8vjNUma1OIdaGLItyiF7DM77irnOkv7ZZiPip5quURNK4fxEZO5
BWYs7eq6nhz2J1ku3pui0Ik379mmFUWVKu2lTwFcEu21ft0je51Xcn3Z/bxoDhFbPEpcZPKyQcqj
bXoyxxLR4OUUpXqPQ46L5q0QU0P+vvJz0zxCFqpMzWxrifguUfy5P5YmOooXml/uQEtI4HNhOmPq
QAVmc5iYQ/57rFN7cDHRxOODr7/xhoYZz4LIiVrwWIfaKY+K5RKmqxK8Z7XkZXYb2X3Uw7qV5ec/
SGHAbuWBnvMvTn4E8VQ6mR7OgUJfzMVZtV1CVtChXqQwJTjN2zza+Z7dL1LR19+JA+OkbqoBfzku
sSV2RPdLSsaUiIYhMDFS77SlFWCYH+ugWGPHSTHU4Y92yIrouKDLELnMDvAc6xlb+N5egRrgkaPs
1FgEkIE2/X+WatqUDJcqLisrmFSis3Cpcqgyk1/Er/LrxFNjjKuRaBBKZzti6PRTDPMT4NhCcUWn
Af0n3Y+KkuMN2ZIkQEcqYfYrSsw1tp3NYcqpbVW2E0gWm9mdR8spWiOY1F3W4U/KxHXKdMoISxWR
KGo0nFwDHV7WQbfz1fTpgkNW5433YX8E8SCsaHjtC/jB0IzeaBgBg4ESz11PbzqYauAqqO01KoS9
YlRmT6VndXaG8yioAkYgAwz2wgB80Y3DYgNGP97kzQTO7xj18ee7GHBF2jRMqchkcRvm3vda5LdH
Yqh1Kq+OQ3uNn1SQF8YjTJ4Aas9QhBswxAbngHEWn4xsFIkoQufivtGlcXEEUlvnKRyOWES+aqMJ
eFR4+rlCBCky8s3/jLQmNoCmTAeHVz+2nAvi5R3hE60TM4mPmxPcYY+nmX8zQjuZPlijPu5hF1uE
45HOKtduJUQa2R3qTUnOJ10Oipm7XQsX1K0Rtn11Ao7xA29ICeYpUmnzxmgNd4h91GGaiwL6hJJT
488Zrrdle7QF0YyX2nREX8SRLW56rc4odi1EmwO/16QVuuUxryAC54fOVFbAdqvkNwe/Q+Pf80RL
bRyaU0mvjsE5VKuvwvqkisREMja2/7Veh8a7sO8oymsqC/j92WYjP78RVemWdC1+JOHxrOidjwuf
kNvZMEWpbuBrEhZ/9OGQUpwrKoGLuIDCdBzj1qHCmVf6+IrnimTVMP/l3vcI0OqlQbM2AE6WE5d4
XuekGTF2pGsSBl9QkfOvyItWONXUU0ohyXnP9wxMcKRWpNT2mmKbWGVn0aG4254gEwkYpbj5wVpl
Q8nVCKJgm4eh3V0543B3sJmV2tX2ad8D1t7rufMo68Qqqjh+/3+BPV2aPbpyCsuz8wGiRawth2YQ
+LMtA321HtI3L1sMHwDXKpxXUUqMTQRpcS4lLwgSB6HLpj2JuRIPm9Xj1EsPAldiZj+tNuPFRqY4
QfwHtsv7DasvFff4ZtarCJcNVf4wZdFpDk3NhVhHopmyiqQd/4HmlAYueBF93Y1LfZ4x3oCR+h/o
96sfQxVh5Zqhpm9u9HjPlWI3PFxHNUIEU3l1aZKcV9u4lW0eeLz7d3hKo+MZC34I17nOwppU1Nr3
2nx9EaQ+SiG7H6mZzWT+Q1PIEsb9HQH51ywFAYyB1vHpgAx167XGSEx7yLaEsfmVGfy281qv+uHX
ugmGieVBuWsCbKeSwmEiHNelBzMv5JMoHgC7cWlXDwOSxQuKlLomtwf+k++yDIbKV6xs9HtKj/nb
fj7N7wm2zp5FLUPJqXIE1LD2YrLHgTD9rw+JbhW4vXJuUmGBzQxOxLF8uj4aQ6TiC01ZeHoU8MSP
BTrxDhNEsoTq0+TiijFG9T5owGJg71PZhhQ6wIELXQxki1k4sRT96nLbU8UbSJ4re0uXXHJyd471
OMEdfpDq0k08mAPHFjIlfu5H3daqM9M05reX57Z2UTqHMXt3wJ1pQEtPz6IORxXaF3xbsRY4w7tL
s2B56zwKSahQ/LcBETO/+FnQ7WrJalwg04/bvMLQZ42pvdpO6Sodyp5VB28cHbC4sNrNDybV14vT
yeoz7BdKxOd5VT+ct2S9V8BJt7yN8NC90GyUA+CsTpngdnSzs5i1Lgv7ls5BOFh4pAJM7/8J8I4+
VkTgA0NJ1C3iVGJJxCsvj82HsD5/wyN92vdEpn3lvwNHP9rJaTaZPzIwx4AbieKAcDVDmit0rzqD
daIdhf3Oxkc3tqQOsVX1f9r3QXPXCA1Wr2GEh9cAmiw8A2a7at6vs/dYkznTvvaL5G2xytdtxot5
w+3RICoURlVdc27YyrBvE7Jy+N3xABn9NjkuJaJyZ9CCfRxvge+rTtHYvTNvUAkmHpt/4YC6aZHi
bklEjYZT1Jl6wPsjjYTVpWnfXezFyeUAINVROraOqWz7VqAwagdin5qBj3vV+HaYGAhXa2FBie0f
JKmDSWzYE09MvfKOxI4loYWwHIGosbZZ2tjJpAgLmve3mMKlxm4pxNsxUc9HP0OH4pDdM1Eitjzc
3IYL7soqNFnK08tZnkK8/v/69fVCh84u2zTmORUnyUFCLK180lDNDs3+rXyH6WBfzmpB8r/OvjZP
BYpa4Vdeb0oztIQI4eZmLAsAmaza6zMB+Dnxxiy1Rm6IuIIndLlGLpMpJcgvxyRvy5jD1Be2ZArG
Hhy7j7t6noEShAVnXvCX8WcCtPa9d4OQVobrbA8NoV6BbOSrpvHG8GxqkmbKGJoXow5hfQdvyo+Z
Z7d95EGnrw9C/KOx+irjJelqu/liUgIpgGuTXRlNjfSuMWsgcb0mpG3X/KAM8Tk3RpF6EhBp4BEX
IUqzgonEM6Pt49ixprubxMHtsiLLGeYx248ZZY7JEoLhx60ZQ14oTpmgJyCYA6mxpIvzej6ULiN6
gQL+Dg2wYfu4yZRKX0sJRbnxRopbZ5tvl9g/f1DiHec05kHRZueL0uoNzuln1y1UDk3lRrJeFv+a
N5YT1lm85zhqLtEYp9LYp1kRga8gVwqp5fyjRcyunrIyWDQAgZS48Iw4K4CQmn/x+JyW82qDqQKs
BsyoePFz+iBdbO9jNUMh80UCE5ij4E7veW+4+SXzAzccU2CQo+IvWL/IBVWl0+0CwiTUzt0jCzuT
905hOrWP+/lB03YfY1bmDFViLDKVZw85cRBq/dazouCygIv2RoZrldKm2dyUd8ycM4dfolqe12cj
3XGTm/cSsJd6UGKyAKbvv0mCvgT8pkxins9HHKgvTm873wxXdWTnHqXqzkzgX03bBGMUxixQZSrv
JQ5SZP75flnte//aD+QH1H/BFeJMsgQg83wHTsZ3R+5lDot8tDQRr0Mxt92gyS5/YkWLbrhoy99O
BT2oeqsO0vSdZ3vDt8alt6o1N/tQzKHKAj+RAE/jVUuaWWu98NmXnrr8vOPpN7cNEr5qdERJm/6B
lkLJhV49vagdRrd5885Wo3LiIFv/uJUrWwTTziURR1HGi4WSE6FLGryUnVyF/gdhVzcwC91M0JYv
WMeGWonfQglbToc5pCsQCLZUuIY6cnSc0Ab+yqhLjvyHqVkE26JwOV3z5b4qdBeQ8GV2P1Wf4DCP
GRcY2JC10He9g9bL7e2ld1fsj97m0CXPlkCtyjaKikIiqUNxY84XHJ6pRGQyVJFrv/mFw/+BnYGn
rHTNI1xWPpKSZZKZ8NzIFfMRv92htAFzpF5g1DOSQMY06XP45P17juohO1ajE6cWONBOTgW2i4h+
ExEY8Nb0Y5RCHHEuxsXrjztjJ3CcpHY8WgtPR7IQ907vqGw0gKjDVOP25mh9foVLMg2B9NZyfCag
6P1Xf1CN2+bJsDUtBgqf0saW7tXPJGtwCzIfQMUgU+X+w+v0A4Ud5i+6sNJu4rdTfXykVmt4UZao
dTznHsqCJdDj5saGLCJLnXbzEyD09eEU0wKA5eUra6OteOTsUq+hOosOdY0sTCXvSfFQQeGHAcCT
Br8ngHalPxm66DL4diflOP+aBy1Z9VlpOtH2rqLjvWL+dnkDxzXP5fFQsx62XW8QVC7g7sXAegAy
5Q2aOp8wf8S/9byPe/sF/6mDSqfZgbLgP9iMMi0GTkMzpxruD10QS1/bgzIkh6mcZOYRFaWLAVV1
FodNaGb+BPgRSXzP/da4EiZsSxWqtr7XnxCmS+7LO+00Bt5yaZf8IR33mtv6lPjPV3LTmsnz0i8s
te5nyfePlL99A2AajyZWKI6ECHexHLzRkVLRsuPJUpzW2YV8WXfmqSnz3l3iyVfYS5HB1zQISruI
6KpTnL/gPuI/449voM5dC+VL0RaOPaHp/QMiTh86dD2/U5o7NP8Bm0jPmNW5FAJ8K0drHlnyivmj
m5MeI0LLAiZWhoKHLDb1M40EK5ba9KOUZRE7s3XRUsjJjegUrt2ksIrQO0xs2KyNiPaR9zheyDlQ
TufPjmPBn4Oddo6O5ecpblJIDDsnLMwT1Oz8Wxm4xvLRehym+nHWNq2qVWoTSTmkXpF+m7B9E3oM
wAitGTSYbCd/3AtPu+OJWanhWzxGkbdbTFuJOy4uAG43mLZHvQKGOfF0knC62355r7olGwuw7iup
3UrMdUyzm2H2PzS2mYx9v6HzmoKBAbSF9BIWDcdoBiMHfOqak6afzBrtT+YFX2JWLw5TcogfQKl8
YLq9j2RkYsroSvPD2lWF8D9E6WVnx1P+LZMnl2yUxzASWUkpWChkVX0HOFUC5XdjKSs8yi3GVoFn
5mpyV4xrSUJrjjIAgU2ajgkedQQdcRR5C+pmj9cUjJAcGoZU5L9YHDUcPUXKtqYfukScNCnUK+yi
6X+wcZbCtM+nGtSLBWGSPQlVUX+K3NAE63PVY8EBhAXo4qyUk3+7Y/8SpPLGIR/AjNpnN1+EnONo
2uwU3mK6gwxhQSY7+GpOm1DRscezzvgxRY6wTPx7FK1hpVENbXo6JBBcKxb8M82GUq1g5L9CDu27
o5t3jHkNT58laz1ZX2DTjgLNtxMxiVhztRrwWRT+4kB0lkpuTrOFZ0VVGsC9/zx/Yw7yFv4R2ufl
CoS5FnPIdCgWJEFEKa17zH5Q6GnAQ++ttmc0FsUN6yfSXJJZs+wZErbKCzNzD/Tn2FNZTSEXaYo5
s/3gyiaNjOis0p5anAIKLaNAW5LPxJz7MC0TDp4WwCc1MBxEcpaaf28xUT+cLs8chPTruBMbdQWR
2JhAwHL3J5niqx+bWy8z5C5LM95qs6onhxEbyY3o6FENiCLWaDc5YoKMDSwdBAnvn/Jv/JuByMLU
SxT/9vEYHj41hohAWaOS2RwgDjtZc5ifySJpblU+tNUlp1CD86QUYH8qdkRTTc14slicPw/MRfHD
nII3u78tEvSeDGyS49GPzOVgnoUtz2mjAPJEn4HpV8fXbrAQDiJ9wu0CbHA3MzlQ8Q5akl1yFSt0
wx4ShEVBQdXGmd5f8rhr4XO8RfRyVWshSGdgl+3/NoIdh+5Q/d5nMircJQp6P5G4gxDM2nh6/qLo
VKBwivbNDtMQrh8EIHuxIEXZZonj+HB2A2iCYU9NGAQTCRczvYhjVqrAo6OmYC7BiS9L5RBTGoDq
S70AfgP24S2gZchtMLp/pWEmEsdgl0DYm5+upFyOZIWRTZC4cLTWbl5p8I5wlk8d7pUmadUy0HAv
oQnOK4c/qrPqrC9373M5STPr0PKog7VnulpUNbJMdsLj5Ff5ptfURqy9+zGaVW76/N/iusVek1/q
04LKUg4B1uMVlYRpIufSCwjQ7dURfzldaL7NBGoed87XYW0iBo4jZ7RTJrrhpo5odyvxZJ1415jO
Cr7FU30ExWKs0Gh8+fMJkXDY+rftX+BFhVgC/gTTB2Q1rvekVgCYkVYBmln+oidP4keYUozLpW8+
498LL1axUyNRBMNj5WgjswhPcjL5KXpzOsIS8W1IvilUT4vbek+nPGAZlv57ObKZ1Z6OAZFbUYw9
codGzxRfmkL1ttoP8qxbx09ajb+CRKCh+EAi+PQIUjqZzIfZwo7zX3s9Pl5HUR5J8mcUxE8PtyG2
/EqHvaMkfEbuc2ZQW2UfZGPp9WvdUpxfzoWZm81nff54FqiFcktTJ1c1kkNY4JbHrdy/2uUGxykP
yzBOuMFl6jgZOU1aZm3vpdMwtrVQhA7pn0or+fTtjk2GnsWxcwbjXMMPe4l+gEecE4AU6Er7e2vT
cJZv34+JPctKb6YISDmgwvhLz0ndnluilVgSqNhnfgNXqgbRQNcVbqwssWmfI1zTt0LqNvpiG5LB
oCYzRWsqc+xSDgqqT6+Ph1lgMPSLTxGnmciVNoQCZKdf6PsyY8Vo11D8tyrWBHeudQ5FyE1Hu1Mt
lbpzonL83trzXyJR4IqLFBS5BKTOnG5zoFAGOmiYedl4DtKmk0XqncXMbmFKdi5YFgrs51fs+NX+
VMq/mUglyKFp4ImbcW/xZuBTTUWUcMgnycJ6CO4y044B6FGta6cCFhTheHFT7JDk4gN8BdwZb5Q2
PHsEwI/LvP+z4ub3mKXGRRXEvaZTTLmoceSnRpWedvvsWGD7ycFrxRb2IzG3TrO+QdaTTTkXd6Nf
GOeHxn31X9dFgDyNnVKUVLtptNvQX3cowB0755hcQtQJqsUWDpFyU5dCBX7ODqRpOZY36NzmT23B
eR4T3tnH8DVblwUb9T1XLoUHRfnnJhuFxXN1l0Ank6sMKERXHg7cA1/vmsUxvdPftcr24elDNIUy
Cv9lSv8QofxWBdhT46Qbdm0G89xno/MX6jDpsFhoQvrUjS+jwi/SEMERUdBFAlHPG1Hvb91IemnN
mGNWc0rglklT7v92fAsjZqUBJGa7Er2YfRJgCWgpOqIsdLCXUl/23GJ7S+9Q2C8/Uld8BUWcq8rb
cC6HHduUw2Zkfg1eosPAmJUi72W+3REXXn5tmkl5qNM6t5xNld4QSqeYMaHp5X7N8YnE3SvU3gdW
9n4EkOUMJw6f6qxG1XNVILNPC93ojKGUO4PNIdfpiJb0Svi0GUZLonasED+PSKWXTzmSzOaYXqLE
hyrLqSig2q8csh1apOunzOL5pclsh5KiQ0tcbHPtG2Pw6QNiqRg9ILhhYrJ/4wMyYdd9tXPOeMcn
qnyo/RP+zi/AAmBi3xvR/jfHvXBwLYpnbQRFOGFMbqywgvOJHCE4MC9JU4K4ZbSYoC+Ivz8wmVEp
AaXtrUDrVlVGJLzCecT9Pu0+VYEkqZPW8y81QkMu1gT0e8KGHDlBT6nc/sxTv3QuZcRPN1iIk8M1
d2PFhf0fTVBDlkhKUISJvoUeHVqXAeSgVxXIe4H0VhUzMVkbFQhclRWbxTsuEdzS8P0gmfLbhVBE
TLL+vkqPVJT9nE27Mv6HRTjZxHQpD7V3ax4J0ZcPugtVmkOZJGQK+m6HuSKs+HUcKeQsrUvu0ZRi
hJRgvThVa5fWdBPGWrjFa1/aYvm14YYV9D2qSql6Kl4w5bm+eIHWO5UERGyxMYVLp0GMS6cO73c3
pG7iV86s/MVeNlxE/PtZFPNzTxQYeexBlAcXnvxAQgECB2xpqVn+/rw3w8b+2olJjv6Eo4Wr5zJQ
bfWNgHSXLmEJqvv0FmF/TF1iC9R7ayLXvoTc5a4vhF2t1CpTzoIwwar1XBjF116TCQ/7LoRnzSft
l6iMjRSCX7kz+Lu+XLNKYVQg1Wx+N/u59yA1L1pDqbuAqdNnY3bosGf1E8faB4Z8qqVa+A9p2ubm
T8OLpRlmiug82sqMhMnRK1XnNr8gEoviaCt8jK5E1cNAuzCdGvRb0mKvU79uqEO555Kt+FbjKzoE
hawmhBxIV4ZmpO23QvKvcFSXsVNLyfYvTFy3xeubX1ammLWhT8MQqw5pweNmLjbkjd/cK6z/YLLP
nEJ/h35IEkbGiEi5cLDfX5EcW/Xg8yCUTAyJXJ11jC7W97C/rWLB2Sq3OeVQXO9GgZ9zZd6ULWOW
UzKTsuTVlv47xzky3clcKZ/2fV+Pvu6mGnSwL0ZOQ0Ho2a9EeOZ2J39dCeTKsMnTmVVotP6LDeeH
UpM6584sXhthF2HMYXco5EKZveLl0tLwXVDgSFNu0nHRA/NSgMKbLhHLfMURPTDixRBLP/UrenPb
QPgXfK9GnntdTxpAgztq5d8eb6nR4exuzM2MDTUWOvWhwFbnIYVnymw4BhbHWl4yGkmajSOWAy4N
myBpxFsaw+2+5BkDIVsXjHaAC6qAIgM1hC39f8I7GxJYxLVREX8lyE16ilztdLmeNBa+chnpCaBP
Dwaynu8LbR2LXayTu+RwnMeQFV7C3/JXrs1pQ/lg5+Tp1ULWMUaKQ3fF1nKU3BEl0IqganHCD0BI
U3wvfM/aVQrAUgjM8MLB2NyaTIJFIxxRgc+XMBoozEiizPHh5A3XQ0kiRpfbTGAMY5TtsdtqQlJm
kAZtltdBE/HjStwSY4ZOszOvPFpFEd3+9UWdsk8lblhND9jEFbqBVy0dbimf6X7aAeIOwT1cWFeY
GJ45dNvE9Kn6TWzILIAc67Hq4Mm8E/J6NEKZKElY3LZYKnW+0J86bQo1j9b+15BM4161f18HZjbS
an3GSdOwNzQYZAbtsE773GymSEdj1gaYLstAL1+l9u/n5IQUNrPVX4feuZ+RqkiSRgb6+B0s7jTh
Z34lUdsufZr18pMIQWEZ+olLUbBezNgikp85/c37xhB1bC4rZRTTKfNRBLlqDTyGMI4ObkmhlQ93
Z7VCdpLAooDQimnOk3sQ7mAo6f0wa7r/xPJ3ou+YfZ9GU3ripFaNXNqR38FtahtqGJSNFpJSphTk
VBvrhUYwKcjjdij1wyOOQ+rpjm7y4y/ga0WpkvHs9ksDDEVijf5595baju7LALyYAjrXT3BNoTxy
43cYNCs7NpAJf+h6Whh7fA2rbhpbVhn7UmE4es4irvHOF1BG+j4QbWaLi677H77JMllh4xeAC5Kv
da0C2K34mFCwm/SsPow32UyjLUN0U5pt7irTTQLVhED7zQfdCRNhJRON5B3k428f6pNQyVRH8Vlm
BrXrG8TrfNh2eIs0ZQdoTZkysv6A1B15S/AU9hnxvOrOghWRed3b991ixEv8S+Xmac58u1kOxZKl
RSvJd5kh5lzNTKrCqjoVFTaW8n52iyuPlorf/DuYAuIAUEJUMsoeJTNqcQfzFv3Ucj1p9IhnnrGt
TH25bThQwder79iVGI6gn6XV0R8bWexu9wtrZO/zmXQWMPz2wmPjFLZP6I8OA5qau9lMtgIRMfIQ
n0C0anrP+78rzVMjb6BUNxGQ66eyFrbfdHe7URIOHoCil/nR3ZRfL6IYdDT6TylSnHozgNX0IMWU
MUUisbNb8iZbpp2dYU5ju3WJ0E65v5OAUX5owj88eGX0npS7D6wmvE28XsEtTrRZQ6qUtJaWgkAD
FcDQD7sfVq3OhjWAYqdLvKtLdLXvbRoKPlkX1Evg7aP3lIyhbh3+bXLO1ZusmSDd1fjcjityEgHm
K7g9NJ3SnYEI3mIl/lKYPQTaMMDEbTh/Kg4YcDa4UVlMBXI6t6l07m5CIdaTIUZkv3aTL+9kBbqn
lyVui1cOQK7EjdZ3H9BKVs0Ds+1KxfDx72ImwcFY9EjIIAnbfDlGjcbH7KeqI6/Vl9X6wffLPLAc
sDryN4FExRZBk1KTlg3L/kJZ8BnnymW9fmBRG85oghsdU4JD/aIKTJSxOEQFweGtOHE91ifY75bh
LhwdGmRtFqF4JJDK8MbYYxrE1OHV1GKv6QU5gUbWUZhi99pWf6wX9Vo7GBU6ZDZZFlOcrJO4mVDo
rBw1SkCRKulpZ67vadXLUIMuX8r+gZ/LLKkRwjO0z6CqdFxXkZgtmm7Hyu4JwnFbp6DRm3aSTOjy
qINEFR/5smWbSyOqltJzar/0iLzKLWQXb3BabfFrKjcklxUvP4beJRX2Q+e+Rnnc86b4soRRgw4K
cy/4k83y9nTp7UuvIXVONvwabfef8zHg1Fj4yi1tWgMQm1JRzqYumK/Eu3fxZIqDeda7cfAFKADk
AKvfibNG1lQ5QsACLBbR67WsPzxCql/JlqdaEfC340GJ6G1Vzjd2y6yrbDiVHOSw7LQ2NlfzgIYw
GygLJTRP0e1bK1F3YCVv+qe/4PfJGKPPFPlS9D1VvON6zuX9Or7JgRWb46ON8E52Clpj6jEHyf1s
MlOJh2saLaUEKcCm1itNwJQRChxbFlDy7eI0W1lp2K7HRux52q6fmPFTtAGafrLUu7CpYCs8abfY
9R814nplvmHt7RvuoF+wmFLj0U7CcdCly2AYKlH4OYkF+JftljDKSWeq6m9JhW0g38LhLBGskCrI
poDLdxsI79mKxWP7m7Mw/xety2rAbRyOaJ0+VJuHwmknRCLjMNJyJ2novKNO6XskccKESoMaQH0K
fsyKqoMyP2LWyTB4bGxZe3Mt45UZUZuQQyXl1k6VgFlhTKLx4Ny0puxGiY30gJDFkXY0hvqgvPyu
PgyHqZb9QkHrvR4zjH+WAA86TeS1k9cpz4lBr/PSxakgWnXp5FUO6sVQeUNr6cs1AdLP2wJdw4CW
X/qmOAAQ+/TTpvr4TLhDP44IlP6ZX01wIVrbMMyeLubvOYieQI+3bcfVklLpJ6u1fWCTAmuXdOFL
v6Qo05fcTpAxb3jXiK9GRYEQ0Zr20VQkwdcAsmtoDHnkX4PNXDw5XX7Conl4vLUzvoX4Y0bN2+M/
Tmabqz1wyVWbtqBx8HsClfjEHNpx17kj5Nv4pTbcPqbCKd7uBX0cNrk2qeJ9iLaTF0gO0Wf++ist
KxVGkUreFprIh1cjAPSRGHSGqv9LkxhRolKJrWcAlcy8rUYfpQUIl7+6n6Mh7g9j8eHkKyoB8weZ
E4FxRMLOwIGrItS5OLosAySBXdiKbBDPQK1iETuvnSVw8EWDc7jUD4KE82bQxCqdLUBON7kr0bhh
00J1PNIrwPFcIl5T60g+TIv4Nhtj2Dcbctmf+ktVP1DBBv42CI5xn3atoNTAYN0K5CFKIVwYR54r
T/+rooHdTAMUHY6u+sAv+IF0+vHnw7oyvXFWSY94ZiKr870UpJXgV9kADQerUkKLoMwWIHt1bXvR
Kxv1kdgHowdCuBtFpnlIZ9mG79XQJKxsTJqccEigF1NrEdb0TlhaRWcKOMqBnL4BZF71O4UH6w/G
TlESchcC8opKiggtONuEtrVm9AmGylN0dpmh1tRkadJ7CVwycW4h7veyOiH8oifb0Lpz5txyr3/6
LWSpg7tJmEi0xEVZ/lF9FEJPaLEWJZcrss0L7d9q2gaIA5sJuHfaLyeDFO46rVF9d+hadwncb0uV
HC9EU06A71TtJQCl0IDV8ymPuvDJKuWDRmssPx/avZBhl3XRNEVL3dEuWjcJR9ssgB+nKAFlUN9/
qH7CoI2RvFCCSrDhAlaunMJzJwfTLy/gV2nMW1wBceZzZsQQnMV0q/vTkRPf5Ng00iUql2qGpynI
ZP7W1+vHGoY8YiTdgxxdcYrl0kkZOqO0TUds4hZeSYJiH5ABRMX10aGRp/Uyj+q64CMCV9lUB4yk
mPHDBoeThNM0R/VCmY518sWJrfI3DWGDwXDYwUPMbp6SUtGEQG/ukVhiQ8J/jnwbINfX0dNqE42s
O2VRN18Gt+dH9OKHwueZKWW0dueYmXtF8iJZG0b5Uyc0sZLB+t85UBWSDWothINt90swmZwRC3jF
Wcs+vzacidt3SeRfYYeJ6wEHhG3Y2/tKgemFsWI/DzkkLHKY49YcjzZpL/Oa1tyEsjpxm9ogkk5P
CUGOMq0//UST0TFeUj/2cRsBx1fsn7fO3lDjjrSh78FAePmxG6GVGpn6GwwTNVfZeXAETl8o0iVZ
GWCUqSk5whsgbSBTTCAOaWToCD3nE+viJkdQ4pcsVt4hSC1YMVe8sVf8XKVdvAnyYs2730BADYjG
V6NwHdI7+dqAN2szy3giTU8wXs7eSpJ66WQqXrAnyxyG63Sbz7NuxiwTISyG0/a2lj8lhQFGGbY3
LoEeegPw3iDpLSXjk0rAehTQ/m7BtFcnYGz/bb183DzzIT+uFzoW2/Q6kNnytIS2w92k66VDEug5
ENihVpxu8vhhoa4Be5+fzRIEATy2ZUtVwSkyowf3LieUQfaIEt8uToU5rsWu+/NjdQrS0Jaj8kv6
fqQ/HN4YQFkNDlnCPf7DNhzuE4+KEZdVMywkvUeda+z3kabPCB6kSqhrQVvHqHWEUhxGyH8LaWEq
czD/Px45bfuCppeidwzn7uBlhkzPL57saXyfWN7E6MJOxaQZB1rtJhoQApvpyY9ICBL4HhCOxJsk
cPq0BMgjHRv+1Jw07EukfQ5Ll9YR3dsPl8jaipXy5swgzVXGeBk82HzJuBOy6zj7fxISb2j0Pf9E
bPtYjPOChDxUjafQ/DKeTk7NcFZ3n9RuAVFp78v15O2XreLMDhTngN30q9uk6e6HDxkIiS2QrXPe
4kXhN8GIile+QxqbrWvaW1k7uKK18Cxo7SMJUpDYLsm2DUMWGFXX3NRDj9dgVDwye2C63el00+q1
Mh0X2zFBwid58xEpJ+aKAct6GmpPBQoLNZVChE4rb7jO+GOq1e7xUCg5rnWLqOmiri6yf8sYJIZP
p9rF5IOJ6zGpKTp1VgrqKevamCd57iUJY6qwc3nRYhncDjvR9cKRzaxpbW1ZTFBAGAuisyrJ5IDI
xvztyqs0ErioRYi4/BPDX4gTcqBSETNT6OU0bCuMbIO15VOyHPmZBUsSQj/2bZD6WfBaoVHeJgSK
eCghRiMqs4XO+TIM9I6xIjy/ric1vLhcyDjmYWWNTKMGBT0CQZKoDL5QSjHxASDqBUv1NAl/XSIY
Y1XIkrXsYwvvB9YLuOB0FXJwCpoHduZiR3OAAOigobAdAVn5VjE3bxUhys6tzHtL8ca07z/uDCte
hTEmzksQYwYmnRwkuBZ/PvBog5fiS/9LiLaUM1C1Jo9AkBqvpxmyw0pxlOfAhUS231tnJpT20Wrq
kw3vlqJ+k2pJMo+rQz5UdHqHruBs2gG+pvwPreY+Qop7YllLUK0g+R3ZOTExhGtmxqVOfBJHFEJr
RLLZHUwK6ahMCq6v0NMwS/FhpU+NqaPOL69V0i1qOxB+Z7wZywJapiws7Xl8wTf2g7ibzZ37Ey8L
sFeXXt5ZctL5bT5ZCSj5i0JjEpOJ5JFyCZdgmkI6qb4D1Plp1FS50jc4litfVuuOeIqap1jXVFhs
sB3b05/QzpACCHjF5cMa/lf+F+CliGuQcI63/AXVom9vThdh3aya2HkPPX+O/yLLC7gNGVzUeojg
r8YbwH8mEko1ZpY8KZQCmDMjmd/uICEFZh7jjjtJ3d0GFFWapwGl2m8m+Z+B4cGsmxDw8JIrfyGA
e/DMZDHnW5Wb9F6dXzi9TtsjdTjbVTWyNmr5fcOvwcwkz8l+QeAhu72slB5cEzqf99MD3cqvREU3
6DNiDD53ph7BW869dHcwp9iC9ufZTbd0PnwHw4JTuQ2/M65S/VV1Rbt42Spkt8FjtOHb2nShP3wp
tb/DjFguJENeiBvTZifS42zOvh+MMBKCUN3zOtDB4RUbdiXb5zh2LUh3T3nIzBMURlrlHdzY4vG7
S8fJ9kojR0NYfoUowCFkYnrH/g3PDE7tWWqigbkZ9LPcdrMG5THDO8J9Pn65BIwFYKrJw3/N81BT
FVqwkjDpTPQrlKndkyN+5H7Qa7jvt95ABFVY2MaeKrC1k3tBIZMP4yZwusGQ8zTS3LhVh2szTDUv
hnfaVLI4jI5Pl+JA4jEKfY7mOKz9yT7YVde+nSBGUBetVShqUsDut3p7xsZHzVEM/15mTeRcPJfb
ez72Qe+2ErJMCRdfdOtZyIeiXp60LfittV7aSZgKjaZ3C+FhN8dohAFoQkukeWkhv39XIdPijBRx
m8psBH1U3S+UEHa0dseVlyzsarAMbc/OGzl3gMXmfD9MHF+/R8LK6Oiyn2RBk2Ar0E0wgzUbnUpo
KzVe41m7Xr0HFYPDwodoCmshHgTSNdNzjbsOLXeeOXIvJTm4hrzIGpYLy6UN+RLzHmVZIFhhUuA+
zglgVgYli1Sf0lLVq+voo5TmRmFY9wqaaXMvMRpx8oxkKUYpl5A6HZxHHi+4mdxh+fsyZQ+IhMe0
V+V2FawsuRspaG7ZtnF9zRy6r4nOMxZG+QX39W0JNV62eKSy4aF1zVIaX7JkfpHqhienJLbyMsdw
RQUIFmh6UMOI/RFTaKIiDfW5QpEjH9B2oDrl0JLWZ2ixauFKyFKHBk+efqNhgRWrMbwQoKx2qmZ7
t+LpPB0ySATqWj9Ocyudozk50rEyZnW2ioHInS8sHokx0gVDgWe7E1jiRQse1XEocNNB4ahHFWNb
GTvWmPNTxjN1UdmfnA9NUs3yxKDv86ZeXj5bpRE0GKdnwXTYGXQCDhoRvpBlthoGilIpXjnQQD/K
yGzstPO1GgATevTsMybvMWJZXfmlWaTVyKtHgllhY52/tyIHTNAmt+GNqRK4ekdZuSwULzh9ZyYF
SfETvuPVnQmBL4CvaC61VtDBIcXIvJam6f8bFtEeZbi/h/xPByO7RaqFZPdQKSGPk6nFMvF/rQDI
4lPuoGaX8aewX6LFsaKjaCbGuBflaEyYsmwCIztOdQOxrgbYPwRKzIp9dZ1K6EvQRgfoQWigtQPv
GHT5fOtrj965QC57RX8iZ41o48ePiVuiKmDezRUIqKqcxLK0So3yVoPU07ef3MyjrrrObbzePp9r
UsR35F894E2KsNgnz81ExIsn07/ps15Gcge99is+hU6ODvWpJDWruZpasEt2U0Lu9m4ko2TSiXwZ
nLDo5EAAJAC5cNBCXl40YZs98ZZuAtiegVkyLdsWVAs8dF/AfMOiEkCFZjJMsPXclfLgR4QcqGeV
JJWfKLvQPaqM7lITe39jS//d66X+Fh1fXFj3IsFwRlGWQ5M9fy1fz8zfrjI8tApOEOPs/y7Egaqw
nDWzpPPufeEUdlhmAt7qxgcdERANxfShjxk79UD0PUbswACk2pMOpV5N3usDhcwW1rck+UFd1uYZ
utvVE0Yp6w5O40q/U175aRpnV3jPRa549hzfqpaZWSpbQiYDAsZWCgtnMrMMMjBB18GzzCNqYAGr
UTMlr0v7cr74ms7+F73mGlPI8qOMkLHzoyovshWu8xcujrdKJSMVO+dlq3mYa14/ozdmgY2Q6qrQ
u7I4umqh9fyJdffMpeDOd1S8mAx0IwxHc2qzGxvIVliTSll5P4Yg7hHuR6bu8kS55cNLMqSAjinB
XrzYelRJt9Lthos6FnLZgD3nhWnb7ScYQ7+fDEdc5fdB6fTI2tpDMYtJOWU/5BGqSG0nQo3npVT0
cAa65+13gQ3cLHzE30bGUcS771W3eYUsXYiuleKxf8B81MPst0CCHCmwuj6FRS1/kmNBgY23wS0o
aoUNSr4oGZDOW0q0NNZwuOdrkwV/v9i3itb3BV4hNcXKs3+qpNHz2yaVEd2QVljCC+5Rs7HRwgVG
KaAPk5upKeGn8AL9kHXZtJYuRj4ZTGyfqDpJL/iht+jrWC+XmZWYvnJpji+qWlUkl/kX+qSYcDv7
n+haOdjAyaDIzUNHbus/92may7c6e2PBj/HmV/vuiYWWjB5qr1LGKBxDeE2/Lzuh6JtykZkyaExe
d65Ut2JB4SXP7DVs6Q+lM+nFcdp+DYe/k1zRW/8LPR2pVUrjQA2MtJA5gadOkqT+7/3/4XatNPWr
Hpx+dnslyBDU50mnJUu7EXL4/JLS6if21fnDTQvQAxfaVYT+8Le6y2Jve+6dV0Dct6L0ZjlzZp1j
8wcF42BgP28IyQraFy6WjuKc4pFIuh8Ol/Utwn2kDU1DrDNyrgQuWTYQcJYZn3s8s8eTXQpIBm2o
hyGsLWqDgcuUY09AmvdHO/VByb0Li8eI7Tg34h39+RIKORUS2BEC6iGvBKjLLNwiMl1/m8zdPNP9
XwCAHw4TFntltlq4gh4Hl/b1F5uLyTK97b/M+GLLGHlWhKwcNLOOAcgx2D8p8llnz0SVefGcKWMM
VjzaWpaBJi7QGbgrZ1MlVx4HGY09JFsF+W1CthxvG1s/DR+wPhG7KT3KHiMZZRJL9OtIaqPi8LZ7
P0U0Ovn2idCEsw99QgVigNG9881ls3NrmiRxH1v2mdlbyt2v5RxorquK/o0RmXnPegzhspwFVIXG
uHnOL0OkfX++u4B7zZZ2tiwlN9Ky+gHzBwYXN94O4rTz5qSIv2/v3XNjan7SVsKXgyDu/63hbuts
d6OhW4268NbBfB91EmjIU8If51U/ToJFroo8izub8QQolYRXxTWe3bUN0s6B7pcSP1FCPfZj/8Nq
CWKdcXcIaPxBVCFSPZ5drScSWdkTsHmBzNkqY7X34WrZZg5kusPHTU52jjWlhH6aeya+cmveHUeK
ayElpkHN+ZFNe8+rldcxc++KRqHW1SJfr9W5lDIFO0qNQ4SQbUPV3Izg9UExiUeLCpgoB6ci0+qL
O6p/lAwjrUtM9GmDfWw0X72PSl1qkZw6AQxd/WfzkDOO1MwyjHZ6eLyXMH6onL7K7fkDMG5JyjVh
SfsBgkh+umL9kD2fJT0lgLgSHr3vaokAL7q35oV3YkZ9ILh07v9sK1yA987k+JaHgUgRg72dE/fA
oNS3rYKYWxHQx11821GOgxyxCk6eZbG/XL6ZuHQIADu1eaDUzWvKTKSHWuR43GKT0xDsS3lKFyyO
aqPvFrnpFGJhmU1QNvOUvGJgi6PjUgF+ZIZVi9O84f2aOItdG+0TgP5abOV/xBn8tTPUxfAuLKx1
eM6buj1W+3lvIeWGgidKCRrNbZfjtk1hyh+5BVbwk3yLC88k+7+smc7y3FuiC/qowj3SX4W1NgZ2
PcDewxKaKuy57rUoSJNomVcJKd3bfOiCGZchbU+oeMUosIx4qax5kYeu3sWGSrGZ3ZQ8EmAMyrc3
vxBZ6591mwu3xewZ117TFXYaLykdi2T0NrVw9qek6+WGxrRbznpSZsV3QC8kGyZ4DLjpfmrfJ9mp
UcVWgwA+giKN/Xkx7+0Dyk3zSAEmu+vprvCCgTYJtrzxd/vQn1OKuYVHCfU42yqRqT7YNo+l1a0X
jgQBFLF4TxhCFsXkCIoJlGwWNybYroUSCG81spUSB51pn+RCu1bF3LtNoSYxeMNbghXve9QPUxbc
ZktHJVghGGSmVZjJMIXZLoxZSAror7c/EpPdZNbOwWjTcug5K2a6J31jLzw3SbohnJF3LX2Z/DKC
WIJTSHyZCaYsahd8BLz8qBYjdV0p8cpBMvdLzqFl/9d1MKcSrkkokfHJvNEiRnhKjXRbpCUaGGOt
tAKail3w1wHpSrYCC7yGemFuI6mSjk6TXrd1AeCLOEk7eV7RoLrFPapzi/ivBL86UfWyfiC8HgPe
4rRVbuRXlVfhvhgaD+6BcMVsMPjxFJF9OHmI/irYGxyMmlvsOYQNPX7Cmfe7gKCnQmQdswJQghGo
4dJjKmMbi4MlZmEyfQuXkkk0dgTgAMcCe1zVt7WNTR4XvvHsrQSI0+7eFdjjk1J7SOm4KX39mICE
KPzwsXpy2rurkLfcO8Emtqn9U686TevfJ4i4hX08iKZfW3BZ+4wdflJ6kbCqjdCVjwZvPHRe4CUP
KZ+f/WA9PauL9JHAMOR6O8bIHg62Fu+qd9UnPtou2e0Ya+dtzFngrU9G0GIMj975IW0v37X7jfT0
GdSADo7Y9DhtEK6F2BpFu11LdfumZacFk87Rk1k4uM75gyV6Dj070dktcFzkyYWBg/NjsGbWU52i
fYUKasftt5Md239Vr+eG+IVbl2FeKzaNaZwo571Rxe4thnpSf32IqaJgqGvkCHnYCXg4F6QLkwtI
uy8wLJRxNti/sDSfMeu+FgQuezIaH8WNnj3ZJMBWQGBqvxEtSqGE49g6dAEcjcYNStQZUkSGFA7h
mGkNyi9dqDK4kBYhdJp9sTVriN1VkCBL7TKo90KbXHyc0USVMRyPjMVo/e+zSX3LlCr6QdfH0YCL
PVol/g4hdxvtYBMxgoiYTOfLn5g+zbjWdvBjVTn/EeIhPQLPoISj1qdfyhzHuvptWAFJ3GcV8xJq
+iXq2xvPTd+q9HLjfraddESYzIDw4RVAYctUb5T9dGF44Lz6rMQcCMX+IkP7DL6ad8kA8d0+vn/v
n/03atnAEYKy4bRZ3RIRFv2UlQOZPzifEIUO4SxPYjIukxKOR9roJybbdmFv4VejNdNO9kZHJw2u
I/UV1k7F69f3QjK8cf066oNRqbbmFmMcZKadCeBLmgsJxr09Fv1Z8VxAL68gf5Sdou5ZLZimmLww
koQY6XJr0jnl1GK2zUSoIrINSICOm2kqEik+2PAaK0/O0Xq/tZ/DZTW5xS6s5+t9ZDRUJauE0vWa
adcqv/h/0EFDj4YhokGCWMfoIAB6ZIzW1d+SEgOMUNqP6rgLe01GQ8FAPf1e7Mt8ruRsA80H0wPP
UGBk1aWkdOjOCPbQy/xd4j0m24PRHENydhMhVE1D2CDU+wWQm5pqG5oV3MwKdCzgpkJksHdS52yr
vBWT6OjZQzwSi5VuyP5FUYDiCFLC47zUVONb1OPX1nW0+N8ecxFU6tKseywcF4weUCn2Tx9eSVx5
XorIbp7TZ3m0BSWDMDpoB+ZnWguYlxv17X8u5SbXSS+eMSSksz//BVDz38jhzvW1x5ULxjMHA5A6
OUkuc7iMVFlmHfyy8CoWfrrZKeWCLLjmIX0vpAabp7kXgA0/BDIsiN3AFvtSWIbnndYuCAzHJgR6
dqF1cIyVDxXi6aH0XlzHBz8hY2ROPv5NNEqDZnjMxrCt9ZI1kPDQDdHr0e+DAolyqHyiv+MMWnX7
08243xZl7F8JFhpil80Dzg5rvEzDhrjHfVm+5YEFF2qf56sYSvfRZik85RAG4HlSzczwALBaGvIF
ETgEbNJ1a2NhtEx1OIqYdX0CMP5QEbb5QtyOOFcJx87PO7j5xoKyYiGh9l5dW4qoksXFIWUTPJV1
Z1dbAIzAPD0C1LdBNOWl21eNBfijm7NuIB5bYj+gArIKy5KAlo3WoH4gxXuRssWXAfYbWMqwHkus
d15osxO6F+Yf25pMEmM1u+QOtGHNz4q8eBEjzMkIlprjWUQMKghOeHuoT0GuLW3nldU0xOGlxhXY
uphrRFBs927an3DkHgbb7BOwySWXgXGteTWz48r5+2nBIL3ms3QekCKo01Y5XI19aXHOmLzDPnyM
uujKMluABPA3r93fwJ9RNvvuJVnP4oHHLnv1ra61WhQxl107ntyqBulCU3kFIE+sM70X9fi27GQL
Wd7QbB00tJJCqVao6HAmUjIRCNyM8n3XYv3ayEY50rIA/+oXxmYDVNQiDjRxICX10ii7WsTpkjdy
BUYe7XC1mk5lbB2P9o8pzAxSiyIjhBnkOg6y9roQLjkGVAYcEea1tagp89xo2cu7VDqz1fE2iisr
41Ihga1b0CVaQyk3CUmyu51j4vs9cbatPru8ltMzpvNXAB1egPEqYUQXKNpnIO4jBPqdWG7SVh6G
NQ+/OLbGIxrkDNRaiqzihaIoWEzKiTiVag77OMc0mgev9EaxptjRqL+Ckj+YiawUEHCThd0SppVl
4dzi12EOqss8PA34jYsyepZ1hzWm4ic9RulszOsSmyHYmBBQ6gSD8g8Jb8Spd9a+NmHzbYVXC7Ku
x5+A+A3S75HgTKX07Bi8DCmY6Hksia5orABKiXalZVfWGQ0IEsL213zgYLAjwYiGv2OY2U9JNsQM
2lw0bnl/tQPQoFgVH9tUb53JtsDj/PrsoIV6tCCurOfTv8lqrUYGALfxny382TmOcdaLEODME3e3
os+FBIhdjw0xAbQ8IjKRM/zDEv4QpEouIcdeCgtJJKgvoOZAQw3e7LdVTlGHVveuDWPMimOFk6Dd
07tdzds0urcC98FrhBuHZza7xxdSAfgMS3v86j5MxnuSXfu3CQfrPXxbmP8uVfcu90HPq9+V7lc1
FJSH9SCZlyVNSxDshCNbTkzSlm8v6Xr1wFvJEZVynZR1aU5OIybO5GOZBreZGdn2dgcrE8xamF6H
Jnb0Revz/JDraWhIqH8m/RrVYRfrMbI/DUvJvpC3YbEjZzWHA05ED+mTIb58dwVjyN4zuS56DQjy
J3wUuAIPwJ/C0MtGF2hY20FwgEfeSSQLqBGS46GoGvyADhC8Apjv+sLHNzFBUWSrFEHdnKr7/RlY
CsqLxDPsp6qQD7b5tW0RFo8DUBQ1DnJCC0h2TG6lpasht8uKbgorMZXSk49+vpq+Wl6Qrq9BnxV0
XiuHqkTG0hzHRmXbwjSsSnnx6zTXUmFKBdeET6j8oH9XkRMxDWf5ohgC7ftb7mPKlctxAJ47dI+a
+WgJL1oVhGoMcoDVlNcY3swaPkyveMSsduaoKVSMwsSioJWHduE2jP6az0zDtvmtge3v72NkIQHY
TI1/enAHNLNqU9CrxlgmjNhIltZ0nydv/va9aDodQTqbGDnzALpPxCW7ZsiusYbb9II1R9j4O6O8
O3c4fSdkATM/KPqJSfT3ESdpovxs6Mvpcmjbj2FBYX3BhSKBikFYNFowTDIW5lnQMb1T2Kxw+VbN
SNUeGsnKxzVDsfjUXtRNNd7Y87cv8sDUQ6p1VNO3ume88Ea7Iu08Zm27C18CxrdI7lm9zkSzEnal
x6DCO7moBVuh4Qqo1A9E9cbeaccspfqgSUWt5j62ozpmj019biPM6jI6ydT80geoDiQxg6vK7WaS
aovhaZFScRyIUo9jOCGoKegTvcnFIjwK33uJTQvd17JLkj/q6zrZlVXqOcKNojJuUc+GoJ1+OXN5
Fy8iIX9yia/4HjugrQYQBiIY0ficmGFUSfWfO94fnwoshCZVCjkqneA08DJMpHWHG5zKLL64nOmU
MP2EtUnqSlnxyNaX+g1buaTf1obx5BpcdZEzJ42K6tMUDTOemZVN0dUkHl1T4WU7nETN75IMGelx
qTmfQfE1mS2Pnsat7K9TyigFuqzkc8K3veWDFcs6c0ap7CIHUNm6tiVXMAuRhwf7vHHUdc+wO1wA
GszZKULvM/0MwaSNJCCuTG1i1Tn8DXMe/P98KKAYovrxGPDOwkFP6l4Xf4b9IOGNt1OsDhvIhBAD
DQgoKmUAP1amLb149RAEav3KY4X98tPpT08RIS4F76ueiJj7IfEZl2wNqLpglzMDUAaj8f3Foxaf
g7aCCxSWEkynHErg0Gy8m8ZMSWLIv1GMYiauPc5vFVd8WZ8G1PzLjNBzczUOZpOAlkq4/wWr9IPu
5omiuJjNTuqG412t0+MyY6FGFan8yrXge/rKeMDaBssKTL9nL9bqlpavUoYK3anr0K34uv/1uGgU
psIVm9A32oufeEyhZpej4/MuIajvkX6rxEAoA9hi98q/WYtdkNigN3DwfWWejEP2Ag8c1eis/2mB
NcZoxtUCcSBD19VPjY76V1uW3VrXcz3bYiJoXfSAuMp9LlGEgsdRxljzVQ0fhF/YGrtJV6cS9tVu
2l1XryctYdD7GTAwedDHo/MLntPJ8dzaBVV4pjLJ+XtxJ0jSYgMbLCOLKD8Q5gBTCVWBuQ+SAgdj
cwn0hmvPQkEah5eKQSWezs0xZE2qUNWhb72CI7zYlDw7fuHiJyAztLP2vFPzs+wE3InwkWEwFOtv
EOMpLN4i9pLub5ypZxihEP1NKi6+ESKrVdwb/tBjZm4SnD+YSC0Gw7ExcptbowFX8sSkaaA34efJ
Eg7jUSswqhck/G7wId4Dx6PexDaRaagiWUW+2oN07u08gLmYSZ0GTsTC03mZhdC+Ermuk4IIyfrX
IkAwjV4z5bFpZUpKkfYQ06UhUbh4EpqFIrNI4WBnDtvdg6JAqTp7Tq2Iaopb/BAag45FHOXcclm0
wTPiELhhgMKCatetjbYneIwW4zknu2nh6eqY2afJlVXtNM37GPXjo9EexlMnLI+RGnLg7E4Rfec2
a3Ilg3pAUdVChvo04LZwovBmeqQ1iRCC8W9GwxcsuDrFLzElIgu8kFub5ArQQjShFaGV6RSuj/OZ
Ub++AjW3nkATybJLm/Hse+0XVjnE8WNTc2IaUx3kralolXYCGQaNgDRJsviuV3OE1/SYHRFJpjoL
txWIUjhCNO4rXsja/PjyWVjoz1VkTujihomGA3G12jbcgwq5ul0JLN/GLZBb9SCJJTzd4dJLoqvN
qrJ/CvzxnyPcr+NPsiBkcSZk2OPZn91ieh881m4BLNaolfZgJQndffhMZfPpOtX5tkjv7avZyBXX
vxrk76AGmCMsPblOPaOhnCNRTwUiYypOmeMvAcnsxmbWYm2Z0wzaf5n29+3H6k4vrghluPhsnli0
SYAl9lvzX3zT/Pif9QHboYCyVlSFkIaooFzXwXuSIVxn9dE3FmuPOGkiEFY83cq2TppBMiXpj1Nf
v0J8jEbefsuxGlcvLNDIZXAJ29nQHopTxiWHvTd0cvY3kKAwSzPSXsTVUB3G1de6pbRSV0RGQ/gI
rLvn8l5IfRUNJWTGEB34dGeD8mZRuSwgtPlWjPn/01BGASOXXps61pZl/eV+NWQeukhUatNCvomt
cGl0RYma23oxf8MacyvKXalVbbz+9Cb52MvAd5XH88CVWT0C4+Ddhg5C2E5CFh7EH+1HPPFhH58V
98jW+ajR5pF+NY1msuOjn1zzdY0X4T6QR8MdJXxL0tVtNjkPrxl9+cOVlXlobIGalM4NXE3WJ3pU
OxJgp262fOlqppow4gtGFsNLLpvDXcMEfFhPxZ2nIJDOeuhuUVcgbEcwd8PaOpVQ2QlswGrLeFEU
Yf5cMeI4XhrSVBj4rdMb59o6xpKDIO4Vu9eRYQQeJbwClccQf3O3JmuW6RAFFHg/3ij0xLBmZqOZ
XHCKwG/eGzNV9HILQMTQICdgTC7JqMMXtKjTvSa9wolyiWQ32jFLn+Sdl+LfJcBqm45FwOeutqVW
xgBQv5110FnzoKiWa05kAtDLjfupVeIRq5o6U9JLncdVvdItxzvgiLY1PNCPYNyRcs4XapZkXBPp
kjC+NHnvbCv3fofdCzX31z90E+5pfSQ3Y02PhTxje66nD7Di6n+S3tL3eRHDlMwSaZxnXCwwenti
3zDYZCf8Muon9GijqB7Q0kXp63cSW+nTxEpONZthFabvwobNZxCXegIh0UW58/fx1SoumP4lIBvi
VydlWrAZnxZcnmMQzCuhr+7uvzNXtxAfePG6zS4ClpEHY2PaK8VJfyWv4hxPV50O/1BLNZ8YWhJH
siDgevbXdChG/nXJj+/3JUw1HTTKID+0r33VdcVVwdh9iHk7YMFWyFA3UVw55UCyBjUPXv0asQHM
L7mdyeERvA3YJEo/JBxmdV6WrLshTrOLHLzVKGxa4gpCaHWARGCbivMjhvUfAZ6j+AnMbVs6YLEH
ekiNDaMmzvWCl4QnrVw7i+NNtlrGgh7eF/mL/g8TKvvtji8q8ZHnQfw2AUZSJbg6N9/Kz4XXKEpN
e6r1B5+nu95GT79rMyHmwzUXxnL6Zn8h4e66k8M4GCNs2XUnJZjQIflhyq+1gFp392kUXw6ko9yA
1z7jck1VMdr4i+t0AxzWKkrRLxXnRDgQZYn9PP9u/47stcjS3FD/ujASSpCQ9TXCiwIei7g/d8Si
+GjA9Sa3XktxcZrZHzHKeHkEn3uAaJ/YP7UKquz6n6n1sHF9ZhOdmT9Nv6I7hpdP75RG5y4zYQKW
zXE/u0mTO17AuTICsH7yoTuTWaiR0ODjZcO9q1WRRFaLqKJSV4GafBj4/3B1GV2fpvo6XTsJY5QH
V7Kzgkt4RnH7BPGv4658JqBD2RrPvSfUcLmhn5MGL1FTuyofgnxG8NLNhYVUIVvPJLfzQAyN5233
iQ1S62sBNVuxvW9835k7NdsFZvDqaB2MzGOMAKOA+3284kT/XCDYKoV1vd+hPYRJVER5M8Q4pQrU
U3XzSEMhL6JXj+VwrFS/nRuQAdAmOxa4o+dhQuhskQ508Tx/zvzzyv8CDBt9LBmd/Y4lz/dHjWFY
aQYZwMkN4EzjbBUejV7Vhkz7cJsYqOJy74yEqmFFqBaD7jQ7vDv2eP5bibOCfSoECHHqQ2MzXWFb
Y/maNzKkuLQRd3MMa7D1onfYjVgNJ2hWz1ovs0RJwikn3TcsUKkKpp3afp8ICFNvjymxgCx+rseN
qeKGr1kVHv2chFAaT8ds4Ljvvf+rooKD0RL7qUzQRUQlCOy38L1F9gPxF/yuamVVDlaiWVT+OQyM
owVmXpGDiPgD6ZbErsAOhwfkctTO4YSzMqvoJ81g/QlUweUwGc5jjLHetns7xx6GNaWoOMc4yMU8
c8IpmhIEDs5wo49E9xJOzUKcwBnRBVENDNUtZs/1HUBH3AYOOGh7wTXCf0quqqcTUBd2xE2Eo8Ux
YDQqNAj/es9L84EEFyT2piEcRJ9HSHkMrNuH7xLv7V5t08rMWcdgBQKYtoJz3nJt9Q9bVLsfPwbV
gCmogtVGDtZrfer9/kvu7EYOvJtr32Cx4Lxkn8cFDQqXye3pdDCETUY8eqGVJ3qbFGuApLV9X0CM
4m1yMn4ENyC/x349ZHoqGYIyiXZPQxmNaI4rq+Fc26bm+m28hed1uD+DIVrjDMfYo8DzTVkmhHjN
sXItnSkY5D7YoyGHucfXNrlKAw6sStdTQkmuuXXhaN07KGP7umUXx8yZyvxcWrdYS5SBF2NV3Fn5
bISB63T3au2ctu2yhSYQoyoN6ukdo73eSH7pw3Yzees7NiI88uKLu74KQHh1vAhsFjkQfa8kYiGl
H8fkX6ROdDfvg4qItlsQUIOa0Z3zR9vfAqzL9WhuywcV9r3BXmu0+Bq0ewR8YJU3fXygVrH6D+br
DMj/pBrRfcosdZLicEPhmg1LS+NBKrQ9Z0qGRn49b6AjBPsk4cNchCPve/xIoz7ho75faVm2V929
zLZMiKfS0IIkmaWi6T/BVI7fLelev8Zn5okhbTPyTEAtYZW40U3dH7DjghD8CZ+a3Bfzv/FYzC+z
4Fvrx0gXV7Yl3l97XMpWJ6wjWIKHT5tufKoXcJyY0lrg1HnfjuqNieARpvKQFvIFWkoanyW782kH
sp+Yw8zArDZTtfKEJAgKxegs+i76YFxjUOeHxuOqw/GRBAsXrFMUt51NGnvdeMh33CRv77j1at1F
B+eEcv0kzX/Vz5XWzoIOhnSGAcLAi0/y3KnuvIq0GCR89wCPK5JR1oqWzzpMWZ+AWxjk2lq1ygUW
oq3qOE6MBX1MHGixPNsSPsViZvQ4oA+N1fTyqMPVDzk6tu1PPHSY+llrh1MUR3sOOfNqw3C3t8FG
FuQORti4U1aPxgwM0vkRpNXxN1cSYsEgvVKP+I/ennIH1NiLMPS8xyzVWk0uoJVMB8tgo8P+N90J
BECxHHLEYgiD9SWy/eRJPUI9lby3qTYhF6AVtyNOvNOrunWzLuvWyFMVu4nRFtRDxCE7ETIHFMmH
F3OFnDx6jLlU+XcVOq15Gx9kg+GbF6+bfGzTs08aoU+TzzIEfGqUknRLU1Jl9jsz/xvnTap2zYJj
Dz58WkDgD3LnNHVGu8tIUZdCni/vN4sL/rQhs8aezL3hVti2Px9WPmXHom4CvMdVN4FRW3lqGJVv
Ju+lbWGueE7JxRL8WWCyEbc6+OmmxFz8heQdUV/yiTmctsxFuaxfOF8EsSZBKbx3c4L0+XPe7p4d
6k0AEWMqK2JbuQVuflNwGUCtiVGbRKVPdktmA3c+mNgd3uzaVREqFsUIzzUVe+Bu2Wkt0AcsOrfT
CnT+Xs+B0vEEkAxE1wU4vU9sez2jH5nYTcJWSeuiw8MoOkDma/i5u9TuLYNg1dUAowqfD4XaW3By
HbEIvryQr3OUzqkt1Env6RYj1EzXTyvIwcJmu8xoMnxJo0FR1eQdRav5wwlx17oy9DvkXgNHDBFO
NbLNSlPagEwe8Pqc8VhtQbtv9Bd76KmD8CU52lP4waWTKgafhO63SUpvkN/GKGonmTRfIoW2rCOt
wWEyF8Mr7im7cMNqpq+0EWRydXUWVmR7tv1wrFrEKbi3Qm1K7s5wn6eRp7ukMhwQp5PMQSXQxQ+d
blKRjuqlKD9IIqMRnS9jfggbGN8sE914hAsacrUERtDOts8RGWcsswuy1Mo5ek73cT5iJg3Bll/W
xKluW0ZAAOg/Gbl6ZpC/QYUWaKyw5GOMSb1YTCMMIcGfyXGdrusuz8TIW7zOXRlRVP9TtcuzSFtM
2arlEN8GguNV00tejinJbv69BM7CsnVzM7LUQMaNBVyQASbnztfbMRpQCQYUjv+4/q1jSUBPMVwt
qegP6djGMR0L6WW7YFmXNLu2Vh+Eh/5Ew5j6Ii3RVPlYIuM9S1cSWCtCdsq5NnHAIyRmph6TM5lp
OCMdTrxOLuEUr5dVJ4jaTEuUROBMnSyARSEhhCIhmpNbGzK1cJfVykD031Gnq7plJQMGx7k+EsSV
zib0Vmkhb1oLh2iYaiPKwLau1DW9bI+vBVhEBHBO6IK6VqBeow13/0JYRVwPMp935xCowcR9vEBR
QblK1kVTpVrumyesdJIlOC4Uf7kvJD7mud1TI6FWmwqvM3xh5rnpCQYB0m5g9ZwcQfcHNvyal9dl
Skc5n65Hn1e/VixX5HKKKsoAIR49UeoW+jQCWVqWIgXjZoWXrdYQdeVOF5ij8xhh2XNcFyIbeTJw
4JjEZVV56ov/Y5zxhcl8fg/iZ9ciGsCU9pKlPNJ86ZuBcR6ynbITCRivAQMUtc1kRkyPNTsdeo1P
rrc2yJdKks1G61xFgJrghNeruAp4+TnvW7f9bW8vYI0MGI26T3KGnczDJlOPr06v1cOsaZxIkGlg
8GmWrUnxhqXINhOFy0oP83uMRNe7m19/AyNfK6I+PH061E3xVz/6JgvpfUFtKcNbByNKTCXVpuI3
+QtV5OpbwMocSRBojAN/uoOZ4mCW9WjCyj+6TV0jnCrd6oGfFKW2rfPZ70WHEURgEpcItZkO1lfr
mzuTb7xNklonxiluj8UuBhkmMqlGwONOAdgWFQEYXzZ4QM04tpqZ8baUZtmB6pWYtCnwTikfta5/
9+KuMkR9TviFY7HUNVTheBsSGfNNsCutuIqfEJACCKJN56ORR83LJAvjAS3YaX3NnwLxQolbZQJs
88wKKqSkfarESrBTbQ29PuZa5Uzn1LLhT9map3vRoERVq6b4dprpBMPrsrTnBMB5RWgRzqrgDHA8
a80MsU1GhfJTkMeVhQTvYwhfdJxsvsqoELFkLZkHuKPHS7hGuGaX/vKVWCS6dQBBrDGCLQ7FMVQc
LFFJANsVxItatHBHWmwtRP1bQ0sBJQUddM+P3y0cJleYMq1/WYyrtrhTMK7x31SAjdf0ERhN+I8I
6kmeeJrslEEAnrk6Jq4LzVFBZF49h+lnwurNUAnXFrUnYhppYxv2UdzabDGDxs5K+oXlkRrDV16i
M4ckwMlqmNds5Fm+o7EhoutPVmSAswg8oR/6WvvMq1Y2ZU9Mpiz5gc87gCp7q5atDXPDeQYdbx6T
WJIJybznGuGxZQvSWyspvtrmDa7l6ZuJ8Vkd92Qppj82ICfTR/TZoQHQXoO3gn1XAk9nQLoyEgTg
GRYDvVpcW9WmskkcjMsM+A0d+1hnzX9uxi9nq2ryPWo2OvUv3bPfTUv6WHAMeGJ1oNvxJShvmqP1
sa4LjRCPzx7vXARNInJ1WFn28CROyXlwhx9z65a5WxQQBoYdIWPSS/zMVgN2oCTxpg18yL4y8rvh
9wVmwZjqT5DqqkcuGwRiZnhbOHZzRjcB3bRcCGpIeC5Bav6e+EGeRe2ndw1V4S0o9tyIerDIzqBj
NKRtxM7Mj5ekMJz9iWylOiiRldjvaPuLdDUXiUuaKDIP70T8iIIP0jgsiGg4xt1pi7YJRKhcjWr6
61y6spixwCjIkqWEgIR8caGVtetImvCO6CUEh836vM5gNlyiiNs/iB4OCiAkWP4sSC3RIlL3DeO/
WxRNWDi0FPR54iUZcF0Hhn/PQe5SK2WRrtqMtXC8JZQnEwmMJL03t2cA/+uLKpkipxopcS8PxLzs
M1vxFSu+vJJwbAL/CQNeNbzn9btcrQCh1eO9BMQ9GA0fKl3pDO25Dp/7d1aMf3OfjgM8GyFcAz6R
wQx4u/tOTzTn060AM/bJMBN2VOKmQbtncRWRLEvKktZQeI4HBhqqJP8T6zM0XBmf6U/p688rt60F
RG93Rqw3UKOKBkGZSyy3fq6b34eXnXzLBJx3I98X04OCpDfjmcJ/x3dR3hoC2+64ByUkBYsYZiwE
+OU8GMqExgi+XrdX8soAhbp5UvkyJxvvOjxDRCR6Qk0Xz04uNFov3ZUZu9gIIOusKuwiyO5L83Ki
axXvAZ0ph7g+g3QAnK37RTICMRUcamxI13YDl5piJ6sf4LRWgZZ5rUKoIIOol2FgpZYLL9D7pci3
JLTq/fkA/QcnpAIR/nQN8sQHrzyhtbKGOr/7xn2fkLeKbZw6tml84PJnBDlXk9UYrBIMMEpXawy2
vEJnp+1zHJj/sD3icfSxH0YNG8NDzwqD8ERfcN99ggVNQlvmCmfXD/7/G70/6VsLEn9CuJwnhruj
lPSnZDYekDEYlPjOAo4GtDovEZAJubHC0GRXmXeba7Gn8T1wEayDR7LrqqD8KZIoMVdkDTyRmhto
Y+9t/UPcU004rY1e/Zx0MNV/zyYuYJRoKBVGICZ5xRhxNbgl6kylxmgOQoaEDipF6iR5t3GZplwo
ZoxpXNk+ctTsfAwD18cMfy/iedyn3pTZ9Hkf++v45/S2shnU+Fg44a4O3BDEVH+1xAxQ3fynTPFk
uAI3nDLzpLULh9vhS0ijmWCBLWYfC1UNTPdG1/DE31wWoLYqdeUUZeg0IlMmQvlkrtAGEQy8R2if
KaXWqw+dahudLDbZPDM3k9/keNqDOZM6aR87gLJgI9tv81oC0nxCElvB034WcR/w2HIixmQEtVdl
90wobZJcHy5ehUs++uMaGrfckZQFAPruSznGIQySA8wQrw6LKzdmbyJqIQqK6qUFZJtLbWTTGQvJ
vyC7yGeWNL2YzQsn/GX6F7lUwgBloMwb92QWmYGS5WZAhLefAnC8jQid2B0952kGh66BrnaqL0UZ
E8XDnTqWV89yrkWPdL4zAntYmOYDqZucN/4Un8IK8RBEn2jbqQHGaFLX0+d8oOEOJJ01/JXR2z1L
/nW0LgQDlObQQ3PNKBDss7wTmwuFweVEUuvtIjxCpkvZLZJiGpncj2CxS2gVlKgvAGxrHzquo6CT
Gv1G+Aj+WY+DEt4oFXodbyApFUr0urvANXifcVzF1ORCGIeIMtMA77ffhbiGowSuOxazNqLbeaNj
f7CgVp+1ZxCpjGgMPB/Au1eYh3/o1CFv4p8RaRSZjYCOHrCNlfUsQ9uZnWX+v6yfQhZpeVvd3YiZ
kg3XEYwLp75VGdYHgsb4p6fqWAbtieDkRTmhVBI+nM1dadnK/xCUqFkEB1jCy/KR4G0ROJ1kIxZG
smINe1QP2vh997GMN9DSpgEnaD6eQxW/Qb2B8fu/VHpkRLgYUsO16FOZbqgyIvnlP2hCaRZOrtE7
3ssgnJxHGr2zShJQAJg7pnz+RcZJup97YlUDFBcWOtWd9VRYVrhzSQhlJ173xu1P41NGFVrwRBNN
CpJjVN8AAP5O1//IYhRq/dZCBNsv3kZgvYqApvuUV9giKe2hb7qjJn6+K+7/BJh6AE1qvhM/+Xip
WYiLMZceVARH5xBnLl+DDKybRXUiGOUTVaM+V4FnsFnDpexXV0FmQipNs2FQpAIt3pI2QMzaOGFH
ADGFe6TgRmWEVOkS6sHIfvp5Z29AshXxilE4FvnBsymXOC9eAQHfOviCnee+2UwMNIZFQqgKo0Ym
quQ3fcyHjj4N9w4H1eRTIKPcAYTT3I4Wi+nsrivJwlTI9sGPLQYI9emot9WCfkypCdX2MXjpM7JY
5f9ZgbVaGpvt8ZhR0hIybj+VWIXczNl0f7V812+/QY5JSbxgyMLvY914+E43X37LxeJX8EADWMx/
LG2D35sal060u4x1bpIfGc36mVriZs+Z6jngUi/+DJaT+kusXvzKnzAYYyYyC2jPLOJAN866fUIx
suHujmSV/GljYQZCv1OCdAvFo5eBgcQfxB4Yg7URKaGpzKiSiTYZxTy9gVDIB12/dfnYGeDYyJiz
Pph1X3hFq0Xauw9nbJHXZAkhV/+mxqmTR/+86NwiB5xxtXFTFhY2QpxCy1lemmGXDDKKbIUV25jl
GTt0q6YlR3735wzEkDGqN3fHZyd92ofEWTO1pDTRGhITfgiDQJhsKF/437EwzCiCzj++dkZWCmwa
AmqK2DefeWF1bE7KITbsO2ZyxJA9xOdr5Fq5ra3p1/1/PqdBVZ8PN7MPhpFyHTyseK5tshezSUEr
rkTs3ZzJvpPPRewBYCM1IOfEnMU6Fdq9L3H1coLYD6H0KwLwsNNgUxTwl3AtGcyu/p4m4Xid2/us
AxcKI7fH73vCUZvq29Wn3vcLKNGx/wvXOOOC8FgTrWzPCBtkibX3ERlrGQhtP9a5fjVvJPvqwxjT
mI3bMOChw3S5uR9ezs+2opsV/6HEvq9MOR/qBN7nTtFu5kscdozcq2ZlVC4IHYG5RRUVg5PDNMqe
Oq8nQqDE0BLRfBiGf7KPhLMgw/vaO4Ln+NfMraWe15NuzmbAQ3qdvnKAjTSRx7A+1EHevag7VV0J
QJh0m37Wa2IHc7ew9KgiANk4B05xbzy9yUoPkg/Lo2qWi1tKEY4ImCpU9SMMSQrvY2KTOh4bOMCB
ji+fbtmQR82yn5ovjLVp6TL3aism2BjEZMxEG1UHyr0HrFhafq0b+l1bJJjMIGbn9rTsLyZWAmmA
F+xjwA0108rOyJsBNA6xiNGABkTaRdj1Axcr8XQSg3bgchxTq9+32q7WLMx7Cxh9jXD1QF8X8UMu
LUXC+IKQCG2LQPI51Loqczv7bsjU1U08u73wEHBK1VN1Z0fOaeZURyijPVVQ9PUqzI4kLuQ+aU2D
6XuTMtx62pc1vHtbE7VQYLX6kTMC/HB0PT2WYTn9lGpFImy5J3rHJT9xe/AtB61Bh4ozw7uI/Hre
KbBziMyypBk/TmUWgcbxrG8mvZErXe+AiSCc4vqu67xRamck34pBpqLAfW5sn+bVkElSKAxtQx9y
zhosbqI/Q+MJ1hqcwHiMG+9HkGf+JhvpOvhTOt8cFuVip4l1Kv0EIVGzWeW6LdWpeDSjDWdpCMVP
pDQ2rV/vf+P0AyqVrqgvw9TwqLsLBgCEoFtjz5rvtikSP97nMDX8dHgTBhPC598dzFNk5i31fymt
zKBCbGfI2+b4JK7TsQystqmCYOVMCzebTP4fKrOToG6kCGZixOHiQdaEYbOsOGFdAJrtpVbvGI0/
J8a4ReL+yFVFUr7jLydbbsuLVmQEHz2u3c480cLjKc5Ln1JepgM5oPoMGtMrZOMvCyozhqgrVdjp
1ga/ZIxRauIA7kOhEw+36EpCvkUVg9wfcRka/EQbplDjWkNvySd8PLJBGWM9DJmb9ZeFPQ5rYca+
dxY2abnD3Zq9HgH/Zy5eXJPBDCSeFxus4Gs/P99sZuPyoXYUQ0Q0zGfrECjSyferTgVi/2gCP3jl
mqKADc1SG2WojC8TS1Og2jq9KcXYT8DUyddUQD7qR83uAWq0i5KYCHGMlL5DSWUdLn7uQORHo/20
QNYTpdSGYjEVnnkYqpzYwVXmT1jd7R7VnSPY7SJW6DOmlQwSdhq4h+mLWM4kdjuVS63qpFarogd7
2F3LxOpsLdCETO07xQU2Q23xMvBGvJO6yLPN8yDPt4XFGglL9EIZV4ea/rqKkKMkBzu7XYvE+s7I
78yzDHQSgxkKXrT4M/8Q2s52bK32qwt4e9ByA4F6hYQT8LjA5YDbTqapwNn5BnVpSx706BDgr0Uw
QkDfpSyeGA4uj91nGJBC90ty7DdzyGdEE91XcBUMbJG56AqidHVjtbxRWUo4e8FT3Cl4u6gsx0/t
420o9xukAYnsvW+rz2ndEAEQb2CrAp9oFFRK79hpN0WqVbsSh9yzpYeKhi0NB+sOqVu7QDjb9wS7
nQTc+hfgvuEhRr7gPmNTLd3pyu/9VpVXiSUJB7wrQPBrhzdvedtreDaRKV91xEpiFS/NBa3J6PV8
e+unufIBsY0u5lGKGd3PcGz+riB8tcrtpUPrLiZQrJh90+JLMsV7yYgGMMIKoK4r1w/VQyzHcc2a
UJmQyw8aM301rRveP4aBnoIAriN2zteQx5BJyatwb6jlD8OQADaWQkLRhQpv8l7O0fVRRVPhPRYa
hMPtCkdHHwlvMmR2J7nspgNnTVTaa6ILPuRjqv2MJ2oIo50ZLwRrHaJs+Z4srrYcs5uyrNJF4se/
ja2wM6K2dQSHXFoU/pm7L4150Bh2hRgLg99uPwv994Rt8Njs9LyH6Ur+nDbewuzM/Alcnb6+dNJb
/4EbqA9Ub3D5xJvzjL2vXxMhbybCXNmLaKQyg8UJqQ/eha20lttwD7I3n/Ykzp2Aq1S3dSGOPXRx
MzokCxm3ZtuWdytORXRkU/Lu/OhtT+SScj8+fcStiqAUtFG/vnCZRuANpLh3ryKbomt7rtB6NgBn
XEVW8s82mGAIhqYMbNPsc6agrUqC14TAzg45JDyu5UKDi6zOKx/R/EXoz/Jt5kwEiodDFqL/X+tZ
da4SQA12yVSkZxqV5gDnQElaDWyAsLE7DeCJiqzTpLP8kwbRBm+ArXjgd/6DDCfQWg6L3fHQUXsF
3mnadaIY7XkrcjiSt/TJod0s/DxHzDhQtvciAtURFSHM2rFV+vWVlurA7nkzf7KuHCpIEv7r2Fbe
s7HY3OfvTE3KTIrQYVPUgdYiqjvcbwy5H7WEh60G9dyLQFSAkvhJKiXQ4s1xqj8vGN6qxAn3zM9O
fwNDg8jWaaEV/97UyGLLB6sI+ERweLsGXhPwfP/PJTBcZUicELDKQ9Z/LPcXTmFEsW8AUdfPhYh8
ddPAostPf/lqH9PuILdCDRzPb7fImf3LsU7bEhOfsZsRY/n52i7SugES87XxGP2q6FAgl/Z3lxAq
V+LOU+uaWAhd/Kfz9x/i5lov+1NxEAZzrlNBQwc6mwiuz8qUFwjQ5Ff3Yw6otZnK+5FE/Zr4VgbA
jrTYzI8/tmhPAP6jHtp6f288vhzt2AhNE91+OOUjD6v4QSlLUcjhh7eXeZM/vgtYHUbMDpG6pAQR
J8q8sc79CoQ3u7n8oKJJ/g1/xvJfQDtHCTGqO3/kUvD7PpDYBXomGjECP0y78uZQlQ2yF3PhCy6k
NDz1Zzoub18zmt1FilCqkvMC49f+zF2G24pBjgOHPya4c2YnLymPoGiSXEuJhPpOVlGjcK4D7KUF
Y+shVeGJF6ru0G/Q7vW9FXjDW3J9QGPUITtLjZwi9R4ZQicX3qCDqfecxWk++9wTj7Nt7oEE9cz2
BiNzD952A/g2dIpOj/vG+Ppm1C28zqMUNh4Om01W57hQk+yI2GtMRS5HHeWK5oxEjhAMqvErFGu2
BsNVoY+QdxNDkXTV5DzUwWXDIjtP7mlqdHMkUlSSXFzAweXuc3RU2qs6AOujh6PHjoqNbtlNN8om
ePL4eqyitjPOIcW6hBb3b2ohQjG7bke/g7sg/gyslqCeK+5ZZvrdQCT4JUsAJv2QWiWvMkdB7nWs
seTmC/MTQUZw8Ih0NcQ24mW8ka91Fx6lzCkhbjNcLUqWOKm0z65OfqUqj1T7SoUmx9jpTQCdIu07
RR7iVF+kzUZ7rr69wPiLoe6XD7E3RHoTxJ7TKyKo4De6fE9j+oLzLn2qHPATge+4yHdOV5iGItc9
MIWp+i3h+c4O/z7QZCTrvZ/XmyUJ4xaP1eXlLceXWx5Wh6fdZ34za+qbkSmJ/MWZkVSU1DiymrfO
Ow7YXAveHtNOgP7lwxsk6a/r9M5JF6ee2TFfxJyXiukZZL26x87OPCkC/LbHSLR9st04JozRlpX8
2FS9W4VQVnDuL5KQIB+yi5okxrPyz4RhnJajxJo0MHdjmKqqPjtZQoUfYmePh5kHsxlDQ42F8Qxn
6Hw9CS08g5gUwjFbuboGRnofs1sOAvQH/dv0sXCeM4Hnhh3Fh9XmQobeCjhaC+7YYa/TS2VNqrsY
Q8S2jcOYt2arhpoO8OEZClkmDqYG1sDVhRatw6TpR6w+UgbCtEfNJncrzS+hFuTH8RNMec8HxpS8
aaiGiBPUE1TTIeX4pHo0qSB83Q0DvHrfGE5YAEuYmhMStSyOUd0ys8F2P1dUkdukQ44jbFBQr1dy
FWG/J5lA7BxbQ9iXqPIAl4nun4sZfvZxLcHSOayhAGmJgS0qCoJyFzNYKkq6wpFvw+TJAYP7zPu4
menE24hV4Wa5A2H2Eyr7Bf8f0TvAmhEgc8tfNanpjZNynNi2mbb9cTQa7SxIP1yLdafE/PrUIPJO
5L/zbusMSRXfs1hp2BCPecdz73lXs5ymnEBNXwzxmh5xIIjQFZDZ8QcKjQUYubFhMD3HWTWHZnCb
qXNYLs6r3ezeVS6Q6Ax+e3fdwofHVbVDcklhGTcKUDZUVv8jUfY+tPBksvL+4UIPXNegLUcL/bTw
RDY/bKHtiNOMh2tN3lGuzgiMwQhWvszC3+lS343aj4XRycgqI7lTkSBaDsAeb6eXmahKlVKYnx1M
6Qej53d0hfuTQHrnPmqFj7Iy70boFpdaUST80F26YzDcvu0NEhATnWUcbGnxbhC/9bH8njz+y5Gf
W4XAo2kOMI//s7wsbVGSmcXVQNqoRCWPiPYW/EREVq7mOXuzm1R5/vApIWhlzl8pmKVPONz+lUhv
P9lT3BYamWDTzRqkpBNgSjZnKLdfLMjJViUHANwdwPS1X/rMVRgBvQupUhAL7XKUJBt2AY0KcM30
ZBcoGEQWRqnrshf2NdbWUDakFPJivVDlIZUN7LMkMlKQaQD92i9ULyMM9alLNKcCB6/CP3yBjOad
Lry5WRsikHt84oMoObyMJMf6FBxUJLR5W++9fGmpq1Wm/EGR5NYFCeBLY5NMIrVX66ZalANhp/2C
LcsePM06lZQGM+LD8sv2YhhT1+IjQJxiyMphzfUToIaFJCmRLwjTC+WMM323nOuFi2W7Hz3xSyAL
1H8WzKgXGGCB5E/L+AyaQlbNRK9eylpt7uzrcPZ58HfFDahOTOmkDLAMOAueCxbVyJQXHG5GwyOI
sCkv3hm633NQY7qnUfomLabg7Ayf4UnV8716ZMp/UqaDFYqD399sAtUKeJsAb96Kgjbs0nnAX6Td
dr9FCktX4t7zcDK+gqHnAYfZlRVQH2oam0PEflA8Uxo7xdkRaHbjNElFcGmQ1wOMT/kqwTEf8yRr
lJtfy4sv5jjrbV5nNFOlfWqW0KafheBXW6Vl7sCeMoy5bicd+Tek7mBIo+CLhdydI95e0n9pZfqj
wgoErUjIp+zdHhGpG/GIL6d4FSM5PvWYiD74LWMaSJ6nGJfr3gYPv+GiGM4AaxnwSUjmSx0W5Ygj
65fyRJRViFs5+nWlDTjdoHLKoCxm7zLy3j6qs12UDCNuOFFzOQdKgqwr0VZ26gq3mXs8WOfdBCXg
gOgdgn9JK8VsFfYnlvz30pCLxE3IWXpriLwnvY3m2KgcP2AJLWFUdC4V6CAW2zlhdVkCK2TYxF8t
10MMpsi3s2qmvANCMBIA8jv7lNE10ix1weNKG3L8xOaq38ebsZbXHy28xjrQrjbSJNDktfBH9Iw2
epXtrMbuWT11WddJT4C6w5qYf2pSBdBvnusdhEaptPNzEzsQv2frKgQOZyNKKjVTKgvDohmIntPN
YmFMFBp1Hbtw3FUc04D0zhaphHzgTgpqZK5fkSrgcJFTZMeMjKpbhqQ+bS4lizVxWgHe9z7RPtSM
MGCTxdpEZAy9DEDsAfu5vJGNmvpnUXK1+vmMRgokVh9TxMdJr6ixDkgk/ixljM/b08PY3ksVHD+2
teEEaljhBOQ/JYSmyYLXKPh8jDg/dMKbfGXWHoqhTgIbgp3sfWXAguZv9uQsKz5Bg7DGGYSxrGMd
efsVLemPUvjUEo7a0tgREnjdRn8OUM22pra9WHdctL5sCuqWwIi4Y7L+DdAdUnh/xbetcCsS0IAW
30u5YOYyVEZRusUAA4dXDKSzAPoUH3m7FdYn+21hs8O+RK4H0WAFBslLaBafwcDnp3bMGUpDbbLd
E/ynmAS94UHlRCNTD0bYBYVkJf4C12hZ4mcInGZ83mNWwLzDLRFj5XW6WDOscxJgHgCU1Z2w6ccd
uU50f9Y2D3rxlGP/D+zR5esEwpJhNDlVTJMAcO7ui5YpMvByhJulGO2Xk7SBfdpsR2iIet+vCP1p
h1vIgAPrxV9tkQYjG7Q+mX+PJpcNmlMPianFgBDfwLA6eiaG+o9A9slun3+Hl+pIqH91oaGRZ3mL
+DbX4AhWScL3o+ZHkLCaZvNbJawxHMbJFu8Ujcv8VCnwVmp+zL3k7mFzFVY/EE8FOQ8S5flEiEzV
+e7C7M2fMTwMstCTXwq9k09lWATzcb43x53mGRb1LuZ6F4C+voNNuGOqX6e07sD5wNlNSVmzYQ9Z
DF9nKti7lvly5D8tCLs9q78QLWZEwv27KDzHqVq16Q5zOnr/OEqc/clGL1PaLodPvMMS6OUd+M6u
Ug8u7UxmOju3RkC8L5xv7AVuB/YVtBpLMk3pWAr0UWDF6k2qBnjXtTgzuQpz8l8gnC/Ze9PlK0Kq
oAXbfpwRG+NLAWrIBKFHGRPRsa6xNnGf1LPKJhRZ0Hicv2isoxAUmvG2Hng4U8aRSSVDLPxyvfvA
EJio+uKqVh/Ye3X1w+wc6bCW7LvfPZbV7BYj0GviIuUAZ6lBRjMqnBV4keU19D2nChWRMa47thFk
0SbvYxpi32V9KEdupMWHzbJaH0d6Rdl2/JTLTx00xOkOJN+u9lR+fjCE7iY8iYDigWi7KBgpL5wa
fU9EXvqnkIZ7DQQPZZ+4u22uTmRv011N1R/Qk4cM9y0cRtttApMpSbUF3CB7jQBDUl8xwUFJXTDq
A0zV3pYnGaqTNXUIAAv+vohn94aT4ywumJtM38GdHqDUpC7L1OL5UeAPa5mj/P9FUDMfSqrr1dfi
fNG71LB7RIdnVl0a3do5U2AeGr84SR19gmeLLkMlFoQ+pOyLJyVejEnJiKvXY/EaShKyFYdXmZHv
0exRo8hf3Hs4b2Z3v26RhJ1/ZEq0x+5Er2qaHJdJsOD5TuMnOVlvQZR/17jGi3ngtiLUnyw+uBGs
kbRDGzsziElnRlsTrqn5siO8E4aSzHotsGl43GBNNn9Zu66bZg6q6Z1la61O3+KajhThK/fLSlSb
R1x/UaXEKMjtC/CgYMKsGVsT7/j09HoUf8sgJGgS6YmlpBSpgnrG22uMCqxtcOkFHItU69ARQN+P
ma0Av2kshLkmQgXcxx3k1kMTrLDqK3BWpJvw2Kpt7ckjiVMdIevJQRpGcXnP6itPS9HNACmpESD2
USWkA5BSc68P8ypd1XNPkU+pMvPskxXUHP0mijyrkltT1E7JlzNh7fJFsYyOE3RxN4aUcjtNbKSS
hsfumZgX3tqop1snEN5EIEW7v6xfQBS5rqFahfMuxjbWrFhVC51p0WqC1yi8kWYEfsBq63UnJyMl
a59Obhb980tTTisOX1gA+oqcenky1jiQ17UOHXCgdzGeLehovIISaTMjT+9D6yErm8Aue6kcLy0L
X7sb5WWhXnqqAZoBJRAA8/H94WfdXZqQhv5ifCiSS3dkeicxHT1CB43sK3TkB4jQxs+p+bFJLCM0
QZObjbIXr7gTTqyA+nwI7uWaPKe0htkkQ2FBG2COr6OX/65C44l8qutyHs9AWS2Is5Rf/IsbmOdS
D8fHBx0IEs4DJYSxsiDMm5ShKBtRkvktR5jEKIZY3p55aTNRRaOkOizte9/8VEBUrnk0cmuK+D5p
9mvmh+HuJ8pOgHXNwNbApEg7nW+v2TkcPgvpD4de4gJl08F2lYtJjIyrMpdnZ0Cvkvdms/mfVA36
Le2KC4cUxlwtAmUVR7bhv6SHX6uGJhjo3i5jBj0vGqgR7BycmnQephZnI6ZwkLJYRe4XLot2bXrx
rWNDmsdNj7eAhW0zd1lHIq/oz3CYGwrae/x8cpss3Np73kGbBMdSYyGKywoGgxzAQh0EwL6CyrsJ
1JAJk9DJYraaV8pkXo51Q6bzGlScq7UQRUsXZqXp4OnZugidAr1OCtSa0SxfiSFqn8X4DOygBX4I
12jOoJ3qwTX3iZ0xvKFCNOZgoxOq3GwNSjFCEqfd9861gRN3QyLl7doQfCKgX78+VsCkU2c1tI+u
J9P/RDdfnq5rX6gbvBVQVr2rEeuGcCGj2Vrg4rCaatn286GC53gVudGa5Fp9exVPqmN6x3oqyZ8o
Iw0hUCNd0PVU+Y4X/p6UU2Hfgl8FAZiCCWPo21uZiHlkgP4CXwrQHJxFBiBpCZFgsIbFV7geR4MR
L2r/QuQFYUGMYxQC+K1JN9zwn6KNqPd4c3LbFQK/1+fCKHp4LInH3Ms4hdw03TQWESwR0WR9Ecrq
NE3FnjYSuJ9xirPcvhXK5JnxZ44eoayj0bh4eBDCYkCzATbJ9Pbd/DPQSDXsoFknpH4cOnEhR+XM
DK9aJpVvLzOQwCk3y8WLHofQxkKDQUKJxUz0NuZbXfeEW+zpN0p+JChSHfoxLsCAjb5O1GtxVVIM
j4tqCuio6V6ITYNyxbd5UTNrEUfrlQLCFVAC9Y7o9/Mo63SQ8XTQbXh6OzUdrOT/0RRVNhd1Gbye
FxRW6mbeP6EAihkxIe6f9UDTMfgPwVFgmwV7QbDixoWdb47hcmoLXvJZYHylEMeu90foRtEbzhaI
+JttaXAse5qFd95cUpSEl82TwU5IQBnEMLSnpvssJSM2cKJ4SB9PMapbxAQVjdA4pq9aizWhLTFk
+7zLYbhJ3oM9B7oi17swlL67/XneTgAhr7GssfazwWGJ+FpDqaXKnH4TIkGo8Hu0Jh0WKt4y1S5e
jjVgxIGm3c8YSDXZ9WdRl+sqwZxasQkl5jRpYDTcDYYkEqHD6hJvleWpbxEkoLiC/0yTctNR/Vah
o1/LqX/p2yNEqdH6gLSHAAjwxQgmfK1IGZcwgl1MAiTanm4MX5xVtt4R8kkeenVxB23jBagqROU1
lTx5khGW/rd4XXJVj4/d72tsMXx1jXyL2TBYP81djyqHgFvdFWfz231MxUYmw5fkL63F5nTJnMLo
9pdz4dvfHpB4v+4KewqK3+IIxLpCOxzW+2kCnNQtSBv+fohL+l8Gd4AYgwub49g/4bk1TaDg3t6d
akHh6b/i92iYsf9BaMdCv/wYYeSlLBwOQHVXR4LCPSsKek2XmS65NbvHjXfPWwtdDnJv0UASGopk
xtd3fB/hjttXEPK9uC3j8SYt3lfq2jwd9EE1ZaoUK3PV4OYY2ZZsA/Q5zqoYJorYrVPHsA+eBEuV
bnOG4dTwy4nO/S8GvdWDki51uVZSHqUc/6FPMa/TLHy0vQ4Q4sI7dvK8AcsGbTgh4d91JO/9DMtV
nRVN/78mxvOEzflYp7zczrjDmIqauiAYGnS9PKtQaVyX7xrdD5fHyeGxEMEd0HO3srbf0cRjjo57
NGWIjqx5iypl2964NFaucrG3MRTRa2z6y88YjHjKMC4j7wwOYORpwvAKMFB/1su+2ufVyCpnCtz+
osES3KYAd2SEh2k1NZHgkvn2yYmJjY+JPgIq43rezAOqk0xDuLDLmumqQgtc+xHNdau9o1zvBhHw
jFeKlZ27aMJk2A4EVbtcMOmuOk1Ep/Js7ZXIZUA36Yl28CN/T9ei3P+r6d/6MA7eXzW6WILocKmU
8mcZYl+54ZarW5rREBiW1LEKJTmQrgg+zSdm0o1UoGnM82Jpz/yylbhe610pwNuRs7CZY2nFfCy7
yVjc4fz6+QhQ7JAcSCZotNOX9X1l5hPa1125g9EhoL2tCGucQrFsxckczDLQrnygGyKXz3y4WKXy
Ud7OAGC2/1Ze7WoR8I2DLXaoeG7yJVRlFtewmdkvAUtDbJrBT4P1kAklDPOdb6mpsWV6e8RGY022
AD0DPajKh6A7/8YhQiRntRL68VA+NxRTwU1DpPV1QqotiTtEmo5ATeDeyWT57nLBlhLRd1MNAQ/q
f9O4G5b1xqQkljGsteCLjzyBKS0+cYA16KTNWCb5l39MZbAlPQ2LbnGXbj4/Bb2dIVPyWuMtHOum
Rvtj4WSRJp4Io3Kr+T317cdLQnbxrmv7XQ98HGZzc59rVIB/lU5N+3CQKnA+4LpYDBPxdV+DOWy1
dnczAu5OnHHA9YLnFa7GSKiIamGn2jiUTQk5q3o/3de35gfFSZHCbCQ6e9/TuhN5S7QyO6THjTjs
SqxiA9lE1EbQ15lGxK8t3rv7MPLobBFkSMI/hUC1tC0n6mCpdWvGLIeE8dGKjJvsGo0mt+wXKb3L
4a0BzhUlfzx+B46YpPVQnMzGNYrzfq+7w0SiBanrSEwSspEIlOSS1AYyuB6/Ndqm/bFmfyycv2cc
CeUHUaFcamzrrhFR0aZM42JPSEgQodwuSMttMNwONbzcsVEHKO7QqfuvWVrZy2KSV/emEjXclFYF
MNUV8lsEyzERzj0ph9XZyTPeqyjHpL0zhKaOk9+k7zNnuOyl/tB77ALLeEnShRzwDdXgnUTNbE9R
RyKDLpfP3alT7pdNP8FhwaKz2ga1S4EyLvR62U4oTwS/6Uqb90tbVcHXPYTsg8LVl6vg6gkA8POL
hlcb6b06kQqss9ie6s7Jedz8JE6SgdULdd0UJpSIknePiikyo2cW0kd9a88JOjscf6wWIZX6X70o
sP5p0rx1Jcu1g8WyBPf551SFuyguppbScpZSkVclI9cpuLefjuJBJOoVdWuGm/xZfStoztkubVlQ
a2VqX0Wp3UkXd6CXhMVx5yvWem48BoRczmlFtfQFaMUaKcZ2mSbMeUgMBCCNbGpG9ceh5nodkuf2
oVte72OKCAiPd18dRcq2MRzGO9dz/kkzL4ztJ97S3B+nM1x0VTKPQz8xVeGEZzziztORyZh+eo0m
kb8S6UDG59NsEYasTlap6aQGPoPzHgVaBc2tXKbbNf9yhxq3eId6wYF2s8BLzvydZxmJtRDFAh48
ypg0k3W+OQh1y/m9SnTSSikMCINQfzAucdI7E+i3sGPfHgW4Jz4rGCkKa3yYjzDjeWU+Ybc/1f5j
cx8ZYqt3GAxjU7mBfOjUZSWX3juk3LAJ+Dwqbf48f8QgOzEbyaeo5aAEtFlrp05VEfzZB658OYcj
fuUUfQJGU3G+dM9EuRu7lh96SYuebYlakodwEWsiqvjRzC1P3rnF9nrNmXWBuwK7mr4vTs0agezu
75uSU2SZwQ3Ei13Jj+bviZPexcC1t1skpDxg5uGitABUnFDH56SqCkr3Vn/pW1hrXSTU74opLVsw
erjaMiuveR2edYPDgfk6/zzvAzxdUl4lbro9RVKOIepjwDSQvEFTrb3buHsHAIvbmGtk5+alN2Ls
Hax0AoiMPKimrwSi3f6Udhq8JoXCIiz8mH2YIAjQ8yAMJ/3sebG+fjrjKM/2ABrrawljJt3quPLe
TeVbkBBvw+uul9NawL8MW7JFKsAfgMkInjng4yWyO5VFNtM5afYS1M7BgQcKMVf+Vdy3HoXQjjd8
hISXKlsFvClehahbJYdmbGlj9wQOUp/BpUReC4pA4A9++Blrkp1lwkR4XduRdl7iIlH1Tylc6kZz
d3hRcc3BOOd5UwW8HaT93hX3Yh2vBLQ6vwsMk8q5t7q0P5tHtYTpNJgiDq0y19Q+jAR4deDwkWt9
7BgWPD4qcnybYTpP5Th3x1MkDSdQoAeEgUeZBxgvgxdJkL9OfZhb5bCZLvWDiSA1pnAU+6qmaESs
Q72AMa/h48IwYzvU6/c6OppM8dm6HCEpaaQWXRSYn+kuoM4C6ud9yNF7ItnaDbdo892OtdQarkL1
ACllxtynDtea7bT1LNQrD9N4BG2KtvRrQVpsXumQE9cRcTw93FDJmujYxcXjUb244/d8g/SAJWCJ
lmR/T09bMiQPmqKk6NsDtZXofkC2rsnjHm7B0C2g1GzGdElmgFvoBXiF/p1CCTCtK6LUooQu7RFm
JyaEqfEevCOeKb8ejGTwr5X9jrmNyhGXH5WUG6TsIZyeqeZ5zbHKCDvPFK/xVyxpZTeG25h1Liuq
+BYFxg3Hd7cbTd6sT3VrlxTBDUv9rbSmh2EQblIAQK9XxNeppN0gDyUwiZgmOWb8guXMUi4FPa/W
YJt4CxO5KmamRwSkC9G1xLzodM5id9+kTVTc+GRVWxCooIqykTiO0CIvGhiMkKylJg/y95Y5el3z
0b1Zm9vIrnJnggyzkWyQt4tuQDwX1wS13dY1BfDWfHjskNIxGAfapWl01nSCzjjHb+R/b0rpWBvh
UxoLWVFqtkVQOIlLTiK/G8dMbz8l6iZAnBouCHCAw6eYhYYM4uc7tn5taIqWf/JOuNRi2UJ3fBXp
RqYJyzsSj/ZLLi96fFPKTXVyXw2Banhr/aMroseET1WH+k1MNpnK2OdLKiSJq2/Q73aJUoxJDxx0
rpOlva93yG7wqcpv1V6dkOrXHrS4cNZysLxolw/nsbsQO4kei12MF/AHtnO1cLc3mpPxwfDctIvE
s6rUCHgtdhW1BOiA7Zr0FwY0AezJJcSnKtk0CdO1h16TOWHNoGKu0khZYxA1PDtMjuLM59iIRR2J
24juxaw5VWexXjk1X02pLMU9MF0XtCXd+svBNboVRGVbicP4N9K4wXnbhDs+JHPHm9FLPo25kg7K
ivmtTC2tkn7LHm//HcKH/rKK9QXmIItRIVwOTasd1UV9iwJmGCGFMDA5flPpTk30rEP58UpcTDvu
VeUm/lQcOkjLPhh6Gefp3xbAC96UFt+7zTNKugngpRUdSSwoGPD7uXL1tItDybzKNSi5Ie0dJJqw
Jb7LDPfF0fjKroGGWbHX8b/Uze5bSHvLsbhbTTT8uYjYBCSgkcZWd4vGzdzOQx9gMo+ZbJq4YbJA
s7mnH0ovhe2dK4zYPt2qhjCfD/lJptCekXZHaD3pKTle2FO9BaBKPKx0jDhtwrgSfiR44CAWrp/e
Px2nssXIthX7Fg8d6WBCmuDeIVZi0HkVVM9o7B8ZEY11U9p4szE6MS++/ckwvpllEO91a9VhXulf
iAYLDZi0+nfz1ZRMLoiLp9srZEsaDAOE+0J0sdRBmZIjGbVzsnTCgptg52hYgCWAWiMyD4Ue8n5S
nQJCYTTttTZ8bN4xupE+r92I5tpMGpGuPM/U49BH9VyPB8o2g4WcvNspmNgJcQHLp83vGyDNjILa
iNpyqU8uPtxAdm2WYc9E9t32LVaiN0r8tlwOygCYFxULcxjo5moaSX9Gfkts9MkG22hAr78qQvtp
1NPRt7JkwNt02w3P+gJ90snuKmYAqCQ5Pz2WRlbpfmx9OIo21suHc1HHkW4XTMyQe1esrTn9EUDf
D5ZIucHBXYH0L3vp/6r+9CYi9YcfakAI/kktIhpXi3G3Q7ZiFYj/OtusjswAKAz8k11tFd99bX62
y6PLdOn5BGUzRejAGyv2h05KQzpgRz9y2Wf++/JwuPQaXIQ6Xfiw6qxCDVsqj59k5zvKTJMOhXXU
iwJ8MeAkqjRo8PajI2TnZBkv5A8TxFV3F16NkyzD8hrDqVS5maR2KsnNmDMa14W0L68kWrWdwBZ/
xLcW3GSR8hGiVcpUz2AFllGIt4jQFmC3yJnKRDCi8FmUtkuS8jydCLdne+x+3DxKb8fngPAqbdOu
6xlCGX+cl4nWxQU5yCSqh0GCXVhBelaQ4F3r7Wt0tkZ97e1dfkX+qsw8n+gSGLZWYUu4+ud2fOt4
3zApurfF7Ot+i1d3rD2ZAUtr4pb6j72AtT9oIDnE4cYYq8kD1HAww9iqiUf5XNpD3tIzR/5QYF2q
gqf4KTpOM6niPhV81JL9vwxkPEgRWVkZkOdiZDtLn7KZBELthjaCPpqs6HMp5LPzwrKp+ducATzR
yz1oEkOrHX2QVNt/PS+qlCTFKGw/h4hRgvEDN7nMWW1uHZ/hfXltne+NHhUoQeUEm85HG26VRmzk
5QW0XcuAWGEb4zF7MHhbFwMyO1BdIVT2FvC4nY+kMPFXjcesl4i1UucD/oEbe7lcE34YoX8sFVLT
FkpbMbJrckbcHEQyOcRpUxuM2z7l4M4zbNhC5ugRMyRasWl9SjSypiwCd+woh5dmMm8MojwougW2
SDIgVTV3gP9eyKS+2ZSqceyBku8jEbPmu7AqIQMnAsIEQq1qusbD5FRYn//wnVC5EINgRPBwmKMO
c78recWfEREpr6xjokb/5tyYe+Uqj5wkEkz3Xgi/SK4fFaIA+ELb+emFQHm+iNbdKjSN/RJXI8YO
seeomqfaldCU/67GpWIgK/MZfJqURFvKRL1KWvuDLKe0O3O0+cTE0vXqSAd1AKM+GEs8YOdi9DIy
qHDnbmp/2ppqAdU0T+j+l2iv2vWEnjj2Mb806DfwaTyv4QG4mqUepQImxHdnSxVDgwkNe4+PCF2T
0Ir72Nevt6HzSeOO8DUH31iAX8JbBwJb+4aLA4cWfkYG1z8yzjzi4arnuhwMkJqGzztiZCjC+ut0
kS6ad8wY80oKnimuH3YcVJ9DIooq/if21rkpG98pao2YhY+OgogmMAMfIRLAmLwYbYYBudH/igBb
hGBtiMqG0RTApyx92CDI6Xv/eKdm5IMLgxiqVwt+EVz80zroY08NfVEjbIcscm9wiIVpExnMPVzp
NZWhsOI1j1cm3hjW6PLshRZr5PbC64JLXp6VVVHTcnDnPqk2xRlom1kVrgtJwmuKYDyLXQNbxRNl
qltZU9hpA1Tu++krDiWVgr3EsfGaec3zXQR9cc4+h0gNdV8OxLUdn0nhdBuXGDSQk1k1nx3Y3pEq
/8hN6Xi+ClxCjMU1EJe8G7GEMEeCXZEYwoji5R0Ru9Cc+v/9RAGtQjCaW/PGP1Iyksc/VKjcpF/c
/pNrLQLOHH1zUj3p3G6XZaUMWPpiY/+2rIexHZ0/t+NYOVMVVARkXmit3BCTIBdugBFZhzEjSnbk
nRKXRM5qzU5o3jdUZi4K5OgxgKsfzgS5eO9wY248m2iq3l0xqiO2MlCIilaNyLLHq/UVAB4XHV1m
8uMi5aBVJCDRpccwo678bpwwidy3NXFhvn9AEyNMTJiC8qn6eXRav7bvbCmRpARMKlixHwpCwQgL
VF2bQVUXJEmf+jQUIWbAVeXAvgjql82YaPxSdqOXHu/qiv9e0TK+MUFqnQ/v9Dps55Z1jdAftFFt
GHBlsa/Rt6olrIQPdU639OOZj6HiHlNa1lafAP/IV107YEGHP0QFabXd9HV3G8ZohTHwDgmXd7ql
PxNut/J+vXIu4UTAEV7PPpJ93FLJ58QRPFnLnPgGwxSVQJiKuOGOspopGTWBrEREFO4rSCaY2Bno
dijbUwSWmkdoaRfS9xsKlL5fY274EHa6SrP0mYswvaSuOHBAi/lBKYsGw1BZTOg4VaPFPZO0MXPx
GU4qdh813g8SQ9UUGzRnaO5I4rIdpcx6jm2kaCiCrFai1MUAfRuN1qfWarXkvdxuzKjzm+esdyeR
n36i0BFFCgcyWBnVw2Ag9oHwo3SF1veR5l9TDKfLqTXInqEaH8HKz4d3SpodsJn75Gab0j25PulS
YeePekO8Mwn0jOod1PMqTmQcnbv8UOnAOR7A73z3iFxJIZ2HJ7zvTdn8Gfp6a+ESTCjuW2KUIET0
xkHMGPyoUQ2DEX9q0Fu0XDUIf7HfacR8nMqRQQQuxV481edz4Xv2OqgzEYzp1fWk64kTCd1sMe5h
EZCjpFHxVMFESe9Rdxaj3qUX5M46SV80e3TsUhCtFvnLX2VFmg32fnTGZt2J0e4TYSwQCuBZcHDq
FlQ1S1v1ETpqaL7Y3AL653SSGoLTkOtpVdLmnFwv028PY67DC4zGz1PEB3SMZzs0FI30tethkL8K
SKAmZm103VLvLmjyym9/+6ZdVelFAIi+rk0lt0g6A1EDxDc8n+Yy9ri0FZMFHcHf2qILf4MWSHTW
D+8xxUY23clv9ANSZUU8jH1qIwopkJi0Odup4LDsQmguKIBhZCGt0ma11b+xuMjeKx1l9uyxP8T0
cK3S0nGEEkvyR/bHSCmR1IlOMqkuu86V4KwKJDABr3J4OQ41mWUmhcypQ6W1YQIgJL8Wv/zVTTll
8+fUjhGDM0g3LQ22xhNz5Y4m1wCYUURMgbTXhnd+mQwKMGXXXRodd/vzSO8FYgh8cwA5KF3ac+RF
DP7CKoa52rjanZ6yLDzrk1Imgqjlc+R4j+uPaUeGmd6+ULyvzJ1d3y8poAq4lgTAzbhpKNZ3a4xQ
HxNe+HgdT6yjYGnm2/vQaYWQez/nIekMigdeiQSF0R09GUYyp+gTFELWXpIU4J/hpioRlC+D6sJs
LQR5knNZO+yc5uuBoSjCI/QU2vSd+otPBcuZcEzE5ZQd4zzy5p+gvq3lvS1tRnDV0AE9C8bZICf/
dOoY7QnUCryY2KOk8sUSuZjxgG1HdGM9h8NGM5fbIPbji/eodGaPtIhCgubsajKu7DaZdAlIDjsZ
r3NdQa+bAUOl0sfGMblJ9cubXY/mSwNzOJRirmV/TbuF0rPD+SGUdrwUknnBMycf6k7h38gYDX1d
m8AlbN1HlTVeHCOcSWjEpqaeA+9d4PY/zAQRewkNI29c8kTwqgWySF0vQYd0SZ4W27FaWP6bRE00
55HQT2BMyr/7xu2luyN6mC2aWh4oRqCpo988Ue5Uf+rFq8J6wpT1UaavZe2zq+A5c84V1l8AH8Kp
NVU7TJf7hIWO0naeAWU7RUHhVx8YFXYIiYq7dysGrTjgijntrSgeP3IrvAYkuEZgszW8JjmCI9OC
+jnF8+Q+1sUWiEQLdVzbpImrfqldMLjICmrlDxPqt4B3wK0eTHZlCQgw2Il0wkYpOlIoV0/dDYt2
tKV4vCNnW9/NpK6t6MeaUJBWy3qTuIzbrec6RaooCfmAYw6ZyPvIYxsVhPzOvtKP/abKqZOAHulP
ysf9FAiERjFdYTeysC3Em5m5XHVbUruC4XrirNwnSabip6FHlyNmECg/OT+5UpsvouTNI00neNqe
1+HetOAzGvoeUai9l71ZTk93p6TTIjp8KfSxqclLPHVTc+8rDG/3Bh9yKmYJ0WO67jLr7RClgKsJ
xANEXGAD4kUE0LCgKmiHz3gWuY/6yg9eD8T0i2U2jrVz7/AgT/57blUvGXlmcOajtzgFMD6L3vx+
a6YYR9bbtxurasdWDlg4KBt12VqCs8cfo5Ssc1YDqnrDfQ4dCn/K4dtbVhAlvT/16BPczLnKjnJG
DH/b8mWgJn3+5IvYZfOebxZKiTkk0ZD0iIk/hUpAbP/7oyeHUIINeegq3U3Z5Z0zCwQQw2yeTjLF
LxiKBmwu+1SaxoLF97b8WZ5ElZw48ff9MhlreoULC+J+rA/7fShpPxHePe3D8NgtMCNuHb7fvAz/
D6O7+5YgE+JNQbGo/z0TDBSPnH/Z7eJ2h2wf9d4V8KELPbanauHh58v6b0/deMqv8zrErEip3GJ4
NPVFk9X+NYzLYyWY5WOt3/Ev4FkvsA50XTYemCUiHfLxIWPLEXuZsYMKL3IPkOgiuo/3gA2bJjM0
d9g/lnfXJNEpDEWqMB8p1E94W8Xd3Vx2FJWZZ2suExwgGRyMbmB0zkpCVSpRUv6IwNqz5wqvs62G
0AcFnM3CTnTpTkeAUrArf3rzYsjxzQlK14OL/HoTCNDopZ1D0790Ee46HfZ4gtFYZme7C7+yN/EK
XXPMzGv7N4cR4mc01mIKcg5g4z6R/FS6Af0pd8Es9W7p38r09h/lGDOPs1KiqmzFtgHH/99twLKz
69vPJwsSD9F6VKzYcYASyJ1Ncf1pB0nc7LuirK5mPP094/rw7gcPFi9D5tmMAGIWycBLDui3oSwK
uTQrIDfskF+UOlyoclu7kHsy4fnCKEZgAofGfxouTSTTnWU7fDe/QMpKu7me+4mEWbrCafDUp8FS
OdXs6fXuJtNQnEVQCL8ZOH2aUcp2T4u6KTkTa4BX3wLjzKhtbxKtbLRVlmehzvvjE/LAsPpyZpPi
wnyK3jhqIWa6pGydax1LZ0j2wWU2gOQJQkNab6Q34PIUSYK/eGEEhTWqqhdis8lhDCVZl5+fRvfP
QOzftAWHvrQ/Um+KIUOBWndBs5lpknwfrL7vVf0sZe1lbhtcW8wghxMXP4ip+ebA4TDyH3HfNIeq
ck9eMlId1QcM/v1DDzPqnhQFQzrwy+N1fNi60dJmKgwBD5L4aGZtLmLe94OXRMVJz+BVr3qqKJx1
WLqX6tF4JYtMffwlHGXwcegaOPhFzUrNpxWWnDaWnc6EJzak6if9EehzC61unRZ0N8zdaDEVtfAn
mpEPZpfgga0n0hyHkHV+vJX49iwtciTVUCOCdnWqU+n9cwsu8ptSnMXai407ycbnL8fLnY6qH2Y2
gU+8Sq4nCuxt/38M9G/x/fX8ijYWpziJUfRUmnSqHYB+rsPjEov6MzHloIY4S2hDHrkqKy/YGZL0
WqmBsUW9vyBnNlKAypOYKgPG2Nke/EXnyvX+yla7AdBTVwydJBJ+n5iXzUAtQPCa2DtDlzH17Keg
S2SZBwQSmY9zh59NdQ7pFSp4g748bkv1VA4pU9u0jbdjojr4F/jIrGl98iH9yJt5ABppO/beHn7J
+A8PrtflOAsq+3Or5mkCpHvsOMT5NgHkazLGZtoXbzDiVDeSlJSsPlpGTKip2eAt9paGCCuRRcZi
WGkJB2iNxR9muKayrvuLR6F//syRemJLnflfogDHXNDlcZ5vcQaLMsNT3WfNykFrnupOAopwPwNy
zKzVwNSwGwXNjaxxcKAsRrs3c1pZnJ3rXCGp1EXMdxAtlPPkLTAQyP8xWfussMT55oGM/O0nUUmq
7UPNDYGaIwoF7q24yFrNG+aaw3Gr/Te+nEUmTof2FEzJJjfcyCtgs0GWAu/E8t4g+H1GcbKET18e
mjtsxAqf/libVbJt02GftI4LlCVOfWUH9ZV5cHXIA3V2MXCKSVap75ZaGh0UIqjbX3zlnBDGJZ1m
hlWxs9s4f4m/BNZMbnKyUwu5nuD4EDtYWcIG0zQo1lMwLKPkO68/3K6+TntH8XpVVAEruhFQT1Dk
5mkYiKtM87JMCP4ckCS7r7kFyysBhjLt7lDo/qlL0bTNUrTvVnWUsCiYwIeFSgPZ4f0yoc7G/KEH
pmjwiyrXoRdXd2isOg94Syr7b8ij9j/9S2oSSM5LeSSoM4SRcwbfdXqPn350ebw4il901Kehhfmq
/1CyVrs0As43apFvCiCtChVP24K4bJ53O768tCkopZGOA5qFLhbbsGt1lsr8IlYpml1xO9vgqHtw
yENg/0PV5D7kXosv80q6IYwZiRlUq3xQ71iM5COmbYtlW3HI/z6emdHW7tyBe/PFz6sQbutf39cr
OkDuTtdZI2WNa6I2WtqwQ44lO3hYLPdxYhMyYIvTNURpDMwnsK7Jdjd6mPnwr9DfUl5V6drW8YfB
qmDfrHKBOk/V+bSunPzTy9xQZnpu8qB1O7pr+5rqbYV9Jl5JuF1FicHh88UpDo1NXWny8gde49bp
1XwENCie+03a8GNxzLu6TwALSBgChYsSEg6zMaMXXh2PGyBYMsrkTJd4KwjIDTZWWwh4j6WeD0g/
WokxAeOCxMXc+kdoGZJWLpYa3b4D453bXlGgnYcHIPImuPkIRs60XhmNy5Df1X4FNgSJ8Gapvh4R
oAySJtUa7goEV09cEYg1EeFS/JvqH+7Ssknm9sA0EWr76QSorDpOOGj47gUUHAqTmZ0u+Qi4lCZj
OsGY0coLGC8oazSnT40RUhdsEojDfBvtlbIMYVsexbZWTJb3jRXEYmoVXJBNZCQVpUKYm0mzz/Z/
s7FIQW5ofFYhDH5Zta/o5CTSKA3dSgwMOXbioMRNqBV/m+yCW/C2ShIjHimLq3Ud/TQ1uIn7zQ8j
YAJVnP0S11MZrVLutYKNkQqlmDZN9PwGx0gaNb2Ru8BI1bzx9tSOZnjZc+GqFm/y0Obn3ZDleJnh
GMvAaw4BboerHKAToU29h43iHQxNRQT5Yj3vm/+VF3S5hK1ryKvDktFtM6q4ePuFcoj5d3ah1YLJ
gAe/V6GKQAvOna+0hoxK2IkxVWEVtq4V+Vf1358B7VmQyP0VnhbEKbH7upPDnKPvjMqbWlXANzQY
nx4MbfKznqtaQWmER34qf2j6824TeJns2JPbbElTxI82xeTCn0hna/SmBJKRDQqlUJJdnGsnJB26
xmUWQcZ8+OzHDH1CDowvZRUXNrnr/bFswUg2UrXGbdQ2hF9K4b7saUJntPxPyOa+OzNMvb2YYPev
0RTh2HjEI73jCdrw9fKyXSueXYpASyMC4ipThQ8hZ3TMviVCC6VXkGe3U9cpOxBXNIIVJstSAhxP
wPp/mT3JOMOKeR0pkt0QLR0zqhu1lIx/WOeusnV0G0W0+jp54gksASg78gEVlloOiEwi3vSC1Gc9
dJyvEaqAR4Id0u8jZtFq5dKypY4r1fDCj7EHODCP3WuZsXP0ER7YoDq0gLnnhd5sn0jTsuwjSP+7
3hSJKu9DqEjG2WeNVYlMw/hXwRSYUMdgaveR8I7c4N6XGkkhekhNLOKw6drF5NvLmHRUJp7Vl73k
YKtRloGEobYS0MKpqOXmLNK7i9Ijd8XiPrTmHCcucU6AYD80vvaCU76J49u7vJFcwCaJsPXwRNDp
mX6j1s9lTNRv7yckj9qUqlL3jGQpt0GmBUJ4v1RF6xu0zdTSQBkv/LHJ90dCHPY7/U1oeXpOGbqI
ruwFq/ubcIkMwIVpIuSaUf8gUrKFP5mtnPeo76IjEGRVpB2KLRdHltJg/YzFwYcsejkx0r8GhVER
XvOZXRHMk4dcc0nlu6V/bN2yhP7GFUnMD5D6vdBzcibAHh4OQHwobtIQDzUW8PhPNRadH74vaLk2
BbqKxtCK/ZHHB24vy6HhVg1KT7aE6jL/lNURTZvSsXlY6HUFEe8dxDfPhgz2suzIfj4efvWHVlk3
VMJRiXyAVbf7I1E3fvXBeQYs7u/DjTKyJz13IZmXMTndc5ZYWM4iGrUXkQJTD4TnDeOPYuevwwHy
2mRRMRgCDS/qqLemzmMyYvTl4F92WdAVQAqfD5MHlc7T6a/Rz7Bg9PHPeouyS+0r2801KM/OzlQ2
sSjtf2d0sSNujA0cGCxf5QnVJ1WcNtE/ZiI2SfZbOuuXM9qxmI1kkYyg0vayLT5uEgwYZix8du3a
tD6t+1kszbk+A4YqcyGO5KfmW1J/IcUcH+teWlrM1X4Oh92Eu2zR1+SarA+VY1D4ax/YER4sAlXL
X2f1zx23aC65XazSJ5/M0ge8VfG0DDzskIzcP8M9FBwBYFE99OW/xrOQpHf6knYLhkvh0nWkd6zW
pT+WTwRYP/0SCY9MGyR/1KKrU6b0rpbpiqUdbs9R9166Kq9/Ut7casdmdBkdPM4hACoRg5cRLDGg
sfa1fbpWyEk2tsaMKiYybtjpsYk5V7Jk5krXxAvk18Iqto1wS9zvl5ULKAAkbgBj26JmHjC8LZYn
pEHxdzyJSX5j6FoB92SwIQUiiyx92Zsiah3qsORmbVHOxfgfr9xQtFAzqmIL303or9hEAgvb5oq3
gx2FM1mxl9iZygPeevxm7dAGAk0i95PMSWSysSbAFBCYiWJCu+UKcD7oIDh+7PWQelcqB3+PdZGk
rxivAyjCtsbrKb/Y21xHPmZkSJ4VTEKPmYomL/qlA1gUoPoovDo6qs8TZHIneyP1K0szWtQ2Xpmm
pTIN2HyL0llyG5xf2CH3ByK5Y7kYh53gUI+002ZmmEf/GXzogtMEh688NrE/7Gh8aOLR5+u2mESU
PU1nVkYStEhyPVaHDwecF7xr5VvBm0XRKbbfdNq8ZDuOSZWxj8b5XT+cLraJcFDrHxfviLqIyPTn
lj3o0uBPWK4B2vvHutQylCg3cW/0hzVSRxYdeQ0wCwavufh22FO9c/pdAtma/XDX5Oc+AVD6wA+W
0yaR3dld9jVpB3umk46Ijd80jclMS5wbTrv1ui8I/bN6Vfg5jTofpzW77gY3A7jtdCwXO5Ei9L/u
bH2iPPKlmBVgH1QcuSlEz/Z4GkegQ1HwX5TS30ErO1VGeK7nnJNYMsgL+DKbwRDCQ1+RGqEiZ87c
JugGtNISf+iXLOePreDqUJ2vPhLFwHxQfF/1LJcV94q2FW8UrBOmpxy5rr18q/F5clMSJqcljksk
6/jGjuIprapWIZySjmy6f+DuBWdOv1ABb8jCDPiW/IL5/WeV3lJ1Vt7Ixy+toSLzo65M9QmodMJW
3u9HH4Kcy3JAU1sS/Gv9iq7M6AqnjH51eQYd5c6VO4v3Mdfn0C0MOksmFtgW76pU8S42Y9V5ZDxs
tJ9J3GjunCZG3uakuwJALjFPKZVm/IwciRN4RgTGqxc+pg5CCOsj+uTF+dY+i2N9ZBvo4X4UDib3
M7fBtHhxRnj5ThrubsA1SUQxjzYvwO8B++0Ccf1IGBNvgfk3PUemnID5232MumJO3PlYa8F2oAXQ
vN7UiQJIFstVvcv5JNJgSOGqH++d8QY9ZHseoqSCEeIVJNPa/7Jl8VMeCJkLIpLwAHRPRa3DtSTV
WzQhMcPZcyOgo33Ta43pxIlo50CTWgimT14FT8D52PCi85I8/KT8+pZ2k57O/+dehEkwTVqHAJmD
k5dJYM2ZTjfj/N7Y3he+rkmnDEB4R7c/OC7p+HBEPLpHgOueZs42DXNiInh81l9FcO/IANNw+p5W
8qiPgYQhP0hzG9fH1pTVq7h6N2CT3KLl0iJ4K9nUoLVs5sQ7pazpovsxfH07i7aZpajkuwvn7oSH
sUDEX+FKhWz2J5PMO98Pykxid8PBl1GidcS44rJZ91sceLi8Sl2WeGG/kLre/3usNk0Jr/geyCPb
T35nPGdlSW5M1ZxCltLCsD1F0scZ8bMHL94q9wyMNnKzWL9AoRypNZ7aG0WKrIq4b0IpqC2kGNGT
OFe0TQm3yaJOrOvzyX+NI+R8ptgDPIuTThmXsAW1MkXw7c2mHRfjVbd1GgLwGsOY8Q3Q3dbDXbdc
qfSvRki41yS9A3YIKhwZf6MZEIG+d7h4quW4hRBApJwo+xmUcCC6jZCesBWOxz1u++NPlgHTYFyz
wuGG9CdQm1SYCyeiSdJfX5Am0OgjymzDWJhl4Z33YsB2uRJC7NncxFjg3vTf7KXGzj2WHowwNI0e
yshsGZYZpTQvH5tAb7S9w1aHK46rXHapxQxe7GcOfBfgV0IkpNNMn3ag3A26QMgn9B18ZAhG1qn0
4EfV5h3Kg4cIZEyWBkBaKB7NJNwLFaspQPmstoCVBF9SUqOlBP9ODrcr7zJ/rsZJIZRRb7WZpfkh
RPXsWjYB8cmNb4O6JW9F0B1757laogftlFsmVnUUY1FNwx4sLKeDtn3S2Z6aIHQHR/58iMjcTlIx
6tVlICbOKAcbvOGrIiKpwnBq0KuSLT34JExQK/l/DIHoCMK9QzoFdBy0puul9OgKvSA6kkpcG1vD
q2sL1FOWwRivzk2gZqyldrCw3VU9Xj1PVvrt/5SmFWxUma1vkfWNoFZ9dZ2QrhI0wSXsX5rmdBa1
PJsYyViT/6ReF9B2I5iMEJm/jnIuc0qoNrb6HheeeykV7hAK4xRfSGKUeIFgwoOhpi0+uT1ehDib
1vrQoArrfapJopVngBFW8TiQHe0LwxM/eaMy2kqX4UwYgmdBVgsv43h3lu/LtPuKvmpguK9mJVnQ
We/QH7QYlvjcIomPf8MMwugZ2p6SYErMOKn0tKMtozPDF6YteXx7dzJYNt23UsHZ3nSDGGU7awDX
9IHIz4KFCKG2AhP6m1ZtigiUnBNZ9Xk5+3P8jqnsj2w242zmTCQa6yeH5IJQKQ7wL9Nj753llh2m
uSSjXK/r6KtUyKY1FVZcaGiRZOimyzs26jxlvB8zjNUq38lqQFib7Gt+HKMbckN4RG86cUiUrlHG
tkFkM5DDsqJ/XqN8sBoubWwXrsALqMaTeDTy6cnklGNr1aWroUSRv6vBizkKHTlmjWATI3Syed3z
aUg21x7b4x2C/iYkGvCHjl+KeV5k0cry/UR/z5vkbnDgWf4WSH9iBOnbsqv4ceVuUYborAGaoD5m
QoJOUa0tO507WvxA7GzZvrdTUTayPIU/8UIUUw+XE96Uc1ZIVZxMuZBecPdeAdmLwxc7C0CrhVOg
mGFIJwVUimKUJTwUyPw1kIX7dk1A64TokmQTQllGztMuCWsOrwWjFyxMmnZwOCG86cr1V/qejlbK
jj6n7R8Tgi5uEvNTVpgd9RClVIHBB+Qf94JCIrRmNh15tmZizPGSu63tF7n8INzDq/iEhWsgkHfL
Ycmt3P/26C+6mLsHh3775uPc0v0u4VKZlohq9syV7zpQSLa/E9CtWFltJ0kuKJYhrWIEx/CC07Kf
NizQiw2nuugjVdohS5BAXS8C28tfAZvcSwQ+uBzEcTdHWdl/INWWrEX+Pw/8/XALtcdp6DXggXcG
uaLK1W18jnYB46KOjHQHYitt90LzBBWaoKbLRoLr26G0YBQ5KkQXRy8qPlQnW18HQ3Np2K4NriWQ
P96Tj19wGgoQ/flTTxNlOkNHCXX5UgQMYPUOy4/+v/o7vjAo35+wc4NIveQuD9eOUhW3Xzzu3d8r
mRoWAysEuJqq/r28Pb/nkmu9Fu4eQmpHvZ7b5c72SUWZX3DCC2OEno6lZfoJdUvQEkuwry27R8yB
Bn2yeLuBdidAByQhEYVItT8fFx0NjFQF9zI3fEvTamkjpqbtbvPfP6lVooDg1hTO0F0jVC8w03aX
WiIhEGIQTlUSmTkfXN78IyKXuFPsd7db/jfEWzXIlpEhXFTh91O0JBEpcIu05/orrlY3chvNREZh
8UujZsa3nEsB6U1guBJsYNd/XWTA2bx9QpOmtP00xHsis5erxMhS1AqjPPIpqp4ba0xnjs8xhiVO
efCDUcbANtNNRV4zNgcU2kV7T/6NEKLUufDB29N8XjLhuXJBgL86kZKJTXKSBVdOIE2Qr9AXhFjc
HtkcRNxMdfEPJMDgBTUIh6qq3J98xsgCn6+gPDnB1e5IfI2yDfHbDHW5HBSh4lzwBbnx5IjmEaoB
YMIFddfupAOmsK/Ko/ZC+lVXaokP0umL+n3BiLcAEQnbGwQdmy+keocIpVtkEX64t7TNQHRQzK99
Py5OjMe4ZfNBvHtKFAeofIgJBVLpKjCEx3IIK1VyZfUc9+TnvoeVRC8noqnr8MWihoMdmDgRi08J
Bm+iFX4Q3/sRv4C13mY95/H0EbfGxkKI5AsaDU2NzvlObtu6BXcvbA6ak7A/q2vY3RUv73/gE/CH
4mcepFRKXjy+5QX+bDOQKVFKvAIKuaxKF1JE82IIPleFi9oGwaj02J7ao9kXnfpg1bnjPF/JJsl3
4S5g4vJo9yLDOItPXmNKh5RRlQ9zR+zFQFYIZv6vJkHYOf0ikeuqtn9O+R3moIuGeVx6vJjOUc+8
87Cztk+2J/1KvxKI9kd1180dijRefwmPekLnNGPfYbpt7etUg+3KbApn6Ob9L8H38rFgN0xdoSu7
f1U24dBIYKn/gW2TOJBEQvR0wsxuH3sob4CwFzR4n95SzvWicYmHBrPBeCRgDGai6kW3RTZBXkzx
/r396v4MsjNYabZOGJbn2vVj1pZ06Q6MPDiKAQ/OI1E12Mvlo5NFmi2sYAeCvF1wPOvAr2NrtkBy
IDhHbFj6aD6Ttk4XyY7wba1Cgb8VOpO0yNN7y6MhInFD240JnjA2wtjtsh+q8WhVXyo5eQmey/Xn
Uf5rf9k0zzPb5IpkuQvAegOcnyn0m2adjDOaP0fgLZ7DLutzH8dteHFHLhxfoK/EazYOWlFSmpIN
zJfDFQ+M6XNZ9owKtzBAkPTX1HQrkmQeDPuoL4ci22OOckMUc1a4t7HUI/VFVczXqTbm7fAKOAXF
y30uDkSbDP1s8zoQmLzNAyL0VbqQ6jcIsIHx1UFrB1B90SWWDXUegPQdi6hpvKgOxDunGc7/C7fb
Fowku+YjrvS7j+7/sH6CnxfHsjBdDJVtnwZTFb2EU3lKSol0gT/G+qkgr/s5CZganaG9WxSiGfJC
h0Vo3Lk4Bf3ZrQlWJ26r5shsbQ+kdS3gdsu1Uue73AxfVdSupRuRQo9uzOlZHeLqZSzPLRdC1eo1
wbhvSGgxqp7qvwHkT3jrmYz/4LJZxDN9lcI2a912bYt+j/z01dRX7E4KGfU4ul5SuGj9cq+mJCM2
uemnDZhy3UfyZvFW6ZNIshIbhhRyRdDjtxmIkHJPWJ0Himzs5f4kkwYxfLGTR34pGRf+PJ14FnQm
QJZisrATOI0yB4T60jd2pJnnB+CnA7WsmIkpi1aJcBbheQueWsWh3GHOQsHJNwhiUFGBHKoQAcbq
6RJ+7Npt129nrkepVJhwz7YVDXNnBq8cFFq0/HZI3fA1PfOwf5UAYoLn9bVoPetiCysPLByaRn/A
cnE4uP/HyFmALT8LPR/93NGjii+HetuOayr4eI8YOyrXATMkOXTfi3OZ6tpWYLiT9OnPQFLmOi/p
X2TWkhysQfqmwNrhaRYmS2bSeHPxOvBNgRwJGfwoS+3thCtB7e138vIbU3SQpj0Ww0TsY3oR+F+5
v1z4EIOYMPsleKBZm8/3SDrF4oQwuZKzLesU2mNgVcXa+/uZHYpMFCYbNI/qluHD6s6Ukaom/EF5
v5O2upjMx1m7rQYJyM7rVfG/ZoAag8V6X6pXaYBRt1Xk/g6lBU0LT0nI8fqPgq/eN+sRWD+3qNnx
U3J9BzOIXMnn61LCVd3Y9yRSp13tXRaKLtrP/nsLWS+dlR/4lVu+4qqqt6JcT7A/HmavxWoP5rBO
QvxlGx8UymBYuIn/5cMFMEDloaxd0EWaszw8uYnCiUqj8vZwGrfcxPnDqUt1lJmm/YyIEgftUeSh
mZw1K1506pdnXKy7qCu56v97tAd6+Kt1vLLdm+aZHknFjPTL8VzoG27lOX0athrrZ6TFP4kFHER8
V1TBcnS2ixwROXzYOJuJ5meiGXCHCNqb+Ox0qyq6/FTeXeFcx5vGsHY1XQowmxkWJt9fjdNB3Eaj
WskPAr4xuOnF8j1eAcbGapbjwaqL+fjwZuxb5wNhqyVQkJHVw/0fwqJjBk773DEeN8BI0stJ2wLg
3KC9IQALHdzrF/GbvW3XY3h1dWNzvZV86fldy1oNl7QN5/fDXw/9nI5fkGqOX2Js84pgo7hyhNHa
DIyF8XFxhNRHJj+yO3xzwG7vxjjganW1++Pb1ysxjMjtSFLPM6Q7bhgsaugUSTVkOXtLePo8gxfs
4iI/jBD62Hjs66el2phDmDftud5pj43tDEFLePwnz5jaidt2FbWTtBDZvY99o41mZbPv3owcKCBj
/GNz8fMLnwe/VKuFazJsxFDRnh53Fx5R4gXfX7qhAItj+9xcyA1Xt1GLvZj9hoscNGTbu+5iiybu
tf0N0VeYy99aSFebodG1+i0KrM3zoOSCv6K2zjtLufy51NmZoIHlUJwaldFUbGrinZSVgXlgz5rM
gkndB4mr41W4Ean9QtYyqPaH6VTIS5TwfmqW1XKY9bC1dXnSWzHoIx6kGmfcznvthtITAGAS5K0N
3IwlANBVbGtBNuVnLZij2AfilCSVTPEXGnkzMBuY6jZSe5iaACWTBsFtKe1+BE+W2532TTCFtMSV
271C7Gtsx5ocat+OjAlvJ6Y17xdXaOZp5JPZ5cN+JnMwB4dapXaV9JfbSp6JiwCtJ9nJi9k/HMBb
WemzWmKea+IBjheMKXVsebehd8an6hxXUhDFykDouqx6hSHHKjTCMfdHf7Eag32PyD0L6XYP3xwT
hgeoNFiBWU1TMeIiIHsvJV+Xz4uIpRbY//I4CTIeEtQELLvr5jlB2zs8n/2EyPt3k4qcotuCtj7S
v35guLQwYvIE1LZeTpXGVkkWVtGJX60ZSsX8RmxMEAOL727KoqhhYLUbLs6je7XWk/nV0okrdqwE
VKy5DmlH8mQNkMbKa0TVmVrp53WQHXaKoi55QaLwQF+lGk4MTU9GD3lpY3rzYgCJzCcv+eg77Ahi
iEyWtCJ932+AFn2EUOWdP5J79G9CRcV7478i4dVWiGqkE9RokL3NWSRMkSLJ70dI+dEbsdD84j5e
EGmcRXYZykx7ieIi11W4v7rR/io/hSKEfShqB3Krk4vxUCDMM/5+iVxyTkV97LOWgKo0KhnUM/d4
8AISKzM+WOTVjnqAlMAy8kDbDV5xw6ShN4qooh1Qe+I3dloIn8gJKVlKS6xjdKQopt51tU32zYz5
pRlM7tBYNxqUuEtFcJEwgyS3eRVZQP9icV5oK8NRe61u7o5ZDjQ0TO3r8tj8FP38+yOsLFqKqbDT
Htw64X73dedIQVrLKzisxeuQdLDKDP3wCF+f0hK2FQ5JeJRgh7nl+v3BDJVRZH6jClFzdK2bbmYr
7pMyM4v8JqdicXIb3iZIaLf7NS/h+AZVfjczGg7Gd7kyjOkx57jFZ0U6b36bwRKUNX7VVZsQl4j3
/LeqkB/7XgTJesQyyYgxg7R8LAuyAe5WXxpEj3V1vPqk/7ShzsGeVYpsEYIjYGyOBlFYr396yEFD
l44L41IbrVXMKWa4P7VAvNtq2IBEZAnJgOAB5u629L+IGgSn9fZdud1AQ6QirRvueYi6FmCVnTMw
kYX6918T6+Yvl0jhAXr3G0BDp29J7HC7so/6daOoRovN6wiZIeIQZjW/7yYEhlr2L4Ng/+7Aqp0r
r3e7I6kvU2ciwYqApVzSHalWUPp+ryPNWOKk1T3ChEw/B4s4tS1ctCXn/DKcwAn8Qx2Tmtze6FAz
qwYSB670j9ujZXL/MT0cuiRM+Ffr2n/lvougfoYMz2xkQzhUXw48UYPudSPNuA82l9ETSe+Ynp4p
RqVybGgQFYVmbtA/dWcue12K8tucWZRfM2ireVF4Dlsh62pzjyugO4TUyztuIkcVbla3k5KMKfho
b3+t3j3X/oOoBI7/IJ2YoFFRezT3ZCHkru2RRcKpq0IPUbUMf/pfKowBSF8qEc3zJhtFwqJ9hzwc
ETCvHIwKiVaqGxsqGeMANx1OSnT6ayICRtULRpz3LcOCne5f8ZJ5ZKxnLTW7pP++sEK4+x5J/WjX
kEYx3NV/TL64DBp2o9InJoe0/nBKwtGUsWv51ljycaAJiSYUvSkhoMffwOatZgLpG1oGXH85pLqT
dtHEA7+ZDcb0T9hprokeQWQjRV8+EzFyR7U0vq92JC0veXP52rZ/AepyP9IBl5x6wGoeUxV8hvt5
V1IUllksVM0Ql+9saCUN2ZnBc7r/tZjZG7sW47M/NJrJCJG8yDuHPCnNC5ne81I4/0c1Z0kMmMBJ
aKLSK9QJ7pRquwBrvFab3ZXhQs5TkcoZegAKhkv345ICdEZ/ZlCUy054nPGVVktIHFBzRfY8+Pk4
p24TWgZke0cYb7NwIoQv+8L89/52wXxj51ODct/VZlenNAiyuzpiMZrJfHIczNQRej0GwbiLI9l/
ABYT6TYMj7uuLBf85bujnVCaPndG9uDT0G03HMVXTvePNhvS65ZagE06z08lvdknTjkoNv3rOf1C
CYAIgIusTnK3xtfWam8zG3xI7BmZjd3VQdlkqCSmwBg/56T+HnR3peqKT/mvm0mjZoLYnxd+e3C5
RMk4s6hpgnxZC4URGeOuGrYAgNLhqrLBVftdsUpudGww66PpCrDLDISLKhPMaQtPW3K9HBdBVwsX
BqFvKXaf50dto4NPuCq52DqQNJ3FBJDOqB8L4Wj1+LVyDmz2QPuC2VmYMuG0TmXQtTz+RJ21RS6B
X3/bY1h4/DYrwMkMpSX0BQlAcXkQSap2Y2CYW8aNPK9j0AB7b/AObFLUzIkC1CW9M7jj4rRfnapF
KQg1VYbn//1MM8VytnohSo2yVDv+GueRqIoEHcG9AMu0l/OIe+L9sJ2CSTcwgyUrQdZahX9F+0Gy
FVvW5dBOIpOyNFpDbzpNnODcua/YfiKTGBrRteKDvoits6p+o+zEJTa0/275zyBBcPIFzjPdGBS/
b37CPoA2yhe1Ap/rmUVYEMYDnfukC0G27lSZyEgxhCos6Kq4h4Ih76/qZj48L3hvQi/lZrN0VY1H
Bo/Gl9b0nXhs+c6kFmL/WZ8Fk895JZF5drYeD2W/a8ASSZfliNDerfh8ywelkVcuLX0Vq1PHiu3C
1X/nWdKVLCfctp22Wow1DOdA8EMtFWhfrS1etdHOGOgnTA/C/hNAN7Nvq0AyIKfoRds8wu1qMesT
8zrQMTlchc0bOL0hE1cl1i9zBEkxQ9+jF3/DinuqAdzStDa+wP3rNHjbKBouLu5MNRdi4iwKNyQz
u6U6BHsOuL+XHpzkt2vi2EsDMg7Vsm6HIojWqBTGX4QpmTaQmF/quISMjenCnheRHCaa8SO8sWSN
GHznWHTCfa2PrWsJDcvkaEl/tE/l081jU8t/6H1So3gj4sWwT5KwJnIVPKqgPyQ/rX4dm4YNJ7U0
IOxMzDiK+PTkBzDXkyjz0jYSbirLWkO7iTcgJgVBIbTEwuSwdWzTWdMvB8ZPLvhhVgVKFZuxAb5Q
1bq09JVjbm971QE/H37+sKjcxYQIlxUrnz4LwNjGqQnQ90u8zwdwC+E8RPUcEG1FCaPEmou+/bFS
gUQ81WuwQL+j/UyIGovtGVZ0OeCNFCUoaC2RylnAw6jQxA8NSrAn4a2EdIcf0K1Ere0VSx7j+lOJ
xwBsgeBXMSEq8OHgVOFheAh8qOgMl5g6xBfrd4eoywVSAJnVgJW0epEy4RUzaUgRSfLWOZtFslPX
5aR2b1FqjVdMY+y7fTEBr6wB3X0fzhXsTsvsiY3lNHNtZiGB3uzn1+95Oj62NWEiXWP+h9ee6UcQ
fEVmcSY0hV8GRgHfbz5IxHzjsnqhQjYEnVOsinU91a6g4powjQ87qqgu4DEeiOnt8M85TiuLLQfx
7BzBm3c/pvJDv5LMKBUSxnNvOjwPd2H9wW4uwmMafzibtozFEshLTdz8NNgW7jvykQpqksTy58c4
EyF6xVMdF21h4NHWZY+Yxv87pp99uyQbKKloKBZF3xETd87aCBglAUCnoECxuIO5ZO0PqdUihpMr
LoRMyaGbjgogsVfBInJ0ZEZPwQJRKxzxJyMuNFid4axT1GwPGCmgYO8+fUgprz/t08FYDgAQIxpp
JGqaXih6rhB93fktgKrfU6afpZTRwQWX+X106bI0JJWlXAC45YDLFtUALMack3izS3WVLGrAn312
za9Hvmfoz/qc44/neDrU4BESeNcRIn6xnfyJFRnTvvIcuYhCbv2caOUp6Cc2SzCyxMPp144BM3h0
/pUAfOwTx3CBceOLs/ppW9Re+DGUCwaSL6lmGhZRfjWIyaB4LGfJsjQBirxuva+TogMIdPy0lwvX
JBn+ImHC9gRKJZ6SZW4QyeetXkNjngM6LvzD2HKNshdrtdqlqEnGrGUDZACGNCV0vBwqCwX9Y/mr
oL5RtrwGk11T6dULIm1c+a6TjIBl5nJ90Kd2yjcQ0L2DZv1AVeqntLb2AHzk2pYeJB5fq/IlWFOV
UhPHgGxAKVzlK5ZMpDZJ16ge0cgaWbzCdcONcumLcsI/CbAp5ZWdtm/hMwhQvPG+vRSUHPh31b9v
3J/ykJGeiJEn/GNmTACippTZE/rDaJ496gqEO+qC5cf0PnG3C6NKHgmAqPt12FmWbo7KCs53NZxW
9qTXvgBuMYvq796gjBIYElSBVWzv9xhsoto32F5nKwxwzAyZ9BPP+fXbhmjBpDSphG/UIrE2RKTA
U7JKUrADdg2g32wb60uX+wunRreH4vuN8JbGhuMRDKL1ZTvDjDCgc2JSa2+mw3AR9yrigg8VyL+o
2gl7Wvyt0S4VsmIFSWL/otIxSkjA3qT/+wy+yTL/iTVtxf8DkiRw/30xEbA3ttvpyEd9MD6k32Ym
wf4hyBpYXgyMmmFzZPsie+/Y6BuR6bPtCFCVfEpSnp6bjM2fYZVNnpfg+bk5i4huDkAGjZ/GNZ8m
lkdJ7UmqqZimR11BBTO7zK+1F1N+VFf/xrsx/z5s82KzoYUS66CiPhw0J/xz23AsAwFkyQFWqEII
EljHChyV3Z7zV3s3W5EpLVX+Hz0m+mNMbM+/uRlYGwQ8RiqBM1k7hvc+wGVGFXEE8L8BTJwRIEGL
m1CPzMAdgKtIy4QZdv1fe9L1KPCGkwT1hfT54HYJuURemcpmJpETb4TJ56t9OCmD9THxrQ9hMl1R
CGc7WUdPXBZ6g7tzR6gHOpKcpqoI0qQ4hpedmvGo0PcpuctDASU5TMq76t7iVkobuaP+wLFsOFhe
XMheGXmsiAF5qa0NRGcD/EY5c1+JtxISa4dVorj6pJIalGLCRJVqtW3IC063Lg+dd7sets18NNjr
QuBX5l88h5lWLUj7+LTbYnANjauaR/XRoBBmMLxwzZi1jSdJyx59OFIhtXz8UisSrlE5L2LjtGb9
JTS1Y/TZYArl5L2dly4fY9NOwrIcM/3J1KM3j7cYUbxXr6/kI+Lg9Zcws4qjjUEIt0DjKfYg8v1/
9AdtAweur2adggQ+SeQ1X73s0yzrTkrTGFRSOGDItxzk8oCcOQK+xA7HKjAFLvyQvf8nyQwCMzyd
uv1IvBr4Uio73iCSrGsGFFYpAgYj5AA3YqDtzXo94Wne/LlaM4hIOZPoUV/fkqk7zB6Ap5lbNVYz
HuazPjx1czHvKw9I/jA8744DIKCsNNtbUc/OTq1+b45q6ygb6G36Wf+RrEUroWyj2JTgzknh/PDk
cDhTYMIwGSkIJGyJqdZ6L1gbhzl5JlqXtxPZQylu3zxfPEQ993nsPeO4pjx/rnBVt6tljQJ08G2A
rDFyzsUSCkW+X7BjymWxoVbOVzqDejdzCN5c+7YrhGaCmBhiVZwQZ0Kxjpghk1+zoLlReetMKS4Z
THD61DTBNnVqPoqhw6BttcRbpXMGkGZiIU5HEoB/DUfn77CO59qkEyC9ImIFm9wLZ+ZibY9t9i9o
p4opwLoq+Icc8/tA6zPCJ+DdCrh8e8k+cP6VbWsW+aMNN/GcUrwNBXrmUsUoLxavt67Gk6Yac1Fg
QWzIscOmWbjn7Zc55UZY2MOm/xHcq7NJDeOGhYWAMDSoSU8rUndPZ+FLLxP9BBABdmVg8a6gbNfZ
m7jVxmHPh7YZlidl4KLJVRdAq/mOyuIoGnA4U2sqrwmsd/YMVsR5vkWDmQkWucc2fxlo0HVKf+f4
wOelsjZdf5JBE+AKFzYN1VoL4tfgNpkmr/0Tm63nzNn1NCRxRUGWR9rflqVpEvyM4gs7DZpEd3gi
U0Deob14MC6HNdnd8w/6smopQYWVzmywOhLVUZXM8guqYvAmiSodyogtE4502dPRT9hcsqgQXYta
MQe07UCQ3T2WRWlciSu5cf5lV0IRvWegP1uWDq9AwMWTYzHNj/g43AVjhi2It6rnpDR+deUmKQ+J
lhWowda9v/vdmo/zJnGBEVlijrbZAIJ0RdwFNCDClKBBDw+EkphY0vSEDF7ex+huF6wtuSH5xiHZ
fdtC1CLTBVzHqb9ZkQLPCU7HqGG1CuIPj/hVxsAjHVM+fAQRmlb1PiIiFlfhIfaey3fy7GGM8tYe
PmHsvWvwukbIKjjqujFTs2C21AIBa7Va7biRPMy5iwG1YRSbyFvd0RKgOSZ47GWJ6KUT0slkbc97
WHFIB9GuPbAlzPj94pLZAq8Ro8kn4VonbGddO5GwGrKitAYbZWkkv1Mt1lmoFKcmtGhwj72rIT15
O/Fc9shBb2QMqTTBrMQHNle3pqy9Lb7ZfBhahDaHh09ZU3aa8RmB6cf007zzCT95+AewdAIre78J
KskcpqUHwf9FS2ClEyfso5dYkUuwu1+39eEoFpIQDuBmGmErSYKpaa7e9XtEHm3Vy8HvcZ79LxA0
DR58eegy33WQ1OBTyipshn88xH6U5GbO5/ZvbD8nDnjM7tplZIR2M/xdhrielCpuRlzyUYWEktZ1
dt4lnHiLZwaYs+363i+NNndS86SjfsPYE+jRG0tH5mhBQHtLSMQqtkXl/iZgdcJprbPNpfXNuvqq
E3/6VlOxBx8dhaB2AwGi9rnAFkphcJmbRKBZ4yDzXekf0ovmTOV1IQU+EUf7JDkxxqrPIHq3rB2I
E1Qek+FjivJoNdO9zD84k5KXDjuaq9be/Xhxau8pTzMmDKlE8nLPo8Q4L6hxHfXFUm9iHgy82UWc
5HVGtJizRKqE5qjo2KsL4dGyOq0UlHromxAIdtE3GQzyQ2aAQqdO4skrC/h+oUvH3274W7taJNIx
A5+NPc1CY1zUjL5HyQG/CDYjaGOf6Lon+BdvtVVqR5a2DQuOn14o5vqpvPkknh16eWOHegsxxaPB
V6mG8J84q3DCpO0//nZ9IaG1xMAfQZrhzjRIGLu4XVoh0xqmsqhUGlNO6zNX65FDNHQiJ0TIn/fk
/+J4Rz3hpKrC09yKPKlDbI+i3NJZr+vn75HyTkBOJG1a1rz6aP+y2nuoKo+NOKqjnvBjdiYOtEyj
xuIb/FA4PilKBG++dil3Os/HHGPiWHdg7HECg5kp1Wos7aqt/ca0arA0Wf/CBfnSnE2m3q2Nm8HS
Q4ZU135/K9SmgxDtyqEZcqPyvE8OxOYAZKJX5HFQfB9C5SyT9NvS9/RzWF7rIGQDYHgQW8/L7zN8
fG49i/wvAWDbcI/Vbt9O3Vu9GBc5KjeT9C3cDnzjtoGyH3NqZOyAEVLP2qfsmx+UD58RlQVvnfcq
n8+SfD0RkO0Mr6J2itbJqpX3ivX8BwCvhqpOHntQh7nPQzd8K5tZrUv77SH3LY9IF3iYJt0UkVOb
7X7pCJjYLEvJIEapH2/BTNf02n9lGSa6EVd6lst/Uo3Uvf59OSAG+UeizzqE5XT1IdCc8jMvW/M7
IBGC2ybGFeIpYKEYZppkYDt/B+iL+o5zBOp2tBQBu/B2LZpkOw8lZ8HnoK6YGKRqLBppZG888AL2
FnmQ63CFEPHkvD6fLcGB8IMmzzPC3C5xGwk3wRdle2jK1PLUUV9dtdXIXh0RAK6vgjCftw1qkIuH
Df5pJk3YPwo/zQPuYfauDIFzdPtdbElFKsbxR+NGf2RgNlsQqDOgyzT/6X8s3o/XptqIZ4BSvoKk
rujOIvLHXUq+bnMUNGy32ertmu+T66seHRf5K456HJq+zlXr/HrnK4vTsvVBdEb5op2nsvpuVuRQ
Gb+xSL7EHtXbmzQf0uqkykpob3tOe3vkkbI7wnZVFGjKlioip+/idJQsNIVtmg/yN1HV3tSapzqh
5sjryv5Bh/lBa5bmspC/VjAwut6URm4NvqG8pRWEQ7YmO67oRzUQQaQW3oCIE4HOXJUNEUuIWOI5
466zY+1n8Yj9wKWsY7AglCeh11DU6dUe2mPxlFHpCiknUdwvCceyLN07eQ3f389uHzXqQEB76Oxy
tNNJ/OUTTOVCWqrT1jZZfk6pRfYd22Zp0vAjbuBk0G0tzm14olYfA7bEqH2zdlD6vZ/6MEXSJRw9
GVd/oJdMmDXD3PYANvb+CaRdc7syaB8cztciokNW3Jg3SGOEfH0DiIGTGMjDC/AhK6iPv1jmRRIk
bl1hM8D/jHwpn0oFSbmT8guIKO31ZKUNovMF7oZHuozxzYL6ygedN7pRAOUxrTSrVXh37wDGLf/P
5qgZMvJkiMzpTSDfti49l5p7cXuRua+8OSxZgwROVW5wL8gozTOh+4Bhip0601znst2QZ+rkVUkY
JcuUr84lw2kZVNzv43z/ckhloxIBj8fE6ZIp0VgAcqJ5Bb6SXb28usoSShv/QGrAXpDCYED1yzxD
7kiXGSj4Q6El95DmwMyCso4KA21l9xzD+w3POmJynpaSo8ISNzyW+eNZZPQEG1Fi+FlECHjiLp/i
3/8r/QGDiJUAHOv9+UFm9CzovtHrCP9sAl42vwxhz7BYh6rwcKOeeEbGiJmRHyT0f9RI7ARD2Xk4
D+qW8lu/tzO/IjEDDYQN4rN2yWuYuBNCUwW3I8Uc+jTFOaUwt4h31eJybevVuU7jYpi+VdQWaCyf
lqwhUsjiDoIUCceBXhg4Q6RNSHsvODhmTgrhvezyia/E4goG2bRk8OToJ1qqR58gz/Zb7kRR2wH5
0/MzOFNGe5R1SN/7ZMMQUgMDaRC0/qB2xj7kQKD88nGgddrS6XvW5S68Y5QHpzw9tx9DB8g9XJXy
kVHHgrYEPg4THHSaOmBJqHfOIJOjq2ZGbXAKWBusevL97Itn1yA7XvkWC7r9IS4pKiFKlqAGKSFP
bTLq+ntsguQUWEOKpWK7Ql2IdQqhTB73i272kAea6UzEpQ33NQaiAqnLnQQn/RjrRXj2A05iwxv8
MdltoKPOfgBT/sv+iHy1dRJ1VxTHfGFUKmEwMdp/WzyqQ+GJCeiT5D104o0lG+BSa/t1T6oD4Gza
3dRYRnTnZbxsCJOTR22HEW1wZlsYAGL2LVuyrpUCueyZEnwTAAcvlhXUJtNq6bQtDJaR3d67qnGZ
2IMQSKlCuEqdzk4eaIqy6FHD90UYRXNnafy+Tnbl/neOUk3PcqIzv2HuTYRcLjFHCd3EoeIB4gMS
kmB+c9eoSTlQ1RvtjeciKHIbwu4OPrHC1YjA5Q8EvAXdAbshiyEzNk2LNrBgNq0tIeBMBFKJuk9q
WZkqFWwfY907mqbymxhdl46Xxk/gKHzLJiYGpa1/S7z/2c0WXhbN8Bzj1Aox5wpWGaXCyOVWyQ21
MQ46xSJ++s7gXin8b2AeeVlGJgoZifwNE55e4xsvxIEW+JCoM1tASuKLXVhuVw1GjPRBz+UYoQmI
nkEkW1a4zvVdDRB9h3vyQMhv928zWjoRS6wvz0lUX25Hck4FRY/m7dtLmhPF3n99My8ff/klOvUk
7m1qj1XC3dUtRtjGoRcwphHHyXF3KwPaDyNhX6e1Pi6FlEvj7ESOdXfAt2APlht4GMV+0KD9N393
2VSmZ4rdLFKyQ+C5RNSgk7Ps93YLzX9rLXtj0Ry4vD6lIHMB6iUqgoiZWjDrT0l4GbpyrEk/tjb3
wkQDUWThOdgxdzCG7La/cPFWROXMJnlO95yySNpmr6k1kSx3gjYqHo5wtRY4SyaDWgOj7PIraYb7
4utfUX/h/OwBq9gAyy7nqLpc99pgBXTeOiEiEaw45wgksBIH147+UhUGPIx8ECC6Woh5R+12keRG
2fS7wA8f0LontH3cw/3T5/AYVloA6MRG1x9H1CPSdEQruIbN9tjv8mpG1BURsREvVqHmy9BaW2vZ
Kxkz8R74urcJcfied8ttMoePDai3QjwJl6CZ9cJlQubzBnpVXHLBa0X7pnCQNaxdmcMvFX3oduO9
z8B7HdvosqiekwNahPgFla3L3BFBdYoOEUwY+4HKIKa5osqm9QKlgBbTnsVEtWVKwpIN64/gyhsM
vNOy5p3k4tJasPZ2dTMMGVcniSoukoVrJZ22wxTuIVHH51yi9AQGznhtQKGWM5ynsvCUcSCAggEV
YgCvsN22eDxq70tsxjwd2qi/5xbcBzmFREIEUgw5h/CW2IaOqlr0ymZJ5DDwfHg/uFH/koRGgmTs
vt5kd6h8MzHANfwCPEogiaEcssjU+93W6P2cjP2y7o3RGfejPe1s2e2KP90fH/II/WVNEIW5e9BI
PVHCqawH4jot/NOSAxz6D3M2a2auPtEx6RY8Q+Suq3yAvzTbyt/j5QK3PwN7QW3eGG8u5y8fM9nJ
C7FGzhuKLEeSGYZZuAkWmv0JHQdxCQnBBWaHEpfPfYOgOsFYzpWnRx+6ZN8R1Qpt9uwJg/zeOnwn
ODlXtE1tdGTUM9Y3jmaKfbdMJry1OIIyFAF/E1n2ZzRqlYW3KRuMdbL51NU5J9DTU72M06bAyka/
cttYIjw9VwIfgf4Yy/jfgQW4B60cVx68XJBUdqcuvAIYAOFFL4Z/iQoZKcJGge3dGZv4SJeE1WO5
lCQdXKcn7LVGGdi0i5VJR3DN128PDwip+VevztG/GqLnhzYLcoj/SNKTxHs94F0JHqlqoETP2H2p
G5phdpbKS/i5m+54aHv5985L+uRK+0dMnJIJUZCdjIvlO2oumfX/kSd9tOyhq3mVg/5ezr7HdeZY
xGkUvPuL3JrqTabT2WWh2eUEnvOWdpFhc4ajCsitLSb/0u+r50oaqdX9qGzjITQiHcbEJW/dEcHK
TtBZQ/Ine7Fjs+8lm5afKXiUDshi8M1qv3H0ph8iNsN+6tLu4eJr88xvwidCc6otQVxyJZqNNBgj
PVtfXBr0e5PeKFiR09vpVr47XAlIwu15/PzCeB1WOnyqteOgj7pysUvDcque0fDTC7okEsajc3eO
0Q9e56DJ3LVx2qKXR0z2148l6JA7z94q7P5fzPL1er2Rki1DQQNBpuk4RKx+nN6OIg+FNZq6NTlK
HK+1B0P6U0CoD7dlEq33CWyv2eWOBeGTdm4C5sSD+/qLEsZMxiuVu/DbaWscSuvNlncQ2GcLAEuv
w9eq+Z9TjkcA0k9azSoy7ga2LW5EB4rbiC00vk29EUf2AGNWeR6JOS7MFKMJSPgZ4I52FjTSbs6O
qOOanjzxisgUTsQVDH6B8p5SYCaA5xddh15UiMFbUEMZ827y8JgCZyJajEL/MyI4Ac4CI45KjXYW
HiHa5QZm3je0Ksj2rxz56/dIyFUt636seFTDimK2KkKr8MZqjA6iDT05wJEbRrKpLFZxlOvaAhRm
042nVlUCMhxNxqLZ89F0BW48hc54pvmoNi98pBEEAl1UWrF+QZF18vdElxpQCyrt6Hf2aF6MNDYf
IHlSL/fF9P7KfW0TFOFTafugfO3e6qBGpmm+Lov12hQUo0tpS3AgbmjrOlzR5ONdLUigGb6CdNs8
OWFKuxD4Dx0ZWI13KQVUUtHom23afJLshO5CcK82fjTAv07Ahr9S/JvKBhjXDURRCcgzS7s6PeyA
UysSEl7Jej3CqKS1BVdboF5jmJ6TebivNZlcKTFv0HLX2B9aalhPkYoXD7EQZkVUd1//DHZheaLK
1Vqu78yQlKtUM+fgQfbWhMeSX4OpQLmbfRRZ5LK2dtA/QKIt1f0hIveSGmQsKmJQh1JWUB8Epf4y
W0zAT6eC2QfZ8JDAD/Uot1IWq4DdAGsslJYa1pUEfJagKI0AFrh5Kqx7H59onYKEnCV6kbqYtmXV
5iuuK5ww3o4yMdjAZs6B8PesdCT9YFYSFM1o9kL8QIoMZ+Lsny+LECHfZe+vTc7fiHjZv2qv1qQi
rEmhphqY75BqNvuE8ml8biVioNjJ8P0ETW26+2tq780bOIBkyjPGlosioFgQcppEJ4CUrTvLViG3
y75Z+ztV/G3u/hMnoSPNrpYE9hdXS+3l4oiCsX7ucm91NkgEJvDDQhBseYk9VBCgJCRzyzyEE09G
yDoTytHn2Jw1LHrl+NebseQhgAmz+JenJK7BoZKE415PsCVbTWL5wT3C4aTgfM/0Pc1YAHla4mci
zqGgHUvkUfVEwSQC3yvgbC6u3urHZYzYv5b21KCMkkjhYCPYhi+FZyL2fCTLkCvSBDD8HiwuPhZ2
vLH23hntW+Ru3R3XdWg752tcIavYEX2PeQBJA/V6sBGcmER2B5gUHSROWsZkFy19MtKZaUvofKbk
BFj+IIGdpafmCJvuYx3WdDqslJjYPmGIl7xtj9Nn1yKJxrt2SPr3VeIEWdDN32k6BbGBIEG80Sjy
vUfytki6ggSK9IIjdyran7xx28x82h9eTWCeeX/OksEdzyI6zWSbcU+XQrT4qbiiEXGx1vnDPuc8
iTgtHcjZedX1pwXgUwKEwtsEDR24EmZYDQWMPcYoRxYUdKgswKuMtLv5YxDsI+OnCxpNy544mSrx
Nzess3lGdO7+V+5r6WdcCY4AD/3tQjbrOpUP2TW+DBHXm4GxT/Aahsuq84xPLYrmzM9HOEoj5ZH4
EMpT6vBBpbygthejgWL+16QgVjz6/f3M7pKB1KKAiW+EgeKSj/XrmQN/4tW95SF2r9lEN7xec+Kk
36X8HAVgWD0KqiEj0cy7T8CTFljZduevAK0sGH5fmF21DxJffpin8fv9XfVyvQFj6OQw8KDQs/lS
+5i7dIOETrOtE4aahYAh3GhOD+acE4zh4OVqqXbCAK6sc+AwSNgLfOEVUX8niuPlAslk2WrVUvmN
o0aP0/pVMgVndywwjCXyztpSl7LDMQ3akeLT+pHOB5y/X+MkUVMYwFgdOuDMeA7FNfXht3Pw0YYg
9UdBMeBcjWBjPWPAmjhpIZgFtnMvFD68TzfT5r7k3R9RC+E98eNI+UnNb6Ri/hrW34p08oi0h5/w
4sST43NtGNLwfGXx9hhKe6hEvjpOhpDCID3GkuP4sywuz49eq318Ds0/+1UhDGerSnr8C7GTkpn/
Ea4OyPGtxFR5ckASKg56QZzvbFbqdsQkibMZLpzhMTrYHsfkCGjCJrc4QcLJjTlj5xXdmTD78cYt
vj/Mn/7JSe3lyj92aAXzOxH+KInuWS+EQWxdUitXKppN4VCnqeZAkJyEkivOK6uallriQBPJ5XCE
P5Wyd33F84D9LmoNJIHAEoo7ja+rwTihutytPd0BmYowNi1dsr9vUm1n6qRMqLw1WNRHgaXkX7Wk
RP1dluarjdJfbXvTQ48osCPblPviNY7uRONntvnKLIbli+B3gT9M8u2TXOGu9tf/42Un/u46mxeL
/JYnPF7WJ8O7kMv5mTlcBP3uf9UrWybQna2VhfKOD7sJinHaLT9gnBD0BD8C2h7MKIkTU59kI3xL
lPGlPDcgz2bNMDN2PRf+vA2sbdjlMYWKLnYkLjuvpq+wdtjnPugv6yh8M/R56ryvzIKlFMWfhAq1
n41weNpfDvEhu5/uiQZxrrMeKxxlum883kSWSsHme5iyIMnmmzscLIJePCOaTS5FtVFG/waT6hvJ
Ws03kNQ7uk8OZlMevoASps5d9XJYPzlU7M9tgMyRNeqSzGx5V86ZSL9ys8MSLvGzQ1SD87ou9T7O
x5fg5ETAKfw4xu30EXxDwl2c0KxnPGCeusNB7eel2WOBdYrOW9eaLiEG+muzfL5ZdJkzueoiLYEA
OXE1wwuKNcpQfdJjSghu5GBfKcirIBuI34Fn58yDFNil7NYT9yw/FJs0OrWnY/NZqPrYaKY5M/1d
w0Lma3/M+I6/5eKOH8f7bMS81O/ve9pV43bF2eaGt3cJmNqxS4kJwXhPeV8Q02626lMJabjCLwN0
xvrvkX0+SlqWOBdsnKfTxKmuAhvJ8aGlKYGNJIsXEWdBFFa4PpxGHPxx+nIG5olIE91CLyEt0ly8
mdSiVc6O9l5XjuL+Z6ZN59KHS78FoJFE9Tt3d9UklZACb8rxTngCxB2dE6tN/TgZWF3sCu8WffuR
yc6Wo+VUdKpHYpU4sdWnBNPxxv0hkxZrn4wSld/W98aReUdYFONwRjcgSZaQ/pPFyBoLtRTa1o+4
eeN5auGlpcEwARMzAo97NCICbsVtrMGT4SkfzPvi3ulWvFe+yoKXyldzzenNf6oTYmMduol3lbNd
KHjqOSd2+2NFQnqi2oTVesmj2uRf5ikz+91Q3qnrPFbSIkybtLBHqYd0C5GPq32+n/Dyn1GnYuih
n/U0/WIbOGbIpnbSjvPOFX6A02vtX+flISCUfHvtfJDYFPTXCR+qsV+98F9l8DZ/8AGSuiMQL4i9
yXyrVuLJaP7YDOXQC9MYKvBMFr81S2ErcOd3/gnp8Ns1BUo3lE7Q60e8/pM29Pjfz/crA4QKcn82
E5NBZsPWiRco2JrHfADbajfg65kTFGVCbzZk1BjKeq5vB2irXfC1llc58vcltuFo+eLsQSgBvgIF
x1GTvJKzEe6Aj+RksAXVqSeb25uGYdb/eouqC8VfzfuR12rsXy0ct4Vz0F55QsghmMD1/cVDD9bU
p6uAz0lvoGsWf+y7itQeL27fqYjIlIJRlMFRs1enfONDELvIJil/Q4D/OCgLElcJ649PurjMRrEZ
gXvju3kq7wfMUMUqQZV5dr5IFaGytVA/b+EbmDkxJe6oNL5Ni0hmCugaXfcaSSbiSEAIchWu1RwW
P/PcN8PD2naTkllBRsmmLQAuoiM3UG+G1CaNf14lfr/MlCcKpMWKEQk8FAkPzs+Z6OG+F0DwWNOU
OJI7OydNl6gcYub+bzXzLwySO2502F+L2GmSYr33onBrtlJETbtPwWybmWn617YS4XmJWo5EVfmv
wBIdT6wixwRVNjv7WUJKd8a8cdHRToAX+cTNVgcKLr/Nz4YgmGoa3HBNR8IoDRHhLEaSPpsF664a
G4rn15Qwbdnsy/MW6q1z1QsWhyRvZYz1tmwnVpDX/IJyRDJToZF2nCwGEUS0fRvvtsybUL/tpZfL
+ejcl6iIZs+xPj8C2iUx3cIulCz3vAjDRm2adibTry46HXk4L5Oc/OqMZipTgBkVzEIPBw9qwxs9
myaNowZu1FrTJo18mnQ2o6fbAfm038TuwSiwwrtOSZ2Cx7IFkKrzUn87NnIbiXTFBqYehRbiJWcX
aspYxH1hLXf7TZoa/O5kR9qVn86AC6HINQDxlCrqH6Tk+JXStPcWnCXxuV7mIqu4n7hNI8oy4iW1
jOYjqC5ok8Pxe6Ui9tX2O+XAXJDI5/gCwZwP6qu4LPKg7AM/SKLG25yzMtGMFhaRpnCeC7gLxYs9
PtiFX+tSMjSVSO1r0bcv/IgVby162bh256We9dUs1KZMIqbndjJbUcNdiAYCb/3bu9Seq7P1CE3J
2XokpADkHg54XXVD9wWi268neBfpYPl4rQBTRG7QJeqIdKjm0AL4AI0moT3YRBb/pUbKLn/e92DY
GVtIKBqLy2/SwtcsPlOV4k19Dd6YCbx/tQy06sVBimqV+vA8sJpJPUn0g4dHXJVDSPB0dDDW9Xsr
DKJgiV/bJoBgnqzYvLle2TCnKPabAz8wopSk2rodYZb4c7t/2EZFCmVycaTIPAlpO5GSslqqvNz9
ZLauoAjSiybPAGVjU2EwaiU0SCoV6v2XOn2YD2P5qcgWwm0+9yfN57+A4na/TmBY+p9qX43+F7yy
KyY86mYduS1sti2RkG76vV9a9Yf3WbqG5QkAYLErGgX5C9Al7xcftZzvxlJElcxKBsKB2wgc9aB6
Dau4+iMwy6REuXer6GGC226bs0cto6iRgg6iGMO3ME5eTwozEfiGBRNYhPwLWu+yHfP9sOm7+kGJ
5TXhSbaWgo28Dkc16J8pLJ7cMQVtPYEwh8anmhyO/E+sLaVNeFwytq0WJjnVdL1XwYSMXgz5Y8f9
zBjTtKTor7+xXUKlnF/g1lXFWLkMNsl1TSJ/wXzdWNgbJY0PQc/1HqcZQDNzZn8/6yoHdV3tp+1O
JDN5GF63JsL4Mok+bWJeY3DcLHZKPLJg8bvMYjkiKltAZM5tc1ofWdSlFEGVux4somevVuarjZ2C
GzLH56Wi84xCoTbBaGWME61fXQDHGvKZAG8SOFH8cCcHUMG156AQbl9lAOKXq0wxlUQkpOHrc08L
zfFI1DU0/VJ9UJa3x7aeArkGX+vj6k/qDDz/7UOE+GpVuFkn5pcmWjguQWbW7k0ZfF2seMGTJyyW
ril6s3Gy+qVcR60ZhD1uTGMBxB/nLxdFUDtGOZz3HDlWp6cACIGT8hQqr8CC6LtT7YZ37WyqLjM4
ATygs4sdaR08S1A8cXUwKkGt26CxKTVoPacVRN9vWH0BM6yOb5UOURI+YNlXwiGveCMPM8HcSZ0m
9AxEWwNxZH+zbYGBdQ72Vpcp2Iyw/1iz502XFvXEdEJX59zJwn+6YCJ0Vp8c52O/siIAK7PNFRUi
nzC2wDjqYopiTMShd/HkT8XFd1tspbkvHu1D7zW9tAvAknx7gMtzoCDG/a1g9r50Ux6r4HN4LXZd
LB1BkrAetmn6DFU2SX/jSdOsrw1NE9S7laZWJc5Xhh0kupMuF0FO3ZmFCeMyno3Cx6UkJqunBi1z
cc8kK4n0DR1vsLbh2rvjC/jIlPQLdkxEGXUHOflursDlXSegU+labBs+gH9hJD3miqWWruoFi/qi
8E268Lp9oL/QNDmyExHw2n97Fh6g+tQoKlw+W9mOTQ8dXge0hEjtmOozCVR3K4GXU21uHK+H1Vd/
kciedHIBWBx7VfWq9NbXhrF6S+feBAkY47QJkwdtmeg7t414I1sWi9eoHx+j5FaxYxMC5vBzf1TD
U7qEBN1rDj0znrL6yIrQadEFYgG7Dp5bZbB3tiQNCMf+yWbx6c7JGJbdlHMoQnUqr7j3S5X8fPLS
xlupzDjzileJOQJKWodsB7XeAjRxRUwj+wl6/1xNoQ4stIBWsFOhlHAbesqIQrLCJKW38QxEUDGS
gO5Bp5GaR6c7WPaOedIUjF4yOrFM79gOdz84JLfO3TL0BGlHtfxBSkE1mc1xwqCD0KJaEI7YYmKq
3yq0A14+Zc5A/ny0cV69fnlybXESq/99yNvv8LbzgSXi3e3QgDQfHmF20RRgEGdHCkoGHhovx4UP
fOPCaSrVjx41qyId8YlA9Owl9uHwv8RbKf+BSNN9Nfm4y3v29qt3xASAbJjnAwqH1qfE0JqSxmSe
L6gIZKjmid77prV3s0bmGoeeaVJzCtVEh1EHKnygmUyAOKuo5VS0GkevBgW01Aegw1C5DyVBxE8l
HObK5WOlCXb4BymLgffTDTO7gM74/p7uNpjALhzo8DbYRWDgygGvor6gUv9sJNhhqmvNJZGNYdjL
x4mDJ58wQEo+OSvT+LpMoMdnwAbvrf8F4wNiSHdzAttXhDpLSqEQfLlpvGLpqtSjAO4lUmM4po93
iP9/R+DtBmbyPTZxcnsYsxZtTc/AYVy7eBfeiYxdmRvxU9Rrhh5MzUW+5eBRFUjNm0bgjAQ130FV
Q7W3l7HXCDLblgBrgVmbcv4j0hdAz1q3laEOI5za9UmdY6NqmdskWOrtljG2tmN5hSo+f9GFyWZ5
KE9Xv+PxxLWaOcq0K1MMtlNAEig97g6S1d3scW++7IodZzQ94tnSyHl5MismmbqtNSf9LUHKnAfO
+VgOf2YrXWOHLwDZ6UJ7fjZ/O30rSWYefeVEIjajfKX+2a00bbThAPYsp9pqiaIN4U8uRd2UB1jV
KyBVDHqbbIhGtIk6BSgz5JZbKa9NRBuvAqxyv+gGKvrhYOnGlQlyq1KAhrIJXECtDy1PyNoTcZyA
+/omH+h7LBcmRpLImTGJWNHi/72szLHtGvI3HzGeCYCHR7p/Y58fXO+0MlIdZLkG55YwHEeN8QUp
k2NO5Xntj7AGmbN8tOFci/ZH0p5OyGMQo9g50WHNSDidl2TrYJMMxcKcpigbFao263d5Nx0N06gm
evtuxVsbbXEwhNUarIm/FvSdOUNuudLi9kK3POIKceDcDlXkHKXsUqog0IOB0X0QdIe27KfNahPF
b8Yxl+U2BiZKTQmWwwRUNAeaFKfPBhd8sVOwuYFqWoDCpg1DCqYaadh9VnGuXZ/vq0Wn8cVOGg3k
4UEnX/t3FacXYl2sSsgIBcrJhU5ofjeaWtqGVkUEpgmc9h97kn+nY2trNGjP+nc5P8rdCJxlikRe
e9Fjl1C1KiBMVLLvABrjHyKjGiK6qf6TE1kJzQUCJdCgZ1rEe6Vob8Cd1g6lrLNUHk/aFfwYEjOc
2CcejFBGVqMj6raf+xzoBdIxP1QoWikgwjcgsEdgWfIDlCRG4lDkgACKCQ6x9JrDn/HXlLh8chUg
CEUHIFjSXddg6hZqp9z08rnj1/EACJDJzI+pu8WMd7Lzum1Yed875xCVgvN04XSGgsnIrrEBFME+
t96NiTHiodiN8Dhn+hNz4wPr/fq/BpbPrcEgvqzfz87QD/gviO5NMDGZ3Tp/FU8aQ8YEl4lieGrs
CpKTNOg1mP/paHHlg9u5Pg2f8om9VP378203mQWpZ1Y6gFKIwECrhHCDhnVKKX+T/pHzCC7FWqBA
tkTwaR9BNIafwqbnoc9rXwWiFuc0lZDaknX5zUUVhooOqpbPBJmWJW1yWl68uxLUNj3LSDemSDnN
lA5xsKh0f0DaNCVLN8AmzoaRJ44fRUAOlC1OmiPlqo35c2zyiv2lh6lRhZCd/l1g5RIma6Hb4hsS
+YRjATiA66BBO5sD7NwGFrJw5TQVWevg2KUwFsuFHCPaHenpnUyO9hvMlofPdkScBbGXi6/LxNW1
KZ/+jQdEzfdZZiwgcmarlNasMf9oKOPwOnfiuA7MqAphr+wKzCw/pKpnwGxuy6KNe66XKmAl0CbB
jA+seU/xh8KNhnCBOG2S5nJa8/8IOu6EtnqHHN98t0eWPkJaaOZ0aHuVnRLWPFDaJQwZZa6SXcuA
LiqV0mxyMnuJizw6Psu53mBEmfmcr7EP5JGI9Fh7e15jTOvhNPwkBuE/p1AR3d5TdUciYdqkiC64
ZPE3Lv9DpYkJHjwhv14rUnMIgzyhTsC/Tth8N6zq7aJtmj26IhF4zIvlOO4WjDNmM9XKXaAHLOZx
/qWY9+CqPfDSSDQJaHCMsuiQyX4NlwmqVBrf8g39TJf2eFtQuFrZREkVwCsnPmk2TRMYIFgBY0d9
480+DRQRdJe7Qx0st6VhwjTJ+aaTuP9jo5IAnaBsRPEkJhrn7LAON0Zl0l8tF2q/u6zplbF8SbAS
my1LBusX8WFWE11L1Bygau83YB86TdZ+2a6LiIDjKqvmccBpRY/6nZVQcdgXNDhxS8JIxllJJ5Vk
8ub5BG7aBIyzQMB/0kMcGkIhnCMQLbkaDCkpQlaRc3n17f5lydv919US5N/yZwxWGNRPbYbK/4gj
F/JqRXnkyDDIMhum2QKAhXdpatxcD5fF+6ZG0ay5m+TgxPZ6AZi2JqgEYOXAgi/ZV2ka0qZC4LTU
xbrZuXIB0OkqdL2Jb/guzKVKAUtspQ5lb0kcGR8DhtPz+xgwjUQJoV2JePHdvGKYobx9JNHLRK1h
aiszTh2F3KODjGiSxlkZfXVG11UChHMSOCK9CYilT/eBEj2bWR1SvsQErX96UwSp/SH+J64WncUU
n9ukhh9y2aRs0qM0dIBmsQbx/1RuykJ/B+cyw2WVyxKDc14EygHMPo8qLILEoXk9rpBA94cKVBlz
sle2e7TFOfY1pYl2tsXiRxYNfVK3tkdDchjqrClFLqb7SLXPPv9x7wQyeP3CenO4LSkgE7NDVQHp
cOWhQV80N3W9TakJq7ia64bQkT8t3jURZkc5FedAtQ1fSnhTXQIwTKtD1xA37A765veAHyU1OVUY
n6FH0+OwZal9Wio3OmEn0hB0anlSl8iQ17WNN6x1pbQO+Iuy9JQYasha5pMq8Mg82h+YgOrFL+hF
Fwp0VAV5KugCtlmfVv8X2sYG/SUMv/9JojhvwGoF1gyqSJHyc8jAZwu/obogfXlUpnpTuy6V75FJ
7e7yW5L+ydu5fzrO9zYm8mBOB0UM9XNuvwwTgJAAL+AwYgP0DTdogj5D6kMptzf3KEsBXvR9+G96
Gphc+dwHNsqPlac1eJ0lV56/5CDbPL2pIiS92una4RDd9q/weTniQXi5vKaodZ+wxIHFtPh7gE3e
uYKT9qiDFooGjRwdGf3SWMnk+6wZDji1hC9j+wl94VN3zJrIH5dbHPL9lZN8kIA1PzdTvEzxFAnt
R9FtvPmUv28mSpNp0TeBnffgPd0ztmIiEZS7AyqoyEnSuLe7sMFkWWNTagDM2PmWrXvXIMMli8bL
MllVj9cBxy/zzodDPrT9/AbFUvw0SH3TDBW5zKablFbkuLi/LDfknEZwkdt7riz+qyFIqc+FSl7N
Z/8g2qeZ3goD+iYLqkr8sfxFqvupj6V+Cg2AuALLJDaiKB0mTttjhdkQgkYYyyMkhdD8W4jxDlmY
9YGXtA6DIkfI1Uf69PibqyrfXK5zKo4QDbG8i9n9PM7/eBLhk1RPpdnpEP4RqSw3kDmJFLRR3dl8
KUhu1ojFdmDH0QtXzXztBxh+dMI9pjz/PMMRkmWvvZwQruXKGtHcqBk8OV1LGxWw7dJDqMwCUleM
8WOxQYuc3qL6mx8F6l3mAFY5YTw36Osqp9jQeY+4KEzv2FyJmnBxyooZ4feZSnISYTJplbs6DmgS
WWm9hIgMVJlIYhGAp7yGA4GeD7R3i0X7ze8aCucXBj9AJLiQpCf5oNs1FjAZxNhiXjAUBY6wOq2x
fdax05smI6btSTi4/jvQG5ii7W/jfd83Vi3dLyXMgzU4kzBosQ8hpuXppuFoJoX1qlb+F7Z2niK1
DXtA9Aa1cbL0ejZgTJll4CqfWPPtjjE1Pctt3GKR4jt/S0NXdDwvCECjXgnX5oKMXBzBcV2MebnJ
aoXbH5TjrK9jqS3mQVEkCWULAkV/lBLdvjGGY6odU94vaJpeDT75RtfI5eMCpYSmds1vw5LmgVA9
+18ndF7nOcrWQlQctBBou+kAsqC3P3xBkBDCVTRjepLznNE7ZAYmMyDXgv4sFCeEReJM/gCrpAr1
lLaHx9lm9u1wuIk5fhiR/wkY6Ja2ZB7hMPb+rRWSmRy9gPFOVfzIsq0N/cYefOiA7u7iiKgGVcXc
Gts6PJcSv7kIwKdu1S9PLxGYLgC0iOrplBcc1g/AR4fMo6rBAu90ldrGIyfmhQUoqkxX3VDR3R0O
UZrV1NJbBBRMXARKkFGGmzRC/OajCS5PgnMPNgMzUZ362iVmo2G4oAhV+nhJxSy4QiqVz9cT2+H3
4gllf1Yot85UzyoLJsTtQFpc+JlWGi5VBH919eRRiphBvmkXM16K9m3sGZieUuvTvOG5RxOY0UZ0
Y1mRc9akWp5rTPDx6xWDyJq0pMeBVP998NiGnimVFg0VvDOoueKJpaELzJWoMyf5y7pgNL3fhmKi
ffGM677WiVpAuE2OHBhwmkYc7JCmRNJxIh0/hPacvlsd6ETos0pyaYkpzKUxME9lU8EDnUiR3JKJ
D1lo8peZGfegC9y5o3MR1ZPZ62AmxcdiqMEBOzivmgCPoLzPEqAB5h73+6qQWIJ2YWrt2x1tsk2o
G381LKB4ciZf5jkCvGLyx7Xv3S57+UxKxx1tsCxOAb8eZUQQs4PtUlqqM0mWMTL8N2WzKQ5m0RnN
4LYMWX++3eAt2Ey4SKs95RKIau0XTBmejGfnp2Ky79XTicjOVYHHMXdDySTXW8WmJ2IWvEBA07yQ
Myhgd1eSAkRRGEIWAev/3JY96XeT/RkPpXtHUX/OdvVXVuamTSUS5YreoEIz53qlbHxztO0EVDtm
1GXajVGoUHVAf93txtCrsYJ9jCGt19KYxuAGWykMUmMuZA7ZvZ89r1fe1jEzaGVIiB0P/9wTdlY2
e3rc4lAZaT0JVePHNCv1xErs2O1DzqK1NZMxgv6i2FzzTuE2PTCgxX9BduvEaDaXX7uVq6M4QXza
+FAK/Hb06y/3TQK3NO2iAUL+Onvi68hXdv91FbBriyPu+wfwWxoZrv5NOGcQZy81py4G7BdK0hFD
9BxRyFCv83O8JkpnRwwdGxao4RPrm1CGEaKVmBPlVJHdJOhEkLp/z/VdshtEiRZZHQZ5tO+m9RTr
nVDcNTRooySCB5Rka2FPl6+Kbq6ahAJU28GIofILHtYuDz5SfUREGmlGDTN+1gh0gw8li/YedmVD
leUdqL6DpEuUIaFEJAsOz8CdiXtR4rdYtgzm3zoAodjwWGbaifJNkdL1AjrSv8VYId+NEqDOVr7C
4vrdatkyv7grygEEdV4DH1XTq4uufg6Wy0asNRTNNWGm91icDMpO9DRVcrh/+3oNNpymFwjokqa8
idIyVmBHqjXiGPEXsQTvShHVxyqOn1pCLdi0umRsBFzxL9jGQb1njnR8TcfVNcMbZKFQUyldqtFG
ueY+zishduUdb2MBteyy8VgbYJLfcIi4hnsqGHeiJ+boOB8bqkLdtWi4ts6qmai9NAUURjkrYEAR
c8XoqmYWvgavwWgHXWb6D4rcqJ5WA4UdDpQQDTLbMshXsazK23f1cL548b9WdFRXylgFhFR+0e6t
RaudTjRbAfBe15spJKPT0tmcHkOH5tDXJ6NS46M8FptBMRa50IJCZEjoJgMOhpzo+zFdH2x95bnb
M/NZj/04Htyh1xYc9RudV7wQUhLBB8w5ZPNSqDAvY2zyjkSaH8D39g8xuxzRXBlnPTh6+Ch8ztBZ
vO+5BU/X5ex0roXnpxWL4KLW+kXawb2ZGO1wX2dSdWJXYIbfU4OeEH2GrCO9FAcoS+kzc3+cOxfu
Sa8Mqk4EoFQGM0h6Nr/p/37y9zpuOisuZ1njeR5mhQaKDE12Iws5kZ+mGksUczpDK41T8EW10zz+
Nn5vHAt2XLPfY5vM1m1+XLeei2mKCD+FLiFOD3dvaqkKDydPzcBMG1n7t8ALWIzQBjKN+OQlrCtA
5+Y2Iaofk6UHYrzRvu76jAkYOyJfG38mVl2j5AVU8OB5sfIX3m0fh8xrtRJ2OtDAWBGt7+fUzZaC
shlmKSAcyZMBUBoqY0s78Qm6N8A3m/XBqRlmF5vPCHYyl1ec6IlLu3w+QWZ8Rrz9cY+Gp+Yytteu
N+1nsGBp7Jg0+bZWYIQrNfSXp32VI4ZEZthMWV4/aWNSTnU8oSrLKIggzcRFa+7fUpU2/0qDVgjA
vYImK/m2lgA++kn0n9Qso+DQMnSrvYlX7TpHqgigyd+9yF5zLeJYuSyZ9AJpQWl/vqP4RSFHUxxR
9gBtG6dgH06crl3z9EnRiyl3ZvIdH41fccvcnhdYe7UPR7GB+4aTOa6v0fNkJ2U6cPK8RQssXy5i
l/XwSIT/IuHT/OvZvPQWuZMwIBSkjnDn5QLpiZoGVRExfukkMi2fn8hrQssptJgAUOd2PmRj+lA1
j9EZRVppcocZWECT+mZq0xlWkqJWPMyWsb3XWl8fJ6QFYwFU9ypRJaVQA9rmzQXmMo4929MOxv7L
IWkMeU+UOdno/pQ4MnEEtXH92jalk+nN02sfS5DJJlIAuBx0XBBx/tQmA8kExxCVT8htsnuDi3zN
e89zXy+dwrFNJLSURgb+fxT9bPKlJH+5KGzEYdmjuD6RB/xl8hOh2WYMrRpQh0+kQ33C/zFVs4mM
CjDeJrhIHc6pREv0kKgm5x95aynhxFpRE+j3kxsHbcc91q3QI+dR+xuXT884LPMtD1d2khaShgtF
XDmXrDE/5TTg3J4ZHCzvb37kW3LFC1R9+k06GD4jDkBtptcRKshxg2+d5R+aF2lRG0//FHg7KPUE
cH/TzwG9fAf9C2YR4rR0OjrfS/2H61Ykt0XFzqFW1qm3AFsPz6DOcKUCxyxPFcWiZkmdDwuQdKfs
qjPkx6yJcFGjxXLnMeMjOsh8cGUZWQwagPezEG/QHr6ipOEdaiOZPQA/Vt1XfwIZGI3kG6313A8z
C0YLTHHdL+rnFZh03POdcnXjfPbpikEtUSCmAR4UtdKuiVn2jFIQhYkC3JLRMkqZ0qZRiEP48Se+
kL8nWDWvrZAc4+BG4VT5FwW8GgdGjRsX9epqb4KbRwPZ9erilwSl9si5mtR7F4NMwfnwEtQGETWw
T6hgnOlnspIfJXtaY04HkD0mQvWtC3vVmS0AmZEkxLq1yO1r3TZDbCztuUjKYaG2HS/Uoa2yWRiJ
LCUQDcNoGGgAEe2RMoBM4iadYI34dx3zZ3AaaNMxSyzIekg/H9/zthXyMI69++fJ8G8L6+7hQrFA
pcBQmhrjoTmYEo8Z8vPYYPCpsZ+X4ffiBcIRVr6F6ctsiu2LTWsPt6/WkQ8kj5D5hARpRM8qeatz
oUz/nrt8NAm/Poq7xG1HapdFs5JBDcT8BOneazYzQlNlPDvfjYkGJVi7KVTEiqZMpxI0ND2luwFZ
jRP7d+MEMCbtRdGuk5ghxrQOp9P7EFXL4mRa45jjAp2m0yeynQrGuPP2R4K6/oTeD1FlPtd9TnRk
zBc9SDizjQ0JbrixkUFSIkoZlVSkC5tNbPiz2u88bFc2Z8r/BIMQ6pFl/r8WzFCvDwjrIPe0Cevf
YiW1vNHPdecwKxkSeZo3aB1U9KJcIglfx21xuoTi+jaqq8a1N539iHsmL+EgPMfaw85hWbGohtvv
juoD7bqOUb3ezm/VeSy+c+FkuIOvh9Z1sjvK66aBVeybCsgnoISyNf0cX1j++TSP8zU6M2xxZZpm
17BPoXBdQ38yahhd+L2dOH4P3amWGte2HE/wFF/nc0cTZeA018ey0YPLECVm2iKDLC1slY3K71kN
NZD3QWXmjkUnjlZAm5eB2mIhgtYt0nVdxCI9CCnwUTPPFMGOeaDbGoBPvWEX5hq3FTWUc5PDXbD5
Ittamcg+wHEwt1pSMX8wm9LU6mI/tEt9otShRq5kPbYUnklF5ehlfMEvmeVXXlFBB4rsZpBAcxjd
f3bNbItX3oZGFgUACZoT2ELqcLbCEMwq1si/aGj06sC+WITzR35cN0PywrEV/33f2Z5ntC6MN2g+
8NNwp+n+t6Px+NIk3VvGufvDKRAlCP0IjUK2js3MGdUqIrC9UupqCavKPdmNxwKdvCgNvehQmnmB
DKQUFbXVhhBJEyeWBfRdACrpUxRjizeaKQmY+G6JJS+zX5Cy9UlX0dVl8yJzGPlSqOAb76ifaCtF
VzNIRJ3vy5kzm8FqCEM8/3gyCTXJeL9Qz+p5/mmLCIgv2tqRvAvPjocTiBXqlduJcxzBc/MmY0t+
zCpp8OKWKLonSBOTbLbKTrD5jM/yiRzgEPLX9L9wn5UZdaYIpPMMjZEYHcAcfLGGjPyYAbIW6kaS
QYnIEWYTIk3+NnM/Y0o7Q6g/TtCco7F3RPbhsWPwK9nj36egYTVJJ1v0ARbDOBlS2Sdz2Oa0RZhW
TFgHbw6Wk8NM2ky90xPVkPxO90EOwmwJd/2fBPd3y6yn7lVlvu8GCwjumsb0jfzPuaoLJssFxsDZ
gXQuX3wNgYIr+wXXi5Laeol3ZfeyN113x029eCygnH68DX1+6vbYn0MZ4H7HnGrSe9f1wWACK/99
gG/q8FaIjxGF7ipBE4Rh+OVLp2rerAT4Z2p2ub492PtmLCDETqkf7fTOpt9LvUDi7lAWkILYRrIC
zi16T1/5NMgqfsk9idr95Fp9nHdzn8Gs4V74nqKknb7iBi7I2Th6IJ7KO+inJzL+bXsoZIyrHTOQ
9FfZ/SaKnozGtDZiNASDXFdNAtNnx47JqUvj2OMwa5uiGHRgDcGILH7v2Z1liP8cSDCKiErbHwT/
OGmIrD/NdiwJ083oUZEejFc4A/eSIUhDOl66M6VJsTTvWHpQGIUZvP39OTEwts0D0Zys3a6KgIv4
7fGr737NCNxemTiLGBMHc8wdRqnMpGFh2k4vOCz1TiE8SYiTSv6ZBzUPuQEfNhJ3/tgoIO3arrjF
WPlM2knGthvHgIVlcdUZPs/iC/fr1vAAeU8yt06RWRA8UWf6IEiqMDs5dY4gSbD9KYYmdaFih+gk
amZrDPhdGFumCtoWIXAQF6Fa+YuRofr6RIK6SMK9i7wgYBLsXzJaojtULc5t3DaKinDZl/ETym99
4CZDzwKDCsyDpfN23S8sptxDhmG0sEDhf7QMYSdOCA1/aihbXhiqCBcPPuT72nAqwwX8OVTcult7
xXXF4+DEZzN4JHPZetykXk5+UBuRXN5kTYZyVVQmJkuZpHiGTn5JuklAtW2RhEyqDA3ZbD5o4hFD
kF5pR2mPGJTsT8nIvWoKjXIR9VkklkOS1ssL432V0QBptGYRBXEOm5+oiXRvWSEYgS/3x9fyM2ZD
NwHMY28GjureKwZuowZ1ot2wcTB/nA+/vlf6yvxZl7PuCahRYhc5x3nCwUsp3n3OMwhSzuZOd5r5
zasK2vCE9SOL6TKlsmSZ/tNGrt3RHr8jPuLNHJEBKBPDil3j8vOOKgicCtutoisuJqPcAe2A5e0F
kB/cyqckS2g18Q84uDFb/0zeEBfhd2QW6kwsx6/q6CbB7fmywGDofMacEkGOJNk4DZufEgG8scMn
UoI4Cdb9GrmI4hGbD4sE8JSz2QpiwWsOmcJ/VMqGJdv/EEX3mPhcLPSSf9nRjmfxqXngs2iEfXUO
aM+8uF1g83S0oy6LnMm2U2BuXge4XMcdpjKR6qGuuWWUGUAHqHgv+o2ZPjh/NttPlcDK3o2IOqU/
d1+pTXKidXlulI2X8pDXgpCpjI+5N8DGTXDAY52DFAIEWidYYcJ5D1OA3HQmgyldwg8lvbkYVc0l
0W33U74fSch0ObaIVwWr8V+Q4uGYXaj9VBm6Byq+pMsZlLxFp9kmO6W220ATQjgM7cTOMhL9KqK+
M67cBgu9ozwuEtBclY9F2JAaZtlbOPAwTUBEgxUxUy4Y4ejA1V2P+bwc08vcZ02lKADV0J0J6YyS
8ZWQaT+j1R+JUvd8G0VZDaIdUT6jpspG5ya0HkribiyTzSxSMhabVv2lRau4riiqCHeltX/OTT+j
gMbPfGU6EzcDJ9iCV18X8CWTHl4e3aTq/To5tN0s7lECXe4/ze+sJTZBx/o+AEUXYRjcGobKJtfL
JN2/9wtbUsxScSQq5YIHSNoroNYn1J1muCh7Ri9SX6G0m2ZriMZzFSNMuEa6OU+k1FSMl9F/skSM
WGnBcXryIvJt+hYYg2KOtcNhpp339GPoWEjhKHjZRUnqBToBhoDH5XmDEgc0FG3w9I2XVMrcx6YN
VvXH+7rT/Vuhn+BvzPFn3PgjmB/sNra5koJwhRtEiFXTEEs2hvVcWCsYBUX/bW8K7JW9PJVt5W3f
Z6ilAZOygEjnQF2JSVsj28Ubwm8ba4HTwL8HwZKyiOmsQ8/LTwvTn8SqjtDj9nkj5W7EA7bexih2
cBmD6nk5pco8EQFBqpOFhbfHvQCGrbHPIdIJFD1eZHPnwHAcr4zGRa/gwC7JKt3D+OwQrR/ykQRS
EALJQACcfXTV4Hb3jmwXdEd+RyCFskQkVI8MerIz4NRiiBtOfE97R9LJa05YM0e416nRoQIifuNa
FILsBdsdhJzyLfldNkc9WG6KM5I+d0F3geXzJ+HIFQUDEtKfHJQVIQpEzJNNvqYIgcS58sRlhGpJ
b0us1v7xLUkyB9tXtTZ0JzD02mn6oaF1wUId/N3MDHYJwsR+xqVchHHejMnqmmC6ed39fIBELpOj
jK3w8aftpaaLL3fYzll+xZM8G8RjVqOiCraq4NLxbccCjohsenmSkMbvg4bzRT/nZE3sBkfBgOw+
M64F2sRIxpff+sdiiP2hz1EMvixym6EW/LXDTWjbSNndvWpRjoI4436mB3FSMTulyQkcEboRJcqt
r2+7LY3rotAIG3fiRa7SFtlV73xvTU/HU/ryfsY5OG3g+xfxrZtCrXNy5Bwl43nRIGu2aIgT3NUB
El/zYWTqDuex3eEnHNNtbHslYn9CIhEMse4F3TuSonGgKOhJmVhBSWb/lBuYaVqqDsFMWS2qEzUn
fJewUMEbyh3FvXa0gZDKH9RNRU3NERYzjzNoJWB0QbnUGM3DEAvgct4AquxZyie6Ony+iAx/FDew
DKpVxkt5BxP8eHTSvT7dZ475kpoPT+XJ6Kk45a4wsgBY/bzh2j2lq4SZEtIBkCvy4B25lKQR1y14
5LGJuvqTZ7s10O92+alwlz0iUyID2NSTmrIz6XeR8tG2ESV21dMtvmeZIRJx4FCL8Kd6elANF7RQ
OaWVosWJzEfaglYe68Y5t37OCEi5pcPTMjcy+JAVuhaW3P4FCqQpWraGck06RqdLFfZGY3cXUP9m
NU397nN3jMzFxAxulQFGoTwr+or3+3r3EYPNLSlFLJP/XFMhcPFYgzfZJy3V9DQk2ITl72IfcvGB
rQpIk0Sdb908h7zp76w5aLjmTL+KbLyANG4rRKltYEM9NXZR4DLdQez1gTnjvPOWvXODc+eUboci
LULN08N0ZxKfB4apjtLk70Vbt6YQFnJ77QQepAkt69JsN1OW9akBCsepOXERpShI3Hckvw92sGcx
ortAsrFbmbOjUOwukUwM1/o0O/lzgvGm+aM7mcyfQrd8jXWVQm9/cyhiEzx2sBXYkvb3AQq7nH0i
reqpeRaVeLSNnfsi/x8NIy/fIg015j79QOjM9G6QCMyH4a6FGJsmgbbWbxXHtaZOK9/FgOkHWLg+
wmpSS1c8Pb5C2CCsIfrtC7y69orhcGfKi49sCvA+CVIpektecD289Wnu7k1EQ9hWDeuHw03nde40
eIsaASKdpdlW3zrCvkG3RjVtgs6MLuQGMZ0yNDC5w5L4bgUo4EQ1L0n31aX0vh7B2DyteDYCQSl6
o0EZtjMjAtRkalyykJQvUoJQfSJNQe9JAeFIC+rNtIIKSC7DP44rbtGIO7rIz7ba3iLlex/9YbnQ
sufQVTAhBGfYqmSy5FdzHrHD7oLZdy2esd0F8EfB0wNY7Y+cDFtC6QYu/6EDhrV7kA2HsVH8DgDO
CQEHZU131eiLnQeYA5jMU1z6fmPnukfstV+DRM8IjY4Iyji6pMmpfg/ZR9ov7aVAmcGTC0icoeQ3
7ipqEUbXrFMEo3q2y9Kk95xkGA6lZkvfRhH6ettOtkRUHCyursvB8R5R4+IuLNMKhtPMq78l1zO1
gH/dNFrAs28xKbZhVRFzbQaKiohiyHuMbJnnVU50VMoRAC2albTpMB9dSO0PhVhel4Dy9pMggOCQ
t46VCgKYVlaT+9PVpD1Nz+vYN6r3Sp7w1cgjQjJTlNt4kYiMjocMcgufZL7+2ZK3fqccuz8LgnsB
OWIhBYsTyITk95YryYrYaesmG1ZJyWCpaRoeArZuPl7UufcdCNtpjFxH7dxafcUf58tK6CXX2V0t
3QFbD8GzpKTDJFg4WEI5uahQQIrOkO8KpJUYS6jH8NtOlcStfDpcTfciyz3tJvx1htY5g15lsgCT
4VA/WEyadOsP8nJENUqtS3Kg2+IPGBzW9bJ7E7a2IHfptCCAKEXZ4PTrEUTGxt1piEqLdkM/7Y3D
Ycxi/R+7h52JsoubRPxcXo+s1qFZR0Dd734Gspg4hF35s/z0K5uil1Cvs/Xh5rIiKQQsUto4kY0s
drw2ofyOLs0x8Or2qz2PzcA/GEYg6yvCd5HBG51iCGopsRaqUL8xnZ07edVK6hDSj12nBUFDwal1
F1K8KjsAvurPQonqogTy23xyzsbplQJk8rUOTU2fVTPg6lPyhCWLZURMsSLxmDvZYKchLwj7H9wx
fLAep/j1XZBzpG6X3UZ+CP29KTrcHraSwNnJnCYRP6EFBbFDE3iYWsn/pkloqO+jNqjCffI8UmAU
n3wzFBNhPXOGrwFDNwUprTrm7DkdMezQ66VWEAXg6cMoP9NhoCQm2mEMYPDADJriDgY8ltvtNtLP
nWnrIOZy0JvKoob0V2oHvcOqJgPkth4n++TK/gTnUu6lD0OuxPTVuePmdHsFMBJNJeGRqWhR+qY7
nn6SLvAhH2T5CfJtx1Mb/6VJFn2p/UL4vT4QsEVlJgGuDBNwJQRHR9Y2jdxdQJkLZzMJ2N4qqbtM
dQRmM/r7pFmtOPGeGkcrDG2V8/cuwG+EA8gPUiiLLKDD5vJga3cUFsLMwtgqgBsmeUMO0iOEdzd2
k/AYuyQLOUI+QTxW9CKsk7wgVZMp1t9gfjfbvDUbzHH1B6s9pMMBeRy8I1Nqw6WmbJA+oIYS/+Gi
vBMr6Ol7CkvT2zGopF7BvOU2dCfKsHNs52w7crT4651inPCrzmCW/w5kQHSuN66SH39N5855EmDy
rzYI5mAguvvZuyb7hf3JdaiLzUI2XZcl8rigYB8aYu8Q6Q2joZwhOOmsJIMb7HpCteyiJ9o1GLPb
1UC8yKNh6DTFKTddJp/0xnIkPM0SWpfN3WhCdVDH4B5Rm9JEefm5V+MqhKtogq7FS/19vkldRRRP
O/QDUF+SetRNwAsLcTkICcaBNtm03x2+01zJY+eb9nPlSBPbtipjHpdQcyJj4tjm1WB/1faO9jSO
AN6k+mUPxlvmFOvP6nj93vhOsVY2L5Zevs3+/xKHvuGFZvL63WcBNCaO+UCOQKYyHUwbBsAv/wpT
DD+lopvfefzl7z71venjBZGHPycr1mn+zW/h26apTG/7njk6H5p0pDJJORyU4F8ngLBpi4xONkit
g+/zP+a2+yg3qX0m4jGxvJ0gfj9Q6RDQ54kpmz1g5zUXsbneI8wCWMqLnrO5GGScH9cduMY4391Z
FoPlI0h392pA+FqxjCb/e7KoOEPkNiZHkvr+9QDYS1290hr8SIZBl/6bGK7ScnFEr3KzeKNVtaqo
DBSwx3zbPjbyK3ZL3cyJEBNsspbz4L7UewNDBf/eFq5OLe0BH/wRfjSkPWgXOqifGvIs/TxmWA3S
oSQxdujTnWa/qb5CY7Xk9ShY6PIS/cmXJwjTcd2GyZ3yVc8bcs9ZuthbOzEkueferre8FLiy9oHv
B7RzhxDUpEvv9xtgGZITXH2PwpaBIGgnqRz6gfY/d6aCL2rixA21wjRvO9UeZHLPhc3dHLB5AtKD
PrQUS7lJB9sIgYViWfl8ql33p3ALwqYRcVjLASwDQkYsdJD/7gCthdlzDcRWu+4w/lCxIeytgqS5
yIMwBQRDRpFbpgTEhx7Rh1+Ty2rLnbP8LXJfsE7a+S2dMbzwJFUTrrAqyXjzOIlniFx2NCDmyxNT
Q9REWmMkEwOYhh6rS5vhCrUki+nfzghIRXiNnTG/NrW4kr98BA3MO1J5qSIQyJmMAj7tZyfbtye1
TqjkeSDq3yDG7ext8R5GCKxQfO0biyWvHGoGJNDEcXlLgace1DVOX6ZG+SwRsCP5Q6hVSinrFYTE
l0DgZnJloecFocjfPAZrALTCurA8kB0rfaaVMry+EST2Vv80/lLCs2lJ1wujl2uqMFq3NJkq2hKx
ZJchhq1AFCHuPAjO/xR5d4tI+ECNNq8cDmVwZqWHhUfBB2Y8BxLW5mcAhJNpNcC3FwQZIX68X9a1
3s9iwuTi7+E2JwLPR7Q/Eq5BTjbVM/wwj6tUvF4BmABK29S/lomcoC1VapkjCbScb9jBAF/iDDYt
BoZxRhsGoJxOCl2hbDk/0nJIW8v3qr9RMps5iPN3WtDaoHESRV2WeIa7Vu4I05wM0bX//W2kMKvL
mvFcItjoSUphO82RScrAX4tD+WWWbO3Kv49hb+AqmpJ433DL4vH/XCIAaNmeNDaWFVgsWlI8pJhp
DHxjlShI64Auzz21uOvX4FvIBcLO8UCokYJsmnXe5ZYLDJGUrwd9uNVd5oqYiqUbqoGZfiAQ0Du8
DCzuEuYZ6sLmZpk4k+UhqgVBUETj81wbZx3bFyPRw2XrOgzHVOxJAhqh5fXrCT9MbyAtDxEWjsiG
9zI4U5xCRvW2+ccYvA2f0LhIVx8aaYL8Km8zp6ZsPtW+hRNbj3U/4yE2rDWCuDhupHPmGKd1FXGD
9NgaqNQnIy9wTDKHG2vDAxpaLp3NTgk/Atj2cpcxQ11Pe9bKd+vG2IKYog1j9RvyYZ+ZN5yeVPLk
4+Zy4MTaIHxnDPCG3GiHDc++04uuSDRQHCIZUYrlKx5Y8IZLOLc7BvXYyfr0qLSsfvVwqyh0mSY8
ab5vgPe3rZRxFGyU/98iBPwtwoQAB/+NDQA89aQXOr/Ng9kLQ0cxGJa6W8d+hdEEmagddfa3F8AW
kXxhlA8o8gziI41vjG8GbVupEty0+SHCGa8qoAOFXP24ivEd06/2xWH8MBuOs9vmb2PGBQ0jaoPz
J21LroYLP1o2rO6uoCGPmu1+rnlQ7k6+eyy0fW1Krop55YcitBPRFC2cqMeOCXGPRISTgFi+INsq
gFEFiyg2uRQOFkbz5YZ068oLsm7VF0pqGVZ4BP1pYqV3BhdfL44pLniNsLJsNCwqsX7WK3hBMow9
NlU0BTxI4V9sSt/dJHyksPierAgqfzhtQqq9IxoxD1obUgABy9gWeZ5JeKx499igGjnWTYb1d0MA
Ty8rGwsOa1bmGKEUlcsz2GtCRTlcnlI/0q5ba/MD4tlsHbxtH0P1RikDSKo065N1GFl1MgGgSfdG
CZBmcijuFj9CvrzU7jUTo7Py8sIg5O3Cm+levbtVGq6EtMkhYvJlzv4pa9LyEmC+yNVu3BaCgodD
LmlR4ogew28eRkjgOHqknL1GJQlB8hPewLwwd7++Ba1b+OKUCwo6n8FTFkLD1UDwJcjZGtdJMUDz
8T10dWyQwtte4glT3JCQkHOFsSVRwsgTV1Wx/y/i9BNT6SCf5w7tbrXZBNpXXDPd30lMRk+62jqA
SPGLHTmhJkju+ta/1GFNfb9js89tz0kGbqAln1ntYNxWcAm4XXP+UI8QuFQj1n0eQxeiKYMqYPFC
thG1S9rIwx779I18iknweXjAMhgg74bJHCZg9Cpf5lTsPtCLnaaNS5lupzT3DuqG3RycTfFUTPvw
hhFseHnmMwyFuqEBnGASm56eHMaPCYK15hryjyHx7UcCSsD6mvQxa4UNPQsuoaAfBISF/wJYwUIb
U73sJGaK3dvbbOaJ6QkYZTHWHAKkZdZcEsMh9f1jDkpQw9lC4+vB/5HQ8Vc5/QWoJNq1MiOm2TLd
gHYeqzSXpAe1HBgUft3zWGTRyFd5eE6YQqSfjG882UFh/ikUDpesb7oSEZ5Bi8Z2ZOnFFVbufX9K
ckhtrJlPsslxOabztkp99o7NQNlnT2pDm3Bfw2FSAp98pEB29+LAkznUTpkANvo4r2LUlJHiBD5a
y3JXnMk30rKk718kPSH+guYuyCRC5yN2derZdgPC9adrDoxSXXSkVjjMf8jTvSjQex3W/W5RJ1yx
hFw/u78WLt8orv4GKi77e8TtJMzhyPb7JPPArj+x/h4sxZHMWWAjMFZr6QUkovFyapAnVJiKx7i5
T9aP6EEuUMBFEud8Ix2xd2mVDZ3/N9qq6zCFB9+eTI5qLni8o2aRUKvfARjaaF0DrjVEXGq9tNAs
oXXPqonB1+8MdSQnBK0/GxlSr2iJZaxDFwU+QPQ48sGOqtLjA/c/PPykkESUyFapEzRFu+h0vmCI
Lc8pCcL2OknoRcBCAWiy/NFV36NgBqT1nDT9A4Bib7PT1YFc+AtsXsRGSBMYTJRg0CkCSrY6bxVq
JeBdf5paYoRnEixiSO4b3S1kuxcRvEwr34IVe78+1KvFYWDRTQEzGN3LQN/mlmRNo7D+tjiW0UfO
sJdFkkd9hS2BskdoW8xjCuiYeuphq5garNVKg3Xl3YmIzNkrDPfJTzYertCLNRmTla+oNkTLWRO/
ALCCWLk+DrOKAyoAV1PeEFFcwj+WaMz/sUMSWIYuTzvTZAVwaJaoTVTC0vr43PMzzWE5LUvr0wxE
NtOlkRq8Bw/+7e4a/SCgrbbpoaXAzX50HxaZ7yw/F06NXN0hVU8YcSuVqZpxbj5GnHELxK4L0QRs
we/YfPifd4mWzw1cBFPHvC5EBwFN2eRpUow70Pzfr9kcmEA2hh0BtVv5uLN+ES21c4aXI7zyyxwK
0CLNKWcZSuSv1W/J/qmiS4nu81PijNyCs8l0v9Ner4YChA5VPlgXUGqechE0GQtCQlR0T07QKOaM
la3vZ/S9yicN+wSflbhtzNDoWcB8AOkkal+zTPdo2P8uWb9nYE/MvX3360NJPkO2eBoeL33HAXqo
T2XkSNQ9+rX7h7wHQ91qDqYqbVXvjvlWOON9Dd0DHbApwLE84btaI3vjxWyl4+lqIUTSePIpn8DM
XaHVO1yPU4ZUx4xLpIEXpvcTLRyDBl0O3GDRxHz/+s6mmRiPhPfleTBIUX/VtU8m9HvZSsCXM5wV
F9cCt7lO/Zkvh5KQA/t7UOGU2+5/F9HS75XbIavYcViLrue1IozEJXk4q93/1chMzT3Igh5l7201
WupGK7u4+o4S/MRi+eVCDpb0FkNtCA22rnCZfGfk3XgV0moVdI1L0623FdDoLb+sHVGwElgK/+2X
mNUkcO6ZgsLapRNZSZPP+97GD6PTY8xqQzygo/FWFtejdZ3aKKmASTqNFAh1qrL8fU4+DqbBxPq3
9DgEcnaKzoBJ4ZrvkY8wyGRnALU5z8RyonfOCLjZ8pkFPMMS36PZBdCx8cZ5a7C3kczmDXXihRAs
XyQO+4NtoT7HWS54fIpJuh407bNwdvD6jRtCypNIHoMxo3LSf+cirBC5H2X8MwA+X9bf90aNfrSK
CBdXOSjNmKxs6pRAc/HZnCaLO2gk+8mObyhKzDGSjcY7seNrmHDFek5//8JIn8hCfK12SW/olwwf
jrLUTr9AmHGx8RUEmPK9YVzGlvDhs82AlA+FinApsskaA85bugQ0bP95UypF//09izpgv2ssRKh6
x4AZilqOgc7Gge6Klc+wpE820Z2ZokW0Uz39SL2Nk3Jtm781KB9ujtyGKaHnSi/W4WfSVWdWrYEZ
wis2w7AsducwGlpBlsmNp4mztm6CXs2FnP52bfP8f0ba4ELIbIHm537kllHEEe6YWNwvE1+GHSeH
YFr+Z6rag6kmiSRJoe0o2m+WZ8igRjdre2iIiR/3GaD05cpBu35VOXTxC1Jbj8DKSqkalpR8BEnb
vxW66w1d6WzjFBFyKXIrdNSvnYh7VjGO2XZK8uDnqvBC1e6srRiDo7niskzc6bgmIs4rfRe3Hsvp
Hx3kpgyVxJ+Olw6Z/45qYRDNi95eqo2S2v1xqi4QYAmAGew5qs1i8mVZYLIry0vvSs1y/AKDT5GZ
/85v9PvSSOGdZv8Y7qAmPVuMBNXL1h/JCw2ym0ueU2u2810uhOpkWt39fxZrH6ElFERLm6clYn6/
GmxBVHFeQtjg3y28GCGY9hB11V+zCZuH3N+nrq1Q+sl+k+USgaSHraGfq4oUfKz1E4yv9skborMv
hVJC0o9rIPUpnRJR7IjfxrbFtVbE1Y/3vIdvd0SW0DUiOo5R+zcTF+4bYij3Uge239A7hRIlYDxV
uDk3y0QLbC9zJlR3vj+wwY+Nno4ekiTB+uyLLHJmw5GeMS7Ii5tflcZD6wJGjCBcSKP0nUtN1YO3
pa28KHN+QqpHkWIIuM1X/yFOcs10H1VAuahpb9vKAbfhCCuKZdHOs6yF6l/OHLbSZgYBLyYWgdbS
TlkwA8HXhb+ZP/GZI6/LFFY0GXBjUrqj6m/FLDsXhzf/jfJ5/PZ88UcN89Pnp8C4cfkMeZJ2EZFC
EYqM+8QS/z6aJ13bMK4p7NsJarRbejQMFcmSEwPLp5wtWuBGa7JvdgBMs626E6n85MP0KlIwHega
evcI8Nof2n9sLMscmi+imh2skRC/zmWUte6TfKjVEos5uilhwdQGq5hLWHI44vRhrn4TadSVc4gV
LS/aVsGHhS/Fk60I2w5gXXaOS1724f/Pz87JAdgcPYTcr2Oysj76u16EK/c4+SCyb+5t0Lvwmzmp
su6xn9gRogo0clnpNhWpOctsfLhrhOYejb414dfs1wY5rL7dM9LIIVnkO/NGRyhYnpNXjIgGX98J
CkFy2HFzyi0+RLWBj2ivMmI66tE4rlYuPTabItYNmfOxssmdWPx5jxEe8FGHa0y49YuRPUHcQPdx
b6ZN8OoW7zAK8kHISaV0ftzXLf8p60yQBuG0dRk+OipLgMKGPVZIi3akz/mj6I/wN8e//dRyd2db
02h4AFMM8Fh6AMa3jytZZvapETXNx5WrFNXJS7IE+ttNotDjQhakkzfVtYMJLtPJGAIq4Uh4GNlr
jc/k+Ym2nhj5grDelE3FMLJKCbd0XfSOF4wsonSWQ9y5AfCuwn7Pe1syPtx6AsSWFzC9lEylE/ec
z4Es3o8oDZPi4bdOHybBjFPKFeeaK7NMNgdXpgWzJAt/DNVjd6FTRD4Osb5Z9cmjEXnsYY4YAJyM
RNjd13+9xY+Dhbw5ISk66Wh6ItqwcFmdgrD3AjGdaokvTRIm4DxNQiIFo/Gp734g/21NhoN1sVTG
+12cv38BQx/bCew3L3Fds/+K5O9WMRbk12OYFvQgK8CzUWOrLbCjVIxh2D+b8oBS2bwqFvVWNLR9
Z96LbNUyqhJqZ0Tc7ta/1iHYy/H7FJQiln7zXeo21YyBw0e0CKCPH/FecqJVR1fiXWD9g70nXQdw
lgW5PCgqttuZXL2EeVxtTCIxDOptJXycjJUruyePQBAJvcsc/92zJQvvsEQcxkX44hL0KG99ADJ2
U6/7ipiDPAzY/8I1143MiDcB2vOacwZNFJQ9aWVcDQ2rtTkq0ulpqN/SuS9uuVi5sr++d9J7Vaxj
p/OR5OS14xQdurU2SwdoVR+5XSLfz2oI8Cv3e3IaHtCZkytYkaUdGxrYWRoLYljc8dKvbrIbTKvx
b/TSU4i5ucWOfa2JQzLHaMdrtO4IeG9eFQT++RciVap0I0dfmv8xAoRByPbsIVTPtc9gi+j/BDMn
wCrKyL7FULzSj/q1GPw5EZw2BgKotgdGP7crj8E4eu1Mk84t/WUwsT18sheCnfH2rNDg44d04DZB
hzvk394+GfqyGui5LlPjBHbH8vdyRloKQtwJaJoS9QlKrMWR8CJRIjFAfNqSy9GVSc+BEFez+DKY
PvB/8D+mkc8tgsl6f+PtjNy0pabqxvRSapx7b2Kium6AvH/KcOb65kAlb/nnbIemngx6Lg3+Fp7n
CrcyFySsXPJS2w/eZZ2oY8oCJNNYBbG07H1BvJSvsa/2oZ8iO91EFt5BGGu6MADouz6kKkjjBbid
+QGZeSyebUneNGcqWQhfkBEfPrTv5KI6ecL/+n5WwPK8OFL0IC64ApgSsqV+3gM1Xad/7TgMJME6
KnNvxQ4VUe0ALCDHzxQhy81UCt+A5NLPgO6dUmXJC4PIcvMs22QMkGwmLJxRZ2QiDTlkQs095zS9
ONMGHIbTr/SEflyVQet6lztDgiI6UZLXoriXu0l9sTmbJW/Zw7iZp6P0Fmm5KoXWnMTBlVAqWhcE
QdNwM17pY4Pqvl8pNDaHpHjfrncTT98775K/1VPNJv4gBtZG38qYjkniB8dLQHug3aXHTqd3BblC
geHU20OE/pLLlhvDLhLQG+1T61/IGNZ78r4VUwws+NrzrZkLVYVeVFCkFED1hqMMAEx2EgYhoZ+9
bGqBJsYhyfgU6lOTUSHSGqOk+VdfxsJYjqZU+vDhXN7NUz6wQW92Tf/WGURQD0Bq7AETHhpTi/Ke
ShFJU4wkRuSMgSW2YDVn39JSCfaF8R5Ko6jMQAiEb9Tn+l3yva8nX4UCZOfyf3QdGBeB5nm/GPQ0
RHhV37l/dYKlJoiQWm+PcSSJiCDV1lgJZvSbDfX2r1hjciehkdgWO19yyHMEDsNzxoVSenNyg8Hx
O9DBBQUNGWyuvg29CzlpwXYGzggY4IfYCbEI3KjAIh6F9xbinOBD9pHHiHGkoF7Ha0yTGaR4O2uZ
kWwVdCDxpQwrQwAdSEqvpHLMlqXZXGZaGq8+XmtLOEZ/0+k57h3FxcgrkMolccpEkXfJowtcPVp9
ubnFpkt5hrl1eUTxXo2t1H7eEigRx9rSVxYhBbhem8mlfXfl2V5C5eXTYIlZ8aJtyphw4Vv70OGX
uLpw49JPQOtJYrm+KFBU64/DpwXLCGI/Tz8YKDcuzcLW+PQyPCWPEe142bOtMlmw3FlY47tCuSCT
3aPDcb0eKOlilYhYXNEZ3vBg9AU3QLyGT1r0Bz8XO05J8EbHdF9XOgXD5ZCcpUy6j0LHGJowhh6z
siI86i4daMngiangBNcZrSuCZvuJfveLThhM85NYDKGhoYXv2Qizablesvsdgio2DmyBSVUDNoS+
F8sdN4ujBQdFQEKyITGxxJy1pP/3BmJK9CyKD4nP3NPqMLaOKqbOn5X9qyxJ5Tfqefnm5AXb+eyB
MWP6QedEtKYikwdBNPwKsSqkMu7UGtoGz51/2mnJ219Ga2oiKr0BLSSDM6k4cUBN49QF/saavIVo
bAEbMzLygyIcG5VxwJMLPVD0CT42UGVsBZPRVnSex2TeIBXbJbeaWqtIAGL8ya7vAZ7RMeaxBMwV
yjIsjIzO9gkr0EfxK4iq0NIIquVUBhkKFugjjut+U8g+GJo5l1Tx+7jnfk6vHlVTTusIFHgXjyJv
/nsXLjpQRPA8zq2dqVj8gUUJxxCMLF8LFbVsdsCZDQauVn/emI0HJBlbkNbRVDdRd64pD9qAapw6
mNtnxqRtNadNoi0dWIaoYFmW5cSxFdz1pZXeLoOI8O0KmzE3/8jB1lEwuSh9MpPlAGBW6l//XndC
hDxhmW6xoAj/HYiwk8/jrzBj3jm3goPoxZkLM46fQbrL7hNw1yafmZB583hG0onrh2OhnlIIIVuI
iAevh+TfY76dgCqKuHKavPXEGBU27qbMltc2D5bMA+OWxRtrHnUkS8aZkaoE+dcJbFCM+hPr+v0Q
VhayB4HSW93von9mtllusBsM1S4GX6a4/XWpNfAeZmeXYjs1Ogv2SltTKUsgV7VIHqg3ECyng3qo
KnFXBgT2USxcbDUpOWzqP9j9A0Lixl5yTBNRJxwaGRcoiEU4G5a06WH48jLLq/oLbwF+CDRMe9EP
ug6eX7hgnS2sY7eM4MsxnZ4jw0c4+7KJ3OTtGhk1/Z/O28iGuSFwHf3znOB7pk0zn14je7z0LoZW
3iwkYwItWE499lIEnIFijQzv414psF+RcXVt8GjS0Nw5Xa19Fu0uPX/IO6D2CU549s0Hx+tfN9yA
rdX9hKpK/g9Uby87SC+7wur4Yn8MihLDFkQU95L6IS77z2ZBnf467nVt+o7vOlah60fpJXjj8zfv
T41v1l/sLV4JO4/TjEDsRZZUBSzs8Aob9VVM+go7qrL6+eB4RsryNEYoODYGjYGFmmSdKN1oSePJ
agYYnNBxXhLRpDiYx+xySg2/Z6grogtOwD2yY+aW77z9WlBXEwtkWYC6+iS/HKIj6P10s5D5pcFQ
3AjpsGXUNmzK7Nukg9AGJXno2EcVE4/Ph37ZDxPg+G+bQqo5Cgz6rGwNcxA6xzsvBKt+CXM54f6y
H8sDEjERNIMRZ+cfLAZSs4/49iU4vedtaJR6jBTXySsOztGh89lBEmx/MvtCcMA9BZTy6EciH9m7
vaKnDVBnnm55UOBjQM+UUal4ei0FoTi2r2bEggNmxqh2wMnhgEkJUuzjH9OXvXE3tS8ekp3VjPPD
A3YVPMXxfhfruUZADvLVdEviCK1jcDrizrV8WXbQbPihi9PO6dL/YD5c4kj5yj03ic+AErBwFXO7
OaxBLnrjIkleqafvHh4/LBXB6BEcnXxsmzqIJdvc9eaG57DL+OxJsQq++igjkBmn13fmoR04TCzn
Qbb727FqPXc1lswDJS9IDHrBx6OeCXtMy+DwniC0/AAyPwnFPPqRu7t/jnKu9jzUsSOcn5JF63R4
bHFxHoUkNouGZWR+7I+tKTYqAYullFDEu7/TDr45HcR+2UkJ/qjXD/WkzjgXSuNNmV/QUaX/Onh/
+1ZonTfZVdoCJzq/f2XT3oLaQhsRG1afcD0PwyAG1/ITGkdqduqwu/bsJ9cINAo3gqA8/LhTCoR/
LdINMgaG8G1pfyuIkNeQtCPTqf9GeBgdi6JG1lPrD+fKYsV4mBJcAn3XuGe9ItiEyVHaTapiWKrg
Ihxr5ab0j0E9XBOHaonLBWHnp27f7H7mgYhb0Gt/tlDg3iqc/9XYBJ28+XnqbVu6HbIo44n//b32
ttddDnofoVW7vKQj6WcalmpR7rY21kUrW4+Qz6rSSqVUmiPY+EiLKvKFYgC1Ui4r9oXlGHlTfvY6
Qzrg5nbaAYMMhemrGCVIAQWGiK0/CX0Rp8f6mnQoxKrtVzhyGv3cFiDbOxnnXu9Mggtenj7goHXf
0vpp48qCg9S5TIOCeCz3Y91rUrDkgxb6tmeW4fpfsPc/S6a8QJ90mXxoE8CnwkYbDtvM2m+k8bOb
4BKAaYuFuk4yTR3Rkur3zxe+Fc9cd6yRuB72ZiVcV8ZAvytfA3kaN0eb8UcZWjYFNUW/lIbxLK4W
HBeOM4sMRoG6RQbXZ4JKbVn28QsFKXxNpzUX6U55bWusB58n8cr5tXMRL9Re5UWc8GfWxkrIWcZB
5koWFDqwWgILgL+ltNlFkldRImWWoE1x7pk2SU4RxZ3//f/0WS6PuZmxNuOIuZdkjZexHckCrnbE
sD4/hScQCiECn+WcMKoCvHA1JnZH5FFNssyIDdJ1pv1GhnhaNolZO/vX1EqcKu1zsowtBgcahzlP
HrZwRWoL9/+eIGZ4xeZ9CgprqY9BPrAcFcudTs5JIwQH82tXGPSciPbszU2G4yFnXu+HqGVTVJ4V
vMwEA0Zg5kISSFX27+yDQqpYDahnNAbZT31tUUP+/EqsAT2NyLQ5DSQCh/1JcrFjA9819yFWnVwA
c31pHNsr5eb+HV5dlKMUe9L/9mCZp1+a2B3AUMA7X7nIk0tUS+47Kgmp93CixBU2SVjgdJtaLpfE
ws1Bw99YWJx4QqcJ58KYcMuU9iJuJUjLAfhm8xqckCrjs9YRd7I7P9qHjgfwuLygJvz2tNoH7tSe
H/86l5NTz2d3Q1+uR9RVx5ix+lnNUt6jiz3k+WGu9nTDKzHF5195GL9J/LZGYPZrcapn6wKc8Urk
1R7h3d/EJz/0Ro+dsGlKNJ6k8hjTEs8kcKvFQw3P3N2eeSwCPFdnbd5m1iSFRs/YuabqJZ+chaIK
FviboO8GKhtXGJh8PejVpUzS9T8DfkRm+9zjWOUXTZcRfz/mLAf2EJg87qSyBiWbaPOitTYflL/k
JZ/N2+wmdIXOwSkVTLBkum1RB/nbBgEd7ZeuaywIiyBWmGQPQ8k0GvzuvsSosy6U7rD0kP7HDN/G
N25Qenfpb7hI+ANrFFy+I+Z6uQlj4FyZu1PzhQG8AkzHZ3zNzAw48i+vRsrR72KaIi0ZLc79oB8L
fix8ySoG8YxMWg6zswq9e/OxhYks/Oy5X7a6B6YwMOe4fdpfW2I9bcmun7udSQCV1UjKfmiNQwG3
cB/ddiFrvrQbqYoAwNJzGdxHWAaXHctfgfeQPVBVt5I1i2Rh9zojuM/HZ9WwNDF5RVEr6Fdu0amu
9fXzGVRXlg6bcTzF4wdPGahEyXfCSn1rhO5MwND7hB79oijO6vbA4POnhgXdJfIYFc47LiH5nXOr
0cDBToGw8mteeLaQdrM7WFcoWItzs3VTo+kynjXLwz+NOwcXqeSs8+v8x0xiNQ1q7tA50obtujbR
lyTlTLO89lt8Li+2evxBT83Y5+gWROcpmy0AwwRPCOXzieHeG7iTTERsLjpd9vdDRynXYvQBZAsy
RVujSkwgbVcav2kRkjH0ivKVPhmSbsW++4PVcGs5nb7LKxaqj4JFMBF7RUhyLv6fzm/6Mkk0aJ2x
yfI79GFmZEEToiPpmWOvqg1mg5R1YR9Tpy3j+cjpxgKqndNxrUfKD9SWx/Pim+zKYt8dEGie9K5R
3uhkab3lRgrNHFwKfAybI5zYAoP7LGoqCpkNmrgGWhg4H3wo+IWj/Xfjxf9N0Qy+QYiIuKlKp2hr
6wyv+a7IqneDvFpRWZNgBsIFKXSIv5pxsROFwVf+UDakaXzZEZbM4uBr7HpKe3rIug6wx9nPxD89
10BHGP+KXjbk3pR8GbGiHMOmiTLNFFylZmcDqeu98xk4sp2nVICbykbls08qUVePAvTZ7Y8dFXub
z1Zw+93bhG0OqqCrXgYk+Ub8BRHbYudhmO1vdKEunIxtxp5FuNEvpmvHCt/M/dqy2v5kfDexNnV9
in8KwViHMJrEUa3g7uxIPm1S4WRBP59QHbCJCzYPHR4KFXx0vyeixwQoQEa/WtpXZxprpprIoSY4
sVf0Hwffcjtdlhl2YPmN5SyzeFkyL57mMaqkslkaDyvpmlxP6DNkfPEclUOI+kzTLQYrvGlBlbLY
q6IEY3KFbMawjsxu8DtNNS3w6OD+hrfRM7bBGSoyRjj/Ucw/nz34yKHilE5GxK9EMI7j1AwQbjHr
uqSeKZ3t6RXVUviY5JTfAd11P7y3xIsM8HwJwmirEPLVnhcRj9YsIxDbH4nqn3MaqPWBb7n7qcl7
pNylDBafwagIb/gXx8SIH+q/R5Ggl+yEzmElbCgbGnnnQ9ZHg1AYDuE/2+A96vwKzRIj2qt+HJPm
+BVGVT6loSU6emcvhYbUnvrWsbMm1FRif4wEkf04Dv7I7T2mwRonOkqumCOcBqdFlMfldUEp4gBT
Wt5XiKM/fYW0ioQBqLLegZ4n8bG+MBOOiSW7BV8B7/9ZZ0Q+vxKqGduwv5KwNyeJcyZmqaN/Kz2R
0HSRpVr7+1zKEExvGQwfRHyP/TdfWeln9CFbwMRWiEMcpzlFX9AhfVhiWh3vpOrXGhoTtwM/pdRg
2PqLhUon9zd8HHVa2fpDrCiRARvqOkQ+m6bZg6vhukPuj93LzIjrpS4b6D/Hw9kE5f1BWTnWRYTu
9OwZiSv0xo00i6+mP2Fe3BixG2GbUnIEfGRxfGIDBU70H9C8U8UqPCaP8rx6djMmnOk5sIbOdo0x
TPhrXczVFRqajwAj/M9VnJKb34sg0eE69W4ZRXJz5nqV8BfSZ2SIUmjAXZe7urZfOwJ2ytPpGF/K
J5TDgGnFbM/aEs/3dphCHa+y/48jS9Ei7Ehe836Wlh4YLAjImjdwrb4KUQxsiHATBp8b1TSpMAZA
PCM58fbdmBiiBTaZ02BOKcbNRORwpuIXzQTmdAjfdEFuMNaRIRc9eb0YUHbpmyGCAtzdU4MfvYZY
Zb+MRgBQHRV5w3cgh+aYppFQQFRoYT/wyMRkOMMGFvjc9TEYGBBUvrQnot+yyWQPdKvLPGbBHrol
j1iyY2Qc/XgnqAX0xBrZoz8jyEydqJpMqmXxBUeJz/1Rc8zh9tgJqffzDQVwU5/69JWvF4oBpDxb
Lm6sXMyaBNgSy6Oq4qpD6EsU2uaV+hU/EnOLfWvvJFG0mY2jA+9brnkXWOV1eOmBVyq4HAOYuzf5
G4+arBHk+Hs2TSIGMKZK3sCDKEoQFmuoKa8VeqO8G50xKhsEqvwYQQC/CR8sVM7eoSyKIpcfXWk2
PLJFdsbN7J45hNDd/5v83fswOkL0Y50EVbzHBKrk+eY0RJabtn+IzO7FOm9igQtwlQV/BVZBlz4N
P+LrB18vDYp4GWoDphBUxMCQVOW4bNN/d47Im+sRCfz6611pOP2Z2+n+RTlZgpWCKomQc1gxn/7x
o2zINgoPhAeY0Z8P/QMmRypFjT3yZNNBcSf2ZoMPhnoWBBb4RHIYmHPzm45XMupZ3IxmddRO6zcy
UOMWWiBtUJbM6atb0Ws/SW6wFYBClEtcJfeNQYtSg+XTVQ+NyBn1E4cGLgGKRi4FzLpxF8ydeHjq
pCJ0NJyCyeKzTOgS0ZTB/vgxfeFndM44cbAoSl1hOy5PnCuTCyiyJ62kA44vsk4BbfAGfWlPQyH3
oeFzcxFPeSucF3A++sWn7eifollXGaZoRUsYUEPVysqUA243BnEb/0/XbfuwthCJE7ta2h/Sg1rg
da6Ghx5uHDepY8kETJOxUN6aajg19PUl6bBqsUayt7Ibat4yOAAjpXMgKDmBLnfs7eM9QYcv8WE0
4nCsvoQJzxJ06aCslgdmmNXc0pPxQLobYVNkHlK2ALNOoVA+H+zdZqtgwL2PHBdhMyD7KwAPdnkM
ylZOirT6KQZ7XjUb1x4UN8ooBx/Mn0c+ZR5cvcNn9wHTpvLntQLzVkjnEtIaBenzLEPWRHxW9fSR
xB2ZF6sSS396CYluzXqHsv/2e1EpVMbRFlp399CYZI8m/KoE2JeHX6diAZbJ9RJPABR7dJ//CPLB
avHLCD7iLTeId7ulA5g7qtOjZndRePfZRGb3CH0Jm/hdGvZMKPLXXFjJ2AfKL6KvVxB7Irnm6EZe
muh4eVIim+cHf/9ebP//nxIptXrePnWiImmeJ+ds0OiwiPdG4k6v7f+6gWCPMvg9X3hGW4mPR84U
4FmHx8fi6XCedvgOQW0dLfqpgyaN/WYwZaQ8ZBSxuunzUv6mwcMs1psisRc8T+UHZvNqsbrw46ve
X1efCWzNRB0b4beHyg2FYfP0vtid2dfHHduu6iuxdkOgpg1agONUjqw0WGnJ3iQoLfcm1Mqq9puP
OdY+OhU0EVyLg7yIFqIKFfw6TRZlBrrAttnUpGLLr31kKkHJ1DEabj5XS9RLT+fIaZ04t8aHhDpq
cAgevS4UJuIXsHff5zqfKGGVbMOo7tcBeTpsc6vPasDmZyNFDHzwqLs1wMr6xOpS38oGArdod0Wd
SASLuHko28w6xUfO+c+YB3/CPjoNs4XO6wUncf8VZTY5ekg2v+Shd2y5UzgxJmab0ZWq5/CRQaOX
9YMWQvZ0b0m+Dsh4uP8NmeDmK/qcsmmgAyswR9N9sVG253gUfRgyij2IkY9Iq746w6fTmuMVGfF8
2aQnaxw3vFgw1YA3XUAX+QESfeyhsMPOkC/6CVjknuR8iFpO0M+bQcQuyvAMsP2iCLLHmtiO1Eut
tfhy+7hguTYl7a3266D2AS+9QhwNOuQPw4IEoSHP2i0WAFQUf4w/auj0Dzy1mjCjwTI80vRXncGb
8zYAdKXBOUojyx5gCqrouX2If4OGFQ3JqQ7y5CdJAvfhp4pDtgeGqHI14L0Mbgc7QIG0e+6+jvBC
ZKmewg+V1iZw9oN4Phn/iFzcRU5FJbc2Beh/SXKuuIyeuOYugJFDm1XZUiAXWz9klNaeUvVx31Ox
DoAtGUMJCQ4Vr2m4ZPr6sXTyjTRSkzPWtx5pdzrWfBSHL7zAv8LoQc7LPOP67s/qJuy1lWRBzauS
3KnQBRHeHqDr6Ae0ZETvqHew5ZZflZlnMgNYn8HVnAihbhKXMPjIxlqMRAEeUj4CX3vo4LTftLfO
m5FmgQsGiFVx5DlYLdYJWqxEbjlEMQb5LEF2sgfMHVqCXBQD7bpG2JRvsJVY9Iq59IxRAN0vtaJX
5q7cN6Egiw3kL2d0JFnqHI6OG8cGYY+9/r3/0feXF7/Rrj2qidLUdAAYmZP5aLF0mnLEf5D7edAg
Uv/cac6Szsqc27wi1g/KPMHEaUgACvjjyGvYFHr1cdbbuvvvnhnqV1jf6GO8/QImnMVPM2VxeCL6
VL6VoNO8NdxcvztcKBNCcViqKGPtPFNDt+oMLi/SYPjaNrOLWAnRI1u8sLlfe6ihhkxx3n565w5u
ZHdwPccHfa+YDdCuZwgoC087h3dBh4qurNP3efHdysFVEgywq0/f8HZNUftfUKPqN5tO8Gna7u+T
g+gcJkvQbsYwnpml86jO3SOyaObqzc4CNE3yR1xG9oWlXfi2orVoCfHBW98z/XCgvwVY59tR+8Wi
TMlpWfpra7TM0XMvXDkEkE4pRh5s8KDlSxdFUOT7a56enLJir7vSp/g9tHC+ldT6yr/TCIGdTmd5
UdKyTQ9hPccpKlB2rW/HYGuMl1mqZx1nEQUo+MD7/RUbCPt8FpyH/4ld1P8Dhgt+6k0zFHMdX3xV
iAmgqzi8WHuihlkSrvO4vo6diOWyRRH0pw0a6TeE1xQy5ykXRMt4X4L7rq9JDP908HuHxvMo5Fbw
PNMmrdldVZHV6ljCY2bXXeu/o7ao/4a5KrhuxIFJTkEcUP5O1v0QTCixHRse6KwlZba/jkMpS0s8
ajcUe8ypea70xh45Ep2aFJ+JXtcM0glvClTp3jxO5nx6br1FVFa+rM6hklmEspWzGpw20MKVrpQk
97W5A00QY06Hl8GPKpylD0qT8wuYUYq3AZ2/V9J7GXoPncI0qUNLcpEcapW4sv8mrxxPAql7C/5/
BYH2lrZpBFurB/mtHcxgMaEr0ziQmOokyXvhyLJGyI+zl2P/rfAdJ83nrriOP31oV9Gg5IuLjDFV
rmUdRrApY4eRuLk8FaRIzHdr35+rs0PRN3IhfNUYPQ46PtS4tKHb1WLUMVmHQcswCgNXtUfVlaL+
aTvzJhCkut1pcuGcc8P9NkdORL5zGMg1AqtR5RR5j8SfPGxBm6tMPyUQxBKAhC1B52+k8FJpw4ft
N3CtjrCMwlxA4ngM/zJgy0TEypQV/RbNJwkoJQ7ZALqxdNH0gaeMBo6L7487H5/qlen5MZgwkmfH
Sq8t3iwDyh8oTkvvwlbdUNHwxyBsrX+/tNfXzEYHMfBqnh/Sau6OOfpJvKyDcToRgHb4ldbs9j1b
Jziwt8Fbt/e4Bejbv8KIzTkW5woIFwhOh70Lf81K66sZTp/sda3/ChDrLCc3IFbuVw8WI58Jiy/B
WXfBlz/6trMfMflrqXIOVpHSuWBWVUvLgh0glJK61UnbmgaQMvRqehhf8IfKScL4HY4uVpu2xqAa
h8Bwqar1Ut8whgUS7T9NIk1cO6pWUP3gsk5bb3jUacEhAHzBem8X0D+uEjzH0Y51eQEjvzWg6h4p
M97BDbQd64M8Y2I3CqEwc7GRvUhM9z4vbyzlpi/OCg9LwPOeGEHqzwToOvcxJd4Fuj/9fEy3VhIc
OSBNAdQ39s0vi5wF5uv6XXa2WQW2Zxvm1egwfn7tlhzIp38zHBkJ4daUsQAJZA9eCy+rfQdIpxRJ
Gtj84WXhh+3lQEOjD38ndSkc0fpwsHQJ+MB1x8mEzabvAG/TxXmvOauFAABuer6fh9JlevO7rx6T
Gj83ejvvUqrGXjJBelqtZTGkYolYL+3o1CdgZYh6NLEoW31CiIlg9P+McwoYcgetlsKDQqFQd9KR
MHeQ05akyzMyQKqcuY+mTcUIMsSYrgyYnRr526z3dSS34FyHu3eFqeavUCGO7KAH/NG0ZwEoxghJ
Hg6vyQI1ZteC1VKcHaflnY3LYp8wVwya+aJIlWiWCxURWk2A19YrnvEvnzkviwWEhmNcH9Zl4XMv
+zwgCezOLx+WdownvRAj3HfFV9xaOBqichxLSW8tDsbSPhAW7Vlej0+y73ts48qrNuI8FVc7AsvS
/Kt74ma99mMAEsWJKmNFfTTKrOGXYcPZZr/vfE/Fa1xzI3HYvwbMdOCsLqTFPVroUUzpophCKxaP
V8CcChP/3Dw8mjBc6IYB3uxEs5H5QD+lCc9tkvoBhALDCq1mpscZtcgL6fPZb9FztbqzhlYVoy42
u8OEe/Ze9oqUp7lIoQz1BlYoP5Yw7YDYNLG823f34NF5EcdinWdfYIZivVAsqv7s5P6u3RP4YeWb
RvXtdbBlL1Djr264Q8TtE3z9GD6szGiTKVUaGpyAeOvJlFzxxTHRyz1EjlFTJaqgPXcFnIlWPbvd
xtd5+vIvVn9os1wp2IN0xEY4tnBX1Mjb+jtlyFVcdrlbtv8dgpaKl+uYPfer/qG6Ppqyp5HEeiyA
FGQT3jEsDPUa4mkVR/XoiuiEi7uTIQiMz3sGXayyLArM1RTx6yKXyuVq7TZopIrsWrSsEFZ/t5uA
LNdVaU2vFsq5/jW/MOdjNXxuCqchfN9AO6D3Bdhz1i/KlAYLPFnhb0ttb/jgjxxPTseG5dmEotQg
W6dMgQjNiMfXROmptNg+vDjPqkhZ1xIGiy+mD7lBVIkQOaLNNZxRgxn52lZTO+9sAK4jET0lTtT7
g253eaTebyrzF7jX3IE/kTA1mFJkmPxygRqmJhCLCdXy0qlW+AaTrNz04VvY3JaFVSFgWBg0m7uk
YneLWIio8bbTWWiwrOkv4wPG43jABQyXciMVJ2pR6HSXgoqFqohN9ApC/wfnSYJVrbZqYCG663fy
pWrPuVx4qfl+l67CxnV4WMtgrM8sm/bIBOtlXupZy50u5IC4+ajePGNZioP9w+bXbOg7ptK6UFjC
ifsCg2vOdnd1jEvdEI/pUVS+38FS7CPyLpOqBuRKALpOT7X2NEU0y7IvbVcIy0tB5Xw4bmnlonHE
pt4IiX9yLNLjOhl89yTCE0+rsNKOciNa6sJAa0467PLFdDADqkSWJMSdKk5c6pSsyQZDk7kVKPrF
PEZGx7bq/k+iZjmmloykrBOwDnYDtFGZ4VjcFeqv1jHXU8sLHg8OzJ8tlxn8pKgTcb/APoFokf5Z
sjE+zETdSh+LNgEbTPtqI8Uo2RaWnXt4mtjhHy9QhWimXOay3ze31PY3jYnk8Rfe9beHRNjOTSbH
NlXqMSusSlwI1d7C61KY4wic7GqUxNjYh/nDIXr/ZUMg1qOp+mWEOX52R9MSJr+HPkYPJWZDaRSj
CfUV2bj0cuM04ZlnsoVgo5YoaUItE4yiWoZUV8rWJqX67247NPNk/D7JeQesCoJ8S6WS2GPkfIRS
VTNBWVcK+7HarbWWxkpyfZYpHbEBbMmvD+VPLA/181gS9uoWXCLTmB8hjHsvq/I68cAgMjicpHPD
9koIFv9+NXdJZaIIh0v6sEP6AZ8u4qabs9sEIDlKAx+CPtJDf6siif3B+NGKqv8Ork1g4x5WOTQU
wdGQphNUY85BwjoQkOh/f0WaeQ1rheWiGUtHhqI5saG/jrAb8Zzqdx03H15Pw9xILfop2VJ7GTjS
cgsoU/3JpDBrNCX8KUZiBCyDQlbyKnucetbK9FT5/ajVYg27tHfgpYLqaKNUre/iqOTvQE6oOoKi
sFwH6XP7KPsMxXSyilsw2brWE7WQ41Jzbty5FftcFHRA0imkqC4JPwl6AxOcts8SUdQsqxabi9ze
LG9kiM6Sn214vdzr27/PS+4ginGYzOpIjIlw1JtyHlm0rSxCFtKWebGWINMVLRrsLWakjZ6LSU5B
PGMcSMp1oDKoRY9DarME5hnwVES0KrY7fURvOLS8k+A4z8tfgAli4MvT3H34kP2VRk89Crvc8Fhx
OYCK1iTsRuPcHJbMv/v6KawZovuwrV7BdY9JuOwCqn3Zl8fCuwcchC5gZe2cFlCbkmBuPTp+mJQN
8tjPJhmfrzSeGG6s7O5EpxJAZ792Cri0MFzAYdPTgbD0tsRf6gXWB7Tnvd53rFJvgt4/9f4AKDuj
VuQ3hIOoByDpXXJfVwEKXaKAqC1gmCApA08i+v4dgfE8gEiAY+LtUQETbCCfGqzfnkVrNIeK/mxI
A+bkDQk+k7+4CmPMxN7aDQ1MKMlQ2cK87E1BpZzitbPNKCbVGrkiXal8mE/Dh2FF4aADX1B4R0/8
KL37Epkq/9nNOjh+hULMDBkaoOayRMZPJlCjYSqfaDEFuj/jQbzlLXYXOQdl40TrUQH1L3i+xvGL
7/4pYfUlPD4Wm+M8jPelixuhQjsT6GetmgKXCJHMv/A9q/JDe+3+wNDL7zorM25Ejy52GgmPWJfR
6/gV2+QlSmwekV+YZN1ERg44u8NG6fHjVMKwNkizto7zrSU2ppXctP4T7xfhVkbNvw3JbIsVIH9T
5CxULomadlie9HBgYbRbxfMbUZ8Wm/yXoYnqnXGywbNINvA4UDlRJ6F7wsTiWbeltBpEUkbry0pE
pjr/Lglcb0cpgNDKt/OR/EurNfPUWcJQbn2oHcJHuVELeTqSeXSVLx/dGldjLrdIGmg4od/kjzEm
m0722hGETS9Jy8EzWLvwQhDHgc6cVfBuPlOv4sms6EueGeNWp6YcWCThnaiHinkO8mNFHGGUopv0
/bXfLloZGBCtKPlc0TU+2oouQkh2Ur31+sEWLzHdQr5mOpc7ahE0SGzXCHbhP3gjUrjQeg47bbvZ
mUtwxOLssjo8DdbxurQRTHdmS2VVVhzqCDrmx2U7Kvsuxe674fBBiit8X6x9WKTN7q2eW5TIQkBJ
QOu3ydbvCJV+6DNH2D3aYBKUIX+jiFo0plbdFFoLJR5P4AhTlm7OCGertZpRIIqwRYErKKgYN5qg
pG3SbcRjvnAgjBj9YF3pXIB/dkzrGEhcLvnlFgJy84kg3davaGkfbEJU07VIqjwd9SAD4Ngsubmp
jKuSprwDP03Il6zOHqZL0IaAkuKj+hjs08IjqipqdSIs3QzXHP27BqOgvpdPCelQwu52f7H900rG
QS9NBg8Dc+pIZSu4I7RPH5Rc9fbMoPfu+rNIlPrQiphbndtm70nfue9SDgryPBGORZKWE8PZs9ih
guK2eeF2ZV47OOFEOxghwgNmrTmNm3mCy5wm3dYhUblXi+CY0Gei9/F1IQHf6I8JW7Y8dyvpSqWZ
M1YpJk0r4iF6/XBskB+19uSCGUY+5RXRmlOfX6QvTqVV6MfDTblPZQcamvADdJMiVpZ/3upzspJY
r3KvqzhQs0VmFDk5HK7aPejz2S/lnen+xVecKE8hJOjcwZ+x33vV8xHfya4470SThoRz59UJlAoQ
21ah7MlLmAfZdlHjhCMTHkusDQr0/J9BIBvK+6ZBk1u9d+uFt+cqCXIT6UzOeVvexOWLuGBuIkrL
R+QUqIjNQ5W9o8KLrk4s5mTJ3zfs5Qb7Jp/MOalGYq10hDpqH2tffrSbS4r53fphupJx4lORRffU
TeBqgOEGRUQxY37EnaYm0xTMz+2+dhJlkHKRq/VvUPx2+5YfudIoWxx0Sn3HZEV1BcfEu8Lo5KKs
6LO9YsLO9vs0QyQTVOoelGaRthbPZTm/bUn1cMGjt9Qo7t9kgHJYJekWUYujf57UOr381v8tqE85
kmt9n71mDimIZU7lERsBkkSM1/+1NZIt6dXh/Ne1/VycOBDhAei3nGqcFuqI2G2aUo4VfuTI2Ifh
Ry3RlF78HeHcuXKlItsDJhFfflp2rHEsH2l0ncOssfmaE+lX4OS6ERvi2SVLSKi0Je7FXF5F2lOS
oCvEKGekzCFgFGy4Twb/4z4QVaEmfqq4GA38aOKKp2BeXO9FKFa/PpHduqM1nesoXwjSlp5s1JDI
AZWNPfEbPZL2r4PFFJkGHlBAr1SM4y7kvmzu/stkdFxV8LERo1COm+MVhGcTtuKY/mxJn9q0EBYI
Wjsdj0ls0F4dpjK4srTMLnYEzQlxDic4QUpCWRiZsy+IwBiw4XQTjNyPuc8rc5ssFNcloXJZJ6T4
BojmVo/3C+bHVpN1UHAs2mhcZFL46hNmQvxuKr/4tBYqHmcXCh3x/mQIEJMVN+AhymLV9h6JLkkO
v8YK8KCyZH2qUNLTJQlSYG05Ow/mlpz15F+0vwkLOeLZ0Zgy84kJF6EMk+/WTn6dpYJJwo9j4nig
ucDAzpHl63jrZejSivHUPhEioFlHlmo0xmLDSiO7oMj2GHbMo+BV725otEMQsWoEaVyNykfXHnSM
HvLIWXYwWgIK+o/Xpc2JlQDJuXJevMoy/d5LXspdCccIpdELXZqXrfteSUrapCKSoN/UWxEJhYVn
c7e82khijBlgdUf6pbFGb1JY+Ox28sjyHpS4ZMxa9Dg+4nnhYn2GJEVTtt4C+EiXHPqfTSqTCiWy
uBQgzTnM+zAB9SdN0zQBLAkE8oiAaxtKBSc7n84x5ZJnuzp1qie222RsMy5HKe7U571xELCZw1Bl
gnq5VHt93adSElgPG5GEfe8FZmOC5coAnGMhshTjc3M1tmAtqSSdZab8IJLkYQyt0FiCancgTUBl
EiVG/+gkhm2+ZBsrz8IW9cDuoH+bRAsXYdXA1W0o1S/0qnVfcPKsldBBDPy2CRtUUh88Kbu/42vr
AzYbB9BIfbK9UGvQdCnHj3yGwBzfjbPKNPVhIgjgFogNa/7Palg8pcvRF+mnMTIADp4eBcgIFPGk
3mtNJ6kkidNoGTBQ4klp1+mdKTZxF1SrAHLjTiSxT28Gxk7zMZYM0yqY1Ha+9BVMmu+R90f/yMXU
MBS16ws2388ytroUO+zVRk1fhKu9x6RYtu/PBZfkYtzPs5GJqMz3C6Hqmt9PL5cyiKHzhgqi++jX
upllyQJXjcpEfdfSgH4YFMx9ldeyyaIZkqHbHTAZkqW3MQkw6PynRwBXAAQ5XlsSCBHCYe64id2b
rOYAP/93rfJ4CW4uk+LhH+QFP1BAyYguaPDFEDv9bFvYirYT9g0q36Lyoi7/D7xzxTfIIGP+nMg6
DbkLVT+9bRNZNtc9J7FKGPsUpUTOkbvTBjOUbTadeHW9VQVW4D2LBXXow5xKLTjIn9C+/cvHN28W
lMZRo8jva15jKvDRhJ+ZEpUUm4i4H8lXx5+pk1HSzXdB+mvq+NkS2Wgq52WAIzufKto8+/l6NRsv
fcHxTVxTRml0C6wSnyUcjKiL424ltH8kglnILYxQ09lbglzfTgBnK8v3BATVOyIYVxi9T/qx/oDG
8dihXaOMRED2ZhdwqGvOVVTP6vCGKI/BNP5zWUYJuyhO3pIpDFJr8M0iQr6YwWG+xeBFpKGfMXs6
wyfe4r7tN+4hU0ZzRMZtzj7p0091c2tJzpPvaAQA4tF3hOfq5J9EE5HNhnc26WBk037K8WCaH9gV
5l7g7AyT5c2repNZdjmlvS3fraXCrSFuF3mwKM4GIcixQkzCbqhdeUoG/YkjhAkJNNvCWja6wpNo
C+XM/mrHrg/Swh6mKkUH4UT6dKQwPBa6/awSqBYu7YBESOG4h/0oLeJflj9VYvq8CWAIITSzlFh1
BZN5SSmW4yyeMHtzaAo2NgUFD/2AUzRxx4qgUNKHDOvU1kQVmghxzmzZzjnLtf8j43tqvzXsJ5Oy
bGiTLVBJrZmwMjG82Jisngc9HkClNtbZuu2oZPj0kxQW3nnU95AvNOjFJRJ7GYiixKwgbzPFx/7l
avA84/TYzT0IfSeVwjYxtKR645WKqL0KpxAcsjIdhQG0fvi1w1kToGBsLUdnph2Yn7VYAifjket1
+RSq6J8sN/E5OruLhYHnJJ7s01AOnTK0UlzBHUub9y9gmJON3nYVLKKIq2VKXHlCNeKE6vAKTBk8
WIYOMR1SSai3GjGRPcHLOoJ7nW234mRJLdALE+qNZvnI1+Zr4WtFrIg/aQ8K7OMd+REzCvYhZcOn
G1Wz3ktkOH/EHfapizadCP4AoDrktayjsNKcPaEua0vPpzEuGZIgHmRx+Ti4eQdhiFyaAbebYM9/
AcCKiH3B6tv/fKtyTQAKNL96F5D54hYGk02NxJs9MEmDoEjOUrS6hQ1yDzRM3CDqiuPckKN/xrgL
k0PPGpG9pm8DAwUd7i4hrbIez6E9YzRALkEOfr2JckriOgorBhNmU8PY/PTh9617R2JthRcWZRV1
dcwgvBAP2ZIhWiXjtrZKlQ+WShfKILmsxuCP7pS0iaKWqav0QYoiteTUumN6H9lNImghSFJBOaKM
ChUI54ZunMtkBGMyzy1DvQlN2rfhOgw6WB5uFqPKgyEoJpcLkUaRUfx44U/FuvwrU8J8jDqXuIvD
wSmrsoD5yXkAaeymkv1uhxq+sRh78mnRPG8PBUs7tbWJvHca09A+IUaa6GdbeNUKyvrfsrAMkNK4
feUL8ytn8CTGtoEQ4viJkVubkCqH4ElIhix2CunXIP1PRmCBpkuyRJ45gBtIhRlyT/hqLbNEZHun
FAYvKDpH8tV9rM6kZEQalrQDw4TUk4tr0WCWJWHTdVIFim+5DuvPxz1XFZypWJiy7XduDgdLjSR7
OLqRXvDK5ij4JHPYHG5yWLHOFYlq4RHosw34A4FX7FqdlAs8ayHvUezhBcTLJ8A2X2XTW1xkwpPc
+lUq8S/bkbK6c0X6ANkbtvpzxa9oCsrSAJ/PgDKQCQa+GqFgk7JSv9XU6UTMTCvqx34I89K++g2r
6O8T60F40+aBfMDa+/0o55njnnn7DHvejre/UtxLR3FZJcJQ37xEMh4DCNI/iZy/i6s0neuqz/dx
vEU2me4WXqd2oZ3azuhhxXAJ+Gw3S572vCIyNPDhNp95nGG9va19oljE7YutIkSg+rIosyeVjZnq
jHw4oW2WX3kXlAjDeOY9T26qAPKzxlxm1b2w/2bI6iRzREfSeIjeHhNWqm/Xh13CYiUgeNDxwwWa
aKhhdBcLgOeBFEmFNQ+ayoz+pA74Vuq4OMSroQBK60uTH1lDU80omCpwo6mCTLy8e5r3mUdhxLyy
9gaQX3/OJzw+yP/+rYgwksU2vWd5Rohv638JQdWPfPVCd28VSJRMbriWV9rENCx6j4fhZWvYnJl2
o1AzlMNN9ufdsTGS1svE4mQklaMuMjUGsceE40qih7Blb/TSd2eZuN8LZ/VcbItBPGoFBB38GxBd
E7nj2/gF7SadqFFDURnNzhWFZHt0dnYNA7qLT5SbWB1wOyxVra7AgL320xHKfQHdKhh6EMxgJkGI
K6OdNEtos5/cvuAZuUjwokGZZ9wVJ8ObzQYcQ6YImynJM3+FZcnZSCyAWt9o9q14wI5nnm+v9ItR
W1QfMaTpRjv4+V48CBXjrfivs/dDWBlEhq7vaMTIk7LVCizRD7/QnIWr2HSNZM3S88SGaAiKP7pu
La7bAElRXHWgU0i5WiArOfHBYe1UUsJmIpw6A4N6BGdPn1bdela6Ck1Fj9BncWRLFEQyx3CaWBrX
1rR3YQ1GVAT95iGPRN9bOpmvK0Tv12thl2gjjVrmklBl5qMlHEj91sBc4SV/Qr7lnA14MvYFW2b/
HjHV1s/AwuU3Y6jUIzDemouDSCGrYSQjCNGPpj88A5C/opt7jgTs8Cjvg/1oZYgGdYTpjLpAbef3
eiilu/1RZYqdvgQTsJ8gTwhHtjttgu66hxz366OAfANUcg8CHm8+tTUKu/j1OPEEFeH1JvjqNfax
c2qRMjtf9aBR5H+372GWuXaDMg1zCvPeXRtZD7MAWyuauK4+LzilO/R0jdk5c9+o8JwHl1xuvIfb
LIf6ibuHl8Ysat0+dzAOhaqXUkfYZYrlR9+QE1vpXnQhPQ27TQh5jsa73wKeRESbvl2chhBW+H+M
EGu5mwhnivPNFr26O/bkZttLMPEOgYV5YWNIc9Fnpt76FNROzpR/Kiw0SsDjw4O25IJhvE4VdJqg
U6GHVjoHAdu/bWrRq3mvTGBcuVz1E6pAchHgVm/4DOFgk0FQoW7b89r0XTMWYK6dzXvyt879BeoB
Jd/dLlcALq548K50OutXZaXNZaGG5/RuGHDWpOeEqLH+mgY/TjlYFChbjPimlW1hK/+ms5lgOxIS
wKqvsTpXLrj6dhYW7YjqtG3CzwIbjNiAphDa2LFSzk5DQqWWoJnsEnOEygxZZ4bzQqx7AIyO4NOs
P3NDWE1RwpKTogiE/cs2RnHVvAbUMZxLrDkqdIvAWsh0VgtI2MXHoluL0wtI+O28sESYeK9B84HG
taLXJBIs7UTOflwAnNFfK//waf15c6DMfjKCZCB0dsRf72mw3a3Ek3YVM+jZijBj4skYpLt66Pvl
AP1yTCVJq4tfwnH2WXfled5Nyn6JeRT1pIvk9shBwFIsmNeC++gSpsWg7LK7eeC/+F+O0sxMqQnz
Yx85zLaDraWgdB1Qynmo6KLwW3WdXBwWz5pqDMT0J7HBvvfvg85sz+OyDeVsKgZ8wAYLw5cokbcU
vvLAmTa+dWHOT+0213ow5FsNkZtijnd65DtqHDTafzC02rGTdop2y/ZBXGs+Jdy6zEYb82X1tMw0
lihTZqvNu33sb8w5ZAjlRr1kXWJuid6Z8ZVMyMSitQx4Q9lrf3PeKCXDH3NSqNXEZzsY942qCnla
L7oizBo6+VLN88jLJDvZ6qbElvZN7L3VOm113zT6HmMknEYoMpvq9Rxnw2JsQSqoFN2887/exhbm
CK66xYwRqwkBtpQcpx3ySkl072WAUeXxKyf0sk5Qv2FyothGox+NhtG4RnmF1OnhnVvsyXDXnud7
8Pkb5Yz82fdY6HgO2BwPF5yPcRuDwNC4h/2Il44qOpHVooZ6vRi1oHRml/TN66c/7McKhbna/kJD
kDK6Mze4eu0VhYIWYl9SJIC7h9NNbpNawuY2fXteQvBYXx9U9YD21T+s1htEEkkonosW1SfIPD1+
1TvVyYKsPBMUJdq86SjPaFeZqP06yPAxUUoJqzqP66C/1ql6fPATz1v8pYOTp3yjFoFKjOc0DYcl
95JfAQioWhxTd1ciwRp1c5bKWTQL5ysDPblY39a7LDI4UEoFQdHbVpQG9KXOb8NtToGKQPkLbsK7
jklR+CLGeOQNe14NXbd6l9qjaU63wa0H/PBqlbXRU2HC7NL6UyFmrreA8yN+qFrjf6TLd5GuIa3R
3YBPcZen1s+54yovEKnY8n6c8WWNOn1c8/IGyZPGstB00fVmfmHhBGfM4GwyoWVGzM4AZO3Za0EW
1rdt9pOhqbPuQVCvfvBCkhDw5zDLX0dqGljBxdo+YXLnO9m7F1EwDFrMgc1TFxcgl1lpxvB1SfBT
5OjAF2i5U1Uech6DjJFJ2cEh6bLUv3AlCWVuVkuzErsMIB3DWqCT1Sb6yLf6FPhgqH0H3vUJtMTo
/ohVTRaYIgo8pB/UwyDS2Fbcx7jvVJSFf8ZrkxPVjwvkKnVfdQUEfNcwFzMUqRbzUrcJffAtWiVD
mv7OfBAoa0OAjGl8epm+mIwaItZ+5SRUaXWSsFchTGJ294XWPy8pyMu/dPW0tjhkd8yBzkIqxj9b
hqF9O9HVu6ai5RrMOuANfAVcVk2Yg1FQqao0nMPc6nrk6aPwIwKMzzy4P8/4fejg3mTIW+f0QhG7
fw5BGkSDyVUaM7kzfEoRMz6JLL5HWgwaorTm/Lt+hTVKaixRv4mvZwZ+Omr3hxwIql9NhC5hOByj
MIpWGbqKbMJIpiqUws9w7aRV98xKZ+gb2UcNg9f54q0SgERNWZf5IQebRmWIXDvDdwiaRu/mBPZz
zj9cG2KRyLn8pHiX57xQ1xumRU5ol7WZ0Fi5jjsV9BWDvr41lPXmdYuuxfSlxvkatkReT8Lq9T6r
KoZFk/w0ZJ4J286NfpdNtAsdx/pHISyJ+YFV1/CLALJuQzT63Wym/IuCc+7k/Br5Vf/Vkiwi6UzG
KiFUCYzY7ZZvEAcVh3PueNbTd7K17M7rwWEsX0dGJ9G1J9gI2UxnKWEkWxv40EBTT5SXrL6epV8r
6XlC12qnOWVslvI4e8+8aHno8mX2MamRZcnitYKFFdXwh3eSNAlumbMp8IaQDapK+82ZKcEoFxtV
NHOjz5gx7zdwlbxqEexcl/AX7GX3cOiyi6LPzkJWNQLPTZ9Mx/lpYq7UX/J9+s8twqMdK+NSK0ul
AmiCN1MoQqNRkwovoG/dO6eiIs+T0mezI59G/2O2MRBOhXi2OwZdEjWJNZ6YqBi4d+YX7oWbgEPG
Szqaz8tFHJbdMTZCGpuk3c/IPdtkNaQdyh1mE6wUk5Yqr56UaQdSXPqaL5IrH5zIJYWWWzB9iSBs
dvJudzYghPuhdyXIzRdpFRAjfw8HShmnRRxhP4EhVwI4s5K8zUh4RLih6F5BMaOqSNoHodu4tr4F
A5HrMaQuaLATAAu2+kfTlDBDUkkxePJJPAJrWWWvZhKQTjVnBRjpJ8gcsvbnruQXaGeugDqVpLVr
hwBn4HTl7JX5/GV55oC6FeDfEjF/2ctPtBHgBXk+aPobn4nqxAi52IJkEA2dk4RknmYA0bjlHVYB
2o3a8l1QUnHaj/w0k58QqPpX3N4Q7Io0cWfUh51zvnDFSCOMR5dZlaUdZU4/EY2/YB8LY4NV7UjZ
zwrHk2ZYIV215UUqTENv1kWu52NGWA8uG85EZCka61/3LMXMiFA/7yXO05cWyTUVgNf3WeN/Agc5
0yZKLg2I6rYRD6ZtAh7yuZZaeMbqmXZVTNttdt1u85ktENZ9YK1XiMXUy5pwTAd0Km4HNqxN1SM7
9v0WyX7rF1YP/QV41VVkfTqGJ1TO4WmemKxtQcpErOjKX1KWBk90LQW5PhXq1lLNlHoI+D8h3W4P
D6JSeQ3kk4dqVdbLAHP/rALUmEOwRxuq1nEj84372cx5DFigWmx0itb1VrUOympkUurI3smnlost
dmvAQk5H/BvAr3pyFCMIgkPemMa8y6zIxcWqCzPCuWwuTEfb4nT4helzMKizstVAqQhkMbDdPj1e
1cO1FyQHyI/OMCmI4rAB8nos0T77RIWxGLgEEm0ybt3cccPfYQz6wYL58nBRx8iwaCJfQQXzWyi0
94eiygRQYF8Kmg9MF6U/aacWI7CG44EGbzhDETQnAhYEpHD9e34voEbxhUfSB33/hGg569mbxMss
PRXkmA2siIOXTGmGsGBTIJz4ZnTid3p9580oh4/fjHYCUwaa0BTQSYehzUat56/7vl/rE4HTvJ9H
wE1bnx7RQTfOAl1maI2Dl+wgG7q8wjIfWOZ93/kl+PTaEDUFJAzhnBqkY/fpF9qZkK9+cTpg/kI1
RzCc8CXyAVQC0Y9N8Z84fFx8vsBPkHyCKIIYcm2biCKy/ln25ZwFUbeRzamwis0nHkGvlyhD1dTN
x8QoyBXMhbSx8IUUa9UGbjLlE9wwje7Zah9DwiJ/tE94pOe9ObCG4ANx/FroZKxlzzCogUfRh5Te
6G1RwzUKRH8KvMzn2rf56fp90uVr/wvzTxFMDRI3jhQ3tBcj162N5wMo4zQG1DonQVUV/wPWORR7
9MdreDu5dkhSBFIT1sh9deoe0h4doytv6141UWYWLQhBRrw3XepYFeRazJlcCgrz7njFu5l9bT9k
EnwKBTQqHVQQlOpGHgX+M4nfG+HlGK5di2f+LsZK9CA5QVO7/dpk71y3oPiU6bJcwujGDhtGMMjC
H8fDo332zy0euEu5QRbuYMDSckiMxIfpSScJhsxqP4n5fKFCnFg5rOLWdYKxZDW1aDdvzgdxssfr
4bx59Sphc8I51jpQoKGsVRZBton3SWPuV+zzKWZbiXdAiaHQt3SMt84FKCb79pRNJKlCPAPZeDWW
hPUIFkWfpvAqKbWWwpQVPsIF4nZC0IkH0iDBx54+uTY6996Jb1NwrFQH+z0Yrv1ln5ODVfLlJ3Ub
tr8KcjnQHPOQamIGSfaZkxEUDFe1uoCUGlCYa5cFsNkLwz16J0fGLauBQ8pXnA5VBpjTsCizG94l
Grl8qSQ/dbBTZP+kC67lSsnQezV7S1iHcE1r6t//ns539TITv0B3wC/b16LeqIMkk4DIs1WPkkcg
Z/czmriyb8gquT0RKyT54Gw9fjh0I+vbHLSzBOWd1kSy3/27ncYMPt2xDBV1j+BBsH99dykVPYz+
ewxPpS2DRGOesJjvf+ze/xnEik3FK6m+eS0HTy4QGVQ7FxcX4/OfF+kSqiWcimoUYdQeNnYeAK4r
1RpHn5tl8yHBBIWyk5f6f1ZnjudIA65/VSxcritgDgvEN9BxBC91nXR3DMBvOmzoCvUmbPD0NkO6
CAYLbpUEurYBvtY5GUrO6F6hjynQatIHHOi5sEwERW/53hKCM/j+Y6TOlbaI7dh0PfkkJ3j/5otM
IjzBci52lCJJV4/qTUCVPl/uonXknN4syGnQswG0vGIfXbL+q1F0NowMjGlz8vwzTAmWPaYARfUx
Kmm61I71BsZ4E4GD8MDaFspJfkx9dqeNcVJuU8jR6TmpbXmqU3cX4ZY+ZReox2+RzlO9Sw7O3Hwc
v16HDhGukRmVImzfctgi7syOsMbzd3IjV8sh9zxsNAdfT2rnLf+MFYIFcwvLI4p6VZzFtG7Ph7fC
vK3UIfSBF6hNhjMkxZab7XcGBricdBLvHr2kbbHkNDXQiZ0og78B+BI/pi70P8CCUjPO47yjZpFL
msRt1ZQgKh4ExnbNoSOYbzX1/qXIMT2gv8ankg0D1rX4TuutM7iJuXf5uAOR5Kycycc8oGwewzKt
FdIwZTZmGIV7UG3Y2dxwO1g/pWrr4qG7RjQ8BnkhvLPgRVpOQJbPVtCytxV/FNiqSUzSu2VuUggP
xpJVf6cmgGOgL3wQJI2V/wrrnRbjiqjersAOkYhuqKHIIDJFYZAdHFDbiGVhsM1TyqOZ4cv/9nhD
nEdbrxdjIOrYHCqS3K552WHJbH77LNl3Dd1Nq0NMxiDPQ881Ip2FAqwYY/zRZNoITlRsssn4vqns
yMSq6WqqcZswzq1fdMGZeu7DUj5jZEOPddS1ZnBlxfZJ6op4rX1A++z961Vlrm4YGDgIPxudgEme
iZmO9FAD8c1I3R19mYLS+WWZdJt2pZQRpcmWPPPgW9116nXr/Pr+g61h31t3Jga13pnbO7kpoJTH
PBmH3C3nVOze4BuoDYpyzfTUxwBbdzOZRNIwa0Bt3OAELSDHEMwwHDgU9R855JHALpDLImdjFc7F
GGOf6Dsz7NalNL710qvt6ElEO4bpBseGvPAAMXp9/7wVCABm9xGfDZZz44Mz8SpZ/Pb8lLHi9TqD
rwB84bA01l0eJdkTJq3KLH78dwh3aqNThtls4QQA7PMwt932ZEIoD7FzLVMsXq68z5MKMG4nhgoq
4at33jzCs4uFuInvf38DBm8t73P+ZydX1qv8kACC6eSfAwlPHIkYghSYfUdESB6JBjFG0LaI66Nz
wERnCidxw3Z9tdNhDBDqaO76evMRqjkbMl6/f/EC9MOF0B6PoUmqsYtuH41hZPx3oI3AZ2h/XeWl
59JWaKwVuMoZka42obFw9FsGTIk7rksgQLWMcJV/WHmqwxFFUNIqkJdqoE0nbVpNJ+Ck+9HlCBp6
XfuPGW6Ya5gvJj3Amzk31aB3KppMZDciTDvEWwfmkaBYWxmIIyK2SPxYxIDvWajlNMGfBKJMOQzv
jEs4NkeYOvmgT9v3ZmBimKYne2Mti6+LzBercWLNfFvQ2fBCxn5E7gzIid5HXPlMjebErqtN8PxT
r9IMuGEcwWTmJHsSht3zvpw9qJlZ4cE3lqKrGes86eNqWaVaNx8T2BE6HAsjqfx6GWQYgyRImZWR
01gqfVzfR5PAzEsacAjuZR21Y+Am59hsDGnH5MTs4kWH2hGnS9g8kjzITrBHNy2N9StovW6M7SXz
0nKPBfLnjDQtRRSyZEWzKPvY7Af51KOYfSwqIysWysXFIL243JAqnSoTG2VzbaK4OnXyOhlulVgI
p1ncvO9XmgDPBrkiY6kukNi7kYjKlRQEug+d46xd8VdNbxFvulq+O+j2SW0PXRBpqzPYyRRpuDyD
x7197CZo6WRKKjj0W4nkek6ULrLcgMvOA3I8E0kB/DD2CkcOdkRUfUuBXYd0ToKVdAlqm5sfuI1k
aIk6dF9ZCm+oQ9VGRQuisM2iRcXvKf5d5uHT+M45AfwdzymUrZm0AoVd/dA1jAW6BJgH3KUmhhAc
DwIZM7GiHZTOO+AS4cDjfxv3UtHZsXBAWVIq0+ssOUXsIbRnxHfWEu3N97Bk73EvI6YzccVfnH3K
KTxvyxzOqLHUdVG28HaPGPkl3u4/nWjKd7kQySbEGfUvXYSSGnZ5ZpaPfelGPpGCC8Q1zZyyl5EE
daUGldt4QvI30nEMPB+Orc5Yfvm4iV/tcNY8v75Q/E5Glgu47WNGU79bkOUZHM40M3h86UUegsn+
6YxKu9jOwbj4tZkfM/4PrQf6unWDlPWVw97T3z8gkkVKZXl9N++tut8gjaRnSrLbnaccRDqrKKLl
bRMviWNXLN0PN98dBWcn+wgwflrejpGC7KDO/EPhjZ2mKWSB8k9g3Tv+fJVQFDGqeLoNGs4P1YRx
68UkP1FgqbdyrpR0s2YU5eiVrdm2a+NUAeS7G9HPcQENMVYMcPRTle5PW1p/3fKc7TvLZHZNfnaW
eEDo47wU7hJ6G8Oo0zf+KbJfbEaEaGa9zoH7YkXc2mo/xJ5UE3y2e6fcFXS3xMmLVmk27rsYnwtL
wiKKMN9q9/GLJrRUXs4l3uAZrVIZUsrE4OyXule2cvI1pakuwo+f0YXap3G/oq8fr9v+IOcECYa3
0fPU+Q3+/x9eECm/tiBufX9zeohd8yi/yGYG9ez4gSibT8NCjREkjYIDfa26zSCAB5qh5ZPFOeSW
JDQs0oZeWPuQ28oqgo2tbVbr2uB1bhYO9wPuE/+iNVbJ93fu6gefhmY4tVnkQgzCWRdVbCk6VoUi
LjoBMkZD8DK6bTKQKvgXtOB9GUrOFBJD+9osd0uOIOxaqXPldcUTAyovLVCJcH4wTm1GQf5LW2a8
SyVYBt2O8eTcAc9oVTRC/iDs9G51JDSrO8CXb5GEWswViCT37WNAzGaDZCVQsfKExcvM72ljXHLS
j9bdVgTM6up4v/Isgb8cemwXrw2V3iTv+PPM7D8ygGW1YnIi6FwCr4M2oDQ/yQEkohEeRXoJWkOf
0vTEdMvrnXg1nJOgNu6u8DKOTiOcDo5mUVUPNWL5KGbXzrzw7jtbnOcAvh+j1Anpvf4jGNKCjdEf
3GdvOY2cSL7WNXBnHSWMvVjE0tal6jLbyTCRnp6NX9/VcHhGNOJaXDrXY1bNMMAQdxQPlNKuyNgT
s7xyhZyE539aHRWigSAYuF70LpmR7jTkDNzbvCugbNzbHUPGgzr+6av2Uv8AVyPIxoCumeboflJB
S0gvSlFBAGzc8MgBxRv8QjYTblEBI/Cxmt2f5k7tAW03qhl8shUr3fzMjyEhAHJYMu3VM4ZfCF8f
q/XUtffFtWGRNIhzeoA5XOCCgeUgA2LK4epWgtKU7ZFXrKByFTgMQW0iVWojFsI/DIdIQLXXopcD
amGDllBDd2cjrv67rbb5I8Qr5dLsZbspQDfl532dG0yd46/j83p8Z7tCjjcdi7CQgmnGgNd2qlH0
vWyP4Vmp/+QqUYYQxnWhGkzLrXglcD5ih7TDDzniDkvk7vspzm/+9jRqoHqo+butmJ99TZNq3eSU
rsxgICauDEJwYsIUlypDJffFhNq12gxEDSJ5vGidf/DClSOu8WOUW7YQQO/t5Rc/vv/fz6U2vUqZ
kioE5wdlmlu6Gjmht+3knONA6dng6AAzB/Z4IHNzY8UIee7BQiSdG9RkQOBcZN1MMY43nJNQt/LK
afCbweofWhZiRTwXNaUQqHBsCg2XJEOpvh2gF0X/Z1U7BfQl1GCZK5h/kLfq/sB5ZAtx3/ccOkMQ
ag/z/F69UethJ8+2jThXUAnaVCY9UPJwo3mAoSCVSz2QXeBi6GzD6jogsHLCghHTL2cJI8UwhLRv
pjlqGOP62edjqczd+wQmXiTmwlZBmS20UdcaAgUsdUgrMyQI5Bgj9U9chO5CSlsWW9lvFVv6wc0c
bbsSh8sJItRpo72jtv4+Rhnx9l2/Y7+sI31DJa8OUFES1aa3AG9ZkicPf5r0Xe/+R8V9zSyo7W5V
Fr5hwCCNDLZ55CZByfLOW7cy33LG72J2btp3SLg08f4gtTBlRVreIBok2cFdmTo2RNjppiw1hesV
f8v6nKPmhD0Q/aGolbIn9IOBRtQqJ0YKH4ICPHuPuO5g421uv878AqbjUwHdlFmcwLbl7Or880ga
0DfdaubY1nzz8AgB6eqzK0hSC2a7Lxk/bdfIh3OmQREioWt59hRyBnxp4aaPcMXnSW2kpkFu72if
AiPVjoYjGqP5ugvNIbQIGoZi/Pj3yMnWLzFrVSJbkfMTGt+EX7sh6upGftgW54D7QK7Mz7MM3Goh
fHuGd/Vn7ceXLxdITlXmCihR7mluLh7PzSe82gqrzqVJ/j/THw+UcP1kfFRdVqIzO0iIbbT5O0lQ
4yo1cZ6VkhyTVicuAJOs72onlXbIy1MnRCwpF7XEWl+QD0kLOqypFM5kgxyR2YIZlxu8Rqmrq8xL
Bfc2nMRu5vbPY2fqPwGzCbwetoclbkbFCcFX4caGmUdtkMzWKqDQ0xvYvrAGzk7MQeY+rVIx6C5Z
U7DBSa/4A9EGsaeV7wS0Rwes6rZIygrDck47fAcZOrwjBcihNY9wLWKPW9fOzuoxkL79C43fwoc7
ABd9JaEN8sqdGKVM1rVBFNGCeMqhDX9dpk5gPYmEe/PAnuSRDQBg2vfOuXLFrll70FuTKRtOSemx
XAz6BBk9qHLx0CDj5kZIr1MrXlNWNvyDMolFvbI0wtaf1vZ6wo9HyTTlEfEoi5krsgKCMms64arU
Z8XiEIR6KEPnr5sRk7FdRDJAJfAO9MtWqGCPugQ9NI/hTmBwjwLAEFLch0JsX2EpNLljfe1uVP/k
HR9tsxveTI4d8Ue5UUdo6BfMTZkP24zj1PVtTH8cp+lDsq6mmnjy3imLB5c+MBY019q4T4wTOyrT
jRQroiYGDaBBC7eotNhN71vcRR2RCpOOFjhXqZwukoHRYaTRc44N3zqZflySTVzNj/qO+U/cv+eU
980MZz0d/KC+sdvRMm4l88AYFT5KKMLXmrlXZQY8WPeYpmr+DECq4w39/1dV/5sB9jqPpqz8XhOj
72nXI9UTKm5Jc7i1+Oz/44SHnFgvPDF7MVA8OiMFQtj/caygUuRk1yhuNp1FzRHNdZ8++ZJ4wvTh
Lko3lQiHTstG41RGnHxcFP454OZ54oo4LbvvPB+Ia9x2v7Mwyps2pApnjhQoe8ywQDJVo/AJytqe
IEZVWmONnL5wI6C6HzUzoKyCn1LB4BZJ3kaOrye+O5ovlFMNC/iglQtfRJGzxy6oRwmOi3qYE9Mm
8cr3SZw9IETIpEB+Fg8qzgZv5oIXx8unpKMRmp3xCZptjcPBQSERL8VsrE2VLiYNo+K4zpvgaK0C
OO1RkTQsi1+6hr+uc/EN/sqs12/nOYaKrh9bATI9pbeeV2qjBUbZPZ3CY6MYEyjsbERIeIkGZ8ML
e6R8bnRHkn9thufk66hzh2TElqrxPWaGZxGFj+fTw8oBQ/bSBnJEKN/7SyLI4SYOzYRw2URA7Rlc
PU9nh/WR1IDwmaUPRV4Vu76xJCkM4X1rlbkprIFZzmN6EHJ7FiR57IqYD+3EOM+zWkbinZRK06My
GJwOibfhH3tpAmhkDYuywK9LLKdMyL+tj032226v53m8okj9cqGkG2lLFZOt4t06Xc0KPsVjDQap
n7Ixhsc5xhPbe1tJ1HsYWvAhtgu7RsWG9JPJ8mjtIIaTT7S+tbGJeFa6cywlpC+EOg89SKCtCWiv
sBdBNiU7/j6HHLCdOPSApyaj9B/ata+2oexwf1HU3ikFJNmDrOJ+xZJw7UKiJ8j0bpDQ7yQvr4O7
2Gxh4E3ECGdDAvCTf7QpLhq7/woYbIkgO9BK89xLwfEYv4w5NRbL81010STVDMJT7k+T2Lwy3WLO
h8sraB5pxnLOTrzPs6dfBvBaDbjVegync26vFZNCTCNVY+3tFBP4jQLA9i61qjdQlocBAUnyCurh
cAVIuMSCVd0GjrV4rYNTeChjRY4JoTk4YjQlz0wdjfBCuhofAa7gq4VViJPo3kmG3bMEo/BGtxNV
+eJHmJD+oqqyM4EuAiXxQmuKfMc/dbCPXItWOeooaa4KYIE+OKcajGGenvPsqXJ8GN3ijpVHPT3q
2BiUpH4JtW4jbNI43KQPcQ68D5i8reOry6UeuYNMnKLRzTEbNK1BR3nHxJqYH/kB/aXuCmSeAdcg
gs1zSWf0Lj/qnbUG2waaxgU8VwiNmqH/xpLdJ7T8itU4cBLw9RGVDbJ/uzxE2ed0VY86X+B8m1Va
qZIJS+K7/G9AvDddyCLQNyszSuw44Yz1X/iWmRTYErCzspqePTzr/19Qx6obQS4DCWUc0zgA9fIz
qqzJKlsZYLZYPxML5HuOUy5B2ZuI7cNzvHQGgOWRsmZHRjlStB+mkPTn73F+uyNDZqYcs0EdZmEf
aDQ1UcIO+3I4PH55Z64KXbZfRnmbdk06YxyoT+L3XHaLjI/uzTNRXHUrn5M7Izsjc6UuxfNw3QTi
eKYIQYDeNngeyNw2/uoh46LkrjYzrKzZQLSd3ghUFLzptpNA9pNNsYuP/HLkNIUABY8YdfBUGfjK
ucnlWd5/QQwPLGngyZi4IVq9VKYD4FSjwico2Ec0YWKlNSQZLWXXwTZ6qt0eST++VjpiSzgutQpp
9qdYM9YySYtINeH8MugfguOY65uhEc+fKcU+Sqv3cG7ekp7oK7Z19+bb2XVCRardPDfvO2+4rNgS
bsKsEL2rEhDp7StKEDsco9KF6bLvV8Ri9Wqz5jGKFDozCvOhUiWEz/nbt0eMDmkS+zpvZXz+Oj1T
xMDfCJPYtM/oC+jKbwxVw+AjCOaCgRvyYjsnOhwFLXH8dkdwvBlPHXR9uit97erVRoCcYORaP7rz
Fkv+ZAVDhzZXF5PX54YkUax+P9KkIo8SLuk19lgjvEX8xeHlaffDHvhD1kGatceSLwgDu9M2AwLM
qYSKyo//blFVsNbA88vCP3b1f8W5Yftu4vclZz1ESXPAcH5Vm7TdaVYFRlZBxxc/xj1Teyc2RRs2
L5EYFyXDCnK+L8RpKVIkq1rk79Vn8W6oT1fakgKurAjnggG5RXy1MxEyy8p/1zQq33uzSdJs41AG
6UspBkXRznv4SF0/CdRM3fMG+xRP+UAWgzS5e0m+brTpo7IyLlB/wqYABRWeJg2e7u2+tc2FUrv9
3QWU2Qm5pl/j7KJf+l1RCLlobEFONFdz801ZErYRDEBJwJ7Qf/2AgfefQwuz4uS2eL66hsBc30zU
5Y83C9spjcWQRQd8XnIqr+RnFgLHYlddr+xweDkpEm9+ycJGNVUzdzzDQLRS8v6kpGjNvO/qWbRw
yIPp6WEM8tmE2/fhYf5Q3bw3aZGzV5LWQCLNNM/F7uqkjgJOoSRO2DDqa49VPgHAe2DXjckcfozu
l6kBXWvs1idXD0rLw3dso6Gn0wCbo+SLOD9mdrEu7EkMsVDVRB7nLML4kUA5FJMbJCstoH8bpQP+
7vqaUKCQACFAVYsurf877jEy/TucBp34dXgCv6kYc3V8pPetyKEQQdKEXeZIrpdZCc3sYYnHVlVt
CjZ1mErdjNLoVHfy52mdCbjTPJBvjfybFLAb9RVXxiXGKJHO3uONSwFJlhg1LiJZk5mxr7rHPzHm
WfI/Yq7rHzdt0DlebhlGQTzC/Ob3YpFZTUX+4TY37SSNnO5MInS7/SL/dUmxytCkb6qOGiXg36+h
VCjYc1lToqbm9Y7qZoVONVtBV3Y1Vs0Bs3gzmgh4jQmALcacPUHNW6e/udfSYDCMbE6oifEwD3Oy
tK99i73heK+yIfkoY6jDmAL2L69lciglMg0rHwcbx/1vGYHwAxX/g7W9mekIo6aLlf1YchrWDGOo
8deIglch7MXFalsb14Ld7Oajdlx9mSpz8ss7MVJAjjzm3VN6OsH5I4em1Qpf7esMt79oR9u+AMLB
tjB55mXxG9y9JlwiAvgDlCbw6ALTwE3Nwfu2ubkLfek6AnkmB0Z6paqjDzU9u9i5z/u53VC866b8
kgYKNnHi91zcjBoTGb51694XlCjG/HCOCUyKZDkMBl1dtRnoK4OY3Diyv2EB7CvIIQItAcBDwhWc
NJsNUPkdjsvZugJMXQAU6MJIY6bLauVpEaUwpNRRIx+jCr11Cb3RnjVRIbsiE3kx1haXu4DJUKLy
C3VzjIeYXd3oJWmvYl/61CGMlyU7P7xFcqlXGjgo2JpLK+NW93fCcO3u6pAIPa+FBHJuTertYc8/
iJPedx6/jat+NqziWLvDYE36fUCPfTFvhA5XopDHn3AMGKEd/MRFIqZwuJ37HHvQjauRnli4vHXm
HjhBAKzMNXYADTxyfBWdaC+sgS8O4gCxCn8vSTYyeKvE5NOUi685vQviswb9sb5ohmyKql1B7/FA
QuWjgt5xNd+WcpJTfiikihILiOiPZJJgeAxixkISqyQ8oQ+oIlp8B9UGMcjd/GIFx6iyo0JfvpSd
20BX8tWqCea6ZTONG2tGdukKk4cDzfnq0gq63IEKDKNOW+NP08IVspopCt4CM2rQYzKcvF8VHChE
seyViS7y1JZeRPo/uGTAa8+vcBvtA6aP+DpE6QA4xQdk0qYwLEgHNxtvKe6mzuMK79b5Gx5wz/3d
RYw/KGOqR3ytqWvr2LS8S4nfuGQTyfUc/VJJHbrWZBdhEuCwnoYuuzq5W3CgWRWOOERPgkWgUBwf
955W1EeP5ApIAOOQpoPx0Lumfox/ngKGCyMPSjaN9SvHUqLthQ7Xqixp87/+wWzgrYUK1SPz0zmZ
JX/92bmtzaAMJ9JuU3OBHAZUq9aVHMYzLa/KlWln4OOtTFionMb6ebDzHQ7X+/UhySsEAmUMuHwt
a57O2M5fwLQmC5kz7yFwGWBPtJ10+0R+gnjTvxKNrr24Jzd8nzbgm+BXAD6G7WELP6I48QUartSs
604JUH3tTN90OLi9/HGZHUF7fHNPUVMnyarvGZpHfnwAvrOOH0h+UKMK1WXFpJEFJNJ7So7XalwX
7QctPbSlXTstHqwPSpxzzCbBnFa6w7t4WiZNvWlVe8hlnSTNjXTTeYXNUO+etl5ASWtR3WNQrqxp
fBeY4Jr+YBW+Xdqc378H9LwN5cA9MCbGKZ0NWm7OMKPNvJQ199h3RrOlP8Be5AjHZo/S2T/xc/bP
gqqRM1JDxI85gsp5Jweq8+IdU4k2xSiT9gKaRxTcFq3X1QAjPqUV26vbW5YvFQ7L5i5UxF/ZTLcm
WvFdaEKMv5uiEUPpXASjPGcjNkkMjOC+KI9OVZaHPoQ7uvTKzrEG6eYqOM8K8ifvlgcLdqIPv9OA
eweEcW+cbznvLhdYwv1lOVRzUMOYgOLFvJxFqLvRwHGjzHjlTuaTDFsiyV68VaHL5huzrDcBoHWZ
p+dkUReAEGkHMVj/+v/gHrk+OfK4qWH4eESN9cicMasfip/JKjd/hsA997RuwlU8L4j4Bo8Rrh2x
5d9QrRIFKukmWtEu3MaQYc0W2dLcMmK31WUIWskslVcivWxtm9eUJAmMtcSLLfZZNxd4Rk088ipp
oqAA9briaBuws08btcLhy+1o6/kEnr2y2m4wP++//uX8Tn4lzvbbxopSBpXXZbEBEftjkCgKSah0
qRA/UByr4vXTyOG96sHDcBAR6rEXAe4hviEcbH7jBJVNP2ZHSe40n1SHQFzkXR2qqVw4dMFYExqy
3+W5wSuj9jTKzIwi5rTFPcYtV9iACgr/RqwHDNhfnDcKjGL8hLtiYYp9h7ZKymQJ5Dm4+tKZusqv
STgDpzPvlka360RMGP0NBz+4xJJlwshjjcZQt/oJDjSJgBAE4hSFaG3HEijKYfMPI9Q+S4vvOtFT
xFGhtioIHgfjxwA3UvNvAP3fkD2LwMnx7IA4UIet1xdwOHZniACE/2AzxmryMTtg6RN5nNldEUbI
OSfAqbFAVKiRSRW1O9t5yxyL/hZeLaC9/udGHYsYHbAEbdkn9i3CAvtYwiXETOy1oKR96piJlDHH
LmwQb3GKHSMsXAwPQlgwOe710nNQtKUKjebkkcN4G8Gs4QZkw6KytO48fHKgQPX7yY9bewvsHxlL
blQFD3J18VMEthwo4/C1kEKZdmwMaK3VhDJrk9/6MPh9IQ80s3r1AqFg9eGdmkb9wqdL/9OAsRtR
ZEDxhcWp2rs2+tl6dkqTUk9d1+vkJMwk4bwlmeHXjoNNt1PERklC9VtuB8tMxK0bx4kDR2tLuN+T
zfPoqOaVA+1UWVW+BHCjpxogk+VViHSrXeQkuihnMeydmJD40SP+m5rZiFSbC+KPgKhcME2s8X7u
Cy9ryWTNfd5jUAHxtZf3C3cFgxSxrGc90y5UnCrjNv0rLMVtoFrCr7Njo0RNNTIbQVqKDo4Lmrx/
F1keDHT/2zWsFTUdgl1Ch2bGS/k7M9VSrFvUP3S8gDp9+F86AFUqxP3OAKxZXYoy5seiyGKtSJws
jSW3nhX5wVQZZXR7/FX9YQPAEjsh2uHGTL2LfGQngl5qvmTa2ntaYq+rRFsHwjieJyYvPawTMjB0
ctzdWZNQ0B5wjXtMnLK1b+zD9twoXl1rBB1+5eVFS0PImQr6IXcRvHo2jYA9YwclVqo5pQxue2Gt
l3qrqdZoRJbIt7VbpToz2fXsQleYRDjtx1fwHjQxLeZ17Ac1E9r00lpdAybyKwma7APIFmvJrtMU
syZfXBcoNkXLAq3dsJLa+iO9i8kngYs364Lo7F9Rnt4WyMyTNZzYiqchzOo6w+XABV7YVV+elUuZ
W/EtJS2HaXAAkEZvd1SlvQMJmWO6pCUgX6kUBaLxmahs38kzhAEIwQmQpJGusvrsqGT7q86ZFoNL
9afWoYMegBrQbWHdXNch3TIMakDtHqwaFkAA6k5XVWo9R111JeIYvc6yCVEVHRjVTiip8JIbzrCF
TXdR3JuZapxp74Ce5HEgq4mCJJkuxWhdrYf8kM4Y12khPCP//eMnsp/8TwO2tFzfCKw/oLFXRXhW
6/xO7rWbQ+tYqsSYfCOQjz4VpfL94M+CJx3sfQJwhGsW2YZDhjTClf7W67TGebRxnO/db0aZi8fr
vVJS3qfQqugtQmIYAxN7IGKOPyEucpIHNeUytJYde5vMGsofhqNBJaviNwmJfxvy5gssaqBei1ok
tNIQUa3UK1gaqecAaZauTAikeM1jfOx1BZ/07MDieYoMo7z9cOaccFlyvcnIv5shZtHiUQB3pjm1
creOrIsoaaR2Q7uly3pyHTAtzwonyJaAV/rcC49ToDJG4JwK5KfBHb+EFlWQZrp4m73ClPkUxQwq
FeLehHCHyYjuFGmuQCWJk96bCWcy5XAPQofOSu5VqsftJVRcN7w9sWxE4c9r17KsEzS1W5wkykNi
tBh3KEUmwZJtU/kE0ubUPZkkSyJRBesrhpl5aWHVbKYi7bogBEFySjjaRNJvcBiNfaame16iMBC4
VChnwl0v/CHXl3dXjCw5IiBw752nWcNn0WmWgaMpkGXWl1D6fe9mpL3eE9pUaFH02RbQVyQcNkGn
zc60zWSW6g2sOputgurPFeX5j5ZbpLe3scHCSfh8FiTh+etheVdh1ovDvHAoA9GU+YuS9agKJwe1
JNDAOn0I6XcWvRwwIhrCqSvbzXpgDXoGHtkn7qFd1ToVh7+qf1xSy6eouFp2SF+A6vaHYNIFbJgE
iSYby+EV3zvNXXpQCXIR/Fg2Yf+msspyyyJzHipC789BO0tLzK4L5T60Tz8SLjrzZa+Xsh4TP6K9
YpuJdCkX+LHjma2Go+RK/M7e3ZAo789WqyQ3NkXVyx1O0Tw6u4nKK5/MRMjUZULWb+zm4DVd6psx
7c5e/S2Oqr2/s+wWjHnG96TbBxbDoplZqAqCtGrIebR/9AlWxKvVMJuXOhOPoARaYf/kFfvatNQr
zCtHy9PQHT2dWHNBBWDoRWpd6g/iIHQkzF+JQ9FToidXiLBLDsqs2sPSL2CVPvIYpnrWapk5qihm
d6shQa2bgbwsnxtlR//gpX+j9h4s9ll8KIzhizYgLgpjX4swNHVpUVlQgXLg5rSAxDi4U0ha3cOz
kx10RGj6i23zoRsPfn8pYcM9cUmdjR8POLpSh5aq6+lus5GfaZfmqJp82/xFREq/J2Bdkr8bt82g
ZQE3BtHtDDu1PuKw3sXBh6ZsiRDokn5K9VAU78h72FACb5Sp7kKRKpxAA6gdDeM/eh7RUppWd9uL
Ne6D/+v4slpj4hwbrVpXTEO2n54agCU2ZgfRQV9+iwnvMWWRpQDgNE9c/C2ylnr0ImMfheskh0fV
3rshYI8Z2D1Cu+nL7sLbAPtI7PzsE/6MHGRq/JmJQY3swMCyNmOWF7hkEmp8ocruSSRKv246gkyF
4J1gFXYVsnqPS5BQxnwTUQEnzBwrA6UbrA+J37ujfE/tTBVDn3umly+rfZ+590fM0/wcbxyQBMTg
lVfXxH64F6lRzQxYi9hQzsqcz9Z/2gxiXgQU4znTocpT/rH0BoX6Vgf+P3sx5E8UmdKLemBfGQjA
sDVtG0f+dzwNkZQN7Pl392G5Jt3wrvExSw0/B4YEeibr8g4IxEKGZLpDFZe8pLAxUjAcQ9Cd0FJ8
KwZLd4nthlkuT+OX4+hFqzVcHpEQibUfdsmo5I4z6AhtoGefw1/RFBf1kQTN4kDXQA4uL3c9xeG/
VTkXpFoaXpQixFVSqW4he4gSX/UXiZt4ZKHN45jxPBQGMTnCWq8I6+9nC98dQUpqNQfb8tPyIGQw
iZbwi03kN6Eyob4/v9Pk8NSxKR7DfdaBskW950hChUEiIGZ4YGeqyMHwP9HaTIGOVFKh1iQv7+Pc
F1NM4Lv3uu6l0cNpbkbuACEoo3lPKwr6DMnmjb2Qn7WTUWKD1myfPiQH7R0TIbyLsxIFic1gR0ot
n0LK+wmTAJmrQNJq71aKVRbyhkx29x7D780zOwpwoti6nRXF2WgIidWf0Y2gqg7b1mR8JSpsOyFR
fuaL56V+uLBn0YyvC2NcxMOPsj59sHjjppNsgPgreleU8xKBaU3xpFhjPotvGrJuQwXcFvIJxgER
W8gz1R5uxrLBDL8OsMjw/OfYQje+/Qd0bpFb/kLhpRNGNT3yZpeHqbSwRCquCjgWF61K1d4hxcgS
aUeDQzEQgn+EDfdVFmrSL7IH1w9vdiwM7Tkr1oep/keJrJuG+luWgpO36Kj/GlRxRmcnOKi3yz3N
Ujf7hjKp90v175BhoYOo7GTyBL3AnATxoBxovbyq00EluGadSeIW/rNQf1inJWhD/RbPd39E42Ky
/uDK9kQeHcGYd+Niv69WM4Cmt1/3uXQBBbBDxc65Q8XSmsBxSzlq7MGMVa35BXoZTgF+EdTKvMC3
THKljvcN7pPS6UqZ9Y6vIR+NDXmOhnrRey4XwmgyR7kPRCMbIyHrI+8a/DBvm1I+britR0spg98y
47XcpyWsVcy0AShGkmdb4YLJqAvxZC3/BvukuEHpz0sxACPeWSUJnkd7pLV1PMi3ps31j9v4V2JR
x6ABGuTqSCjEkFqVr7yqr6ViORyJ7QhVsse4Ju9JLRtHXcrH7JJrNT7b/AIdISRoXC7A2bHNU0Zd
Vuko6QYRP+jOrKz3dhoJKwZjVu5pf0WCQ9cNi1sPpENLsz1AuEhJtrHfy/ceFqikVyHalz/+dgQv
tvpiI/Feth/E0dUR2jy9QuGOf4Wo62Jskwr0JkU2MYf+4l4acYybbRDYb4unY2csr1qX7TjhurCI
rCu8Kfx1kUT7YZvoeVjA1ENoTXFf4odzC9faHm7tlmSeydw5s5DEnfFlK5PT439nyaoOd90SnSZj
VlewLApPbIVMmHO2XKI7WVYoBPR04rE6kZT5zUFWDDqY4yr4GQ0BKsfc8u2T6QJS+M94/OKgLkeV
Im0XR5qQzLJ29Iaj2WpXIM5WcEQZz47mUVUam9pXUP7mjMzL5HKaMdmkOliH+Sf1eYtceqq9PRLo
e/Sf7ToUF5AV/BOmM37XtTiisv46tBAgD0jmh7AIAaJbczE3XgXAw8KJ9EiYsKgLNQEdfkYdbK1b
g9HyKhZcxPnFhm068mYZPD7A4Hwtl5ilT+wQJ/2ID36KlAZXVRoRCc4g8CvtBVNpwS7SqaEWUJR9
wGA66lc6wj1FXipx++UZljyPpes7WRXX094lE65TAv89X3w2n+D25NyOqJwrxKtnVYAHX8mryVUR
0mzvGzvNerfPAlJUfw7PWEVZVxnB7mg/uYWYwkzTITPIu/tYdNUD1RKCUwAMyheGAjN59myz2xtF
fnuWtX4Dru+qbAugxNJgtKgcVoJDQAWfFhF6pxaajfhfrS3QD5/amLFXvn2sE5QgSgvlgMfVVExo
NrG7O4BOVrVtRZGLOvx2XcoYtqeVGtsUy4O6eduxi2653ea7z49vtcDB8vyO1wdXoDJmmLVBqk+q
8kqLSZpoyRInHgQaqzH23KcmMauNe/Y38gCoIoQq62GYcplcL91MyKHbOq3uILiHoR7gWfY2ueBy
ZW6llhRQOnaSjszlmqzQmf3OIYi5dEDeVILQq/xi+m4LyuLsHiKIHxR4/A8onqqVsnSweERrE/NN
wLcL2Yp+s5+J5KJ7WPAm4j7MYA+/Zuc8N9eAKNy0A9f+3AWO20daR75AV4bn3pYPru0eeW5sKv8J
m0UBDmNTEMyf2MAzpm3WYblUvV8avb7BvDuofZtwksuK7JMiVD3beQNtmC/ADAd5/WswIU3cOu/X
tQNQkt61usUCjTDIgoyHwA5zeShvqG328yygo0USsD8GTIdtivNnmYITaSm6+NI0sj7EcaCPlE39
g91sZiJMSN4B7vlG4ED1/C0A8etELNKTRIhQHaQHVArZ3aj0+nt2keFINB1Rk/gpnqpFj2Awrqft
xEgLFMPQ0NntPkE39nQoFafO4tHlTK/kQWLeVJMCrJ1rLf05wDJdXvvAmqzTY1lSDm+rt/hF48Fx
AlQVZ7Ao55Jwu6JT+eXlpedAoiwDlmoRUCOk/Gx/IMkLPapnp7ttkIzuc2I47ZJgXf+XV1d8A92D
CPqp/MVusIIav29zL9sP3b44Q0WW5Fl04niJ8NwoA5hVxVZrB3ATSou7I8/noctD+dHEXXzw9iL8
Fe1t99wQ4sFBJjwOs2u7CUjHKwds21OdHQ18wsFKU2hOJMVml8ZRQumefbZXfVcCi+QFgtpr7Fwe
1ug1mRw8OQk+Zhsou0VYQQ4+7YpFJuCAAtaLAujwTsxreJ8h0r24I9QERbpeycL4etq7TtG0x7z8
1/+JtJIDsnhu8t73Mfs/gZ6ACmMEGO6VtfG7LWN2xQK3+XPosvdY10QRVjHex0bGoUy5U9iLUm5G
9EzhizfD4sNZ9mbWSh4xz9Phf63HCmpvTm9o+Ugkqws2FEsNqTlWuxN/yNFcVgP79D+dnfjF9P2d
6ACDAn3WawMOMU0n3sAQEy1PKHQQx1RjZ5tjFbKwbe6wIW0NmoUgPv2zunhpkdLocqiAMRqQovpW
mhosRLwSmFytsZdynyju/SOhb96nbIjYPfCGwMl81ksq1OcLBwq1m+KmSqEZDC9K4fZwvJHiuuwW
/tL5WoYpwBE1osO04l1eaQd/v/OuzOnUgf0NX8KJFjlzHqt8s6aU9YQ5hG/NYqOhPMpYUACpY7An
OY5pfBgi9AQWyDa76WERrh3FGRgI5+jP6YJcaBe4vcLOxejAj+91n+Hy0n2VED8n57LC7Qhx6DYS
hA6/iqojrvwMeA6XJMxnxVKDR7wTrDQmkaYvWj9Q+DCaAWnbxd5gLo4C4DlVJ/RyckSZzpKPusqO
Vq3biWUgZUWH/9yrNPa3WWy6T1Me7r0sF2lMsQtUdMZCBl88fd22kqeO6LmQLhyO4D5B/laJhsfS
inaSm7NDEoCh7R4nu9om9H/HcAPu6cUkvnQp72ewdLhvWLC4gfBKVozc8PoAqZEHWAz//dHH0gtx
juwuTphxhnjFt4w+YdAlJtQsxQYQcnurNKe+eJsTlHcxLlbP0xPpYH6dRGRtZnKgJPe7AxsbB8Cj
Ml/c/2STZ/a8t41mLFu1GZ3K9RxPAokf0d8K8owydx5T5uqdanAu2oD08JUxZh7IRZjmG6nvH2Q2
6w35bySSP0Hx4WQzA8r5qZdOkHa4Nrowqi4dwME+LNtWNJqHUgLx9bjmnk85jtonxSNSs+7wfGNj
Vk5/JKKLuT3Oss9JyTg0tk3epoRm8U5PtZGoM16VwnEEk1C5EpnQMpUakWfPHKm7rHG5d2tEXxJf
f66HGyjNRIjEtHR4j/y5Fme6nxrbZPY7gZ1hakrNA/7qmEGJj6w1J7yhcQcTsuq20HDifHwLmxbn
xx2mNumeHg+xghmV3GQCSx/vt9msEFhB2mraiHkPROSWZPu8DJwr5unJ41pYhmtLDsvCXS6h+LVZ
PSm3PsNSEnFZSQQRYAQbD6cYPFWdBXro/uKtB+qS/oSAE6mv3i/DqNahIoRCjxq8fZas+WwkJj78
9rTbX30B22/NswYdpQ8vOUtbHmwtix9752JYM6Fo8LhXTiwbrgySe/4M2+3uTuwbbBF8QBj477gi
66zTLXfEmH2ASSFcnIDDPTcfr+zI9fCL7pWUvV2QojGrpUtYh8JzHtIuG+kKQUt5rzXbSLWzh5M5
526xQdUlrGFYpSbpTVMbgSeUYpUZ/NI3z+3+J5yvKX6yNypzs7owlMP7yL/xDhK2cNGucKuuXqw8
Ih1mf+hoSI2L6VpGQhhGbeMSGSVuINihJjCsMpnuz9HI3dwmr7Jm2tsm0jVCG7J5Dm+lo5lkvrkf
zdoCTDiamQFOt5xWbTIawl3KiToYnZ6OSf5eWX6+EWaNhhqmCMPILuUioJkHrisFs9iAz0cmL6Zl
elDfj9CIy4JIYsUvLS7B3tfIpdj62NcPeGpALbkHPt+wm9WnD4cLh4xy2XKhXsUuCTVlruardo/P
tWmf/BME+oOIH/s9PlvrfYkYYU7R5fWiupm8h+HoJ6vYYx2tHl345GsJzUye/uzxbL5blpzKiIKF
vZxzA4e7OfGdV4fscUd7EUasmzRSdwgBgCSoiJXnV/TEVtr6yg1FFiVYKAZglf5ro38Ce7eh0GZi
mxu/T/D9BBXJygvtNmmDu9n0s/NR+rFyfoPZkWBhiqoXDc8sYsJIu8VrWxkYaInjx8/GqD2qJwQ5
TCNmf8Rcb0RZARQs/VBZXEMy2jJmF1JtMCwapqzbVn/uKl9OgGoKTiQQhol7K4WamflGXcZ2/K/7
0dsF7flM7SUQOvH7ZspecuAZ0do1yYhpC7DClopQile2Zi3iSw+E+5RwkxabYu9eDQfpSzNzwD8l
cOvbJO8RAZ6XiQ3l2PoGCrKgfunNiJ+urpzv/ZbAsvmONulBLaU0gxAtajRFcBbF/wkSxC2ENnrp
7CxNMdgBXaBhDORpxQaEbdlaDvj3+gUfhkzrl70E9UqgaJ2Y3yBAezOb8f9IcSWljfGlMOM7Q+Mq
qgZ0fPfPHjVtSivIeNbmi1SlRoabfxBl2GzBtKWD19lcgmycDT3kFbE5z/dPSGuAaJYIy9FW0Oi8
sazvLefdcKxhlkOVqt5yZI6+3sh8G6aceI4AKfIM9b33B5u1z7+oCuIQk5dLhU7e5l1AMUqRtVQF
BbjneX8jXxtn67mJMBuTCK4GHVha/TuVMNceIOalxVBnkGl2rREgJxYVmjOfixMZbn1AwlUWqMku
dXi+tYlVxXsJDRDeMLNpvH7Kw9svGzl97QvdrvPF/8eVaNFctHrYIqudNgRcCjs0CRW8jgqe9GMT
ol90+SVxudEdo4Q7SD972SrlO9azPfV2eQRMB2Q/fwIqPNKq+mwJze44X2PuYfJvl33pNybrbAyA
2wap1Z6upwpe4HV0KIfcYTPQ1ZGOn/Q22MLlsKSomwBgm+bugJHtKWU1in6C2AnMJlwzErJ/ZeQn
lk981bG7qQD/nnrJfkAmM+JKScT0DksXdYPVCZj86sFsQcZFtVMfZ+Ego04Z1eA19f/VCsy/lWij
GjwJrju81ABlgup6//ps9y/IZ213phxZ9DsiotegADmCIrRXQdlB95t4ZnvdPwfOns/tctP+ozeI
t5pYtHcJjzSTmNQzDGGQJmMoMKBTz1zon25KxApL4ipD2PgRMH2eZkEbc0tS4FaEp5kSmI2S2bDW
hq21Tc3ujt4SFOGutoHz5+D3vEclIUZmXKoktAXSY06ah2hIbhizFN5xtQBsDGEXhZC24u1B4k/H
FdvpQue/hhzbU6umGvq++uRWXyJv9rV82JRv0WSjt6ARfPVwlwpjHUC/NeElnAF8Nuw2w2q8jD6i
2ON2U5flcV/ZfWEUtXF0isgtTL8ce6NyibZQYOqQRB4N7Z10l0e9lNuyRhcb0YSDUXn7P+xaL4eD
MqwiGlRtv/ovsqVXsx79PRr+QlHBW6J7FZ72aSTtZ3t/DtmhHkP/irI0QEhOkblx26dgsCHGHbt1
68H8GP28pf/3WChSfzjRLTYT9jr7QhBIfIcHDEkH7Y77w3McdWowAuNerbL8QtEY5bL8G4WYz2Pg
id3hVprwat4+UsxtH7yjkSsZG2CeKVkUPJX3w2ORH2TkmZZiMECat2+mQ3iyYKM9avzxmijAhrzu
P41wBIvPWrKqg59apSxRoBGiT60B3z442gjZyYFa2lRdquicHIETVrkVattWKANLpzvcqHuilskv
cVh13iyZ4pOKyP6MHcwd80xEBMG2ebftNUPupbGCHSnioz9NF4fb8XlRcjoQjsLxhsbB36+23ARS
d4O0+J6HBGNwyR55Ic8nNoSMT4b3bh8ttoy9E4dQF4Z034iT2rTQt22LJGBRd4VkTtHvdP9/Y56Y
hz0y59pZVdEFsVMl5l5rObooqPdzFeQJkZ9Ea+KEbYu+OoarelNXr3WvIUn60RPhnt7g6HaDxpmN
2E71Kmh/85DnPzVA/+FiMbFbX5ZLR42TPsklJZDu/sfJvQEscMLKsgsx8Jpz9r/QI6NLpvPuUSwR
kwWkFnMR2HPxDUKLD1hUPUjump3bE3SMbuTGGtEJszx612fpsu5RbFgKnwuYcQyYbVCOD3lbu6GF
v2VULhBVrWtlrxLAtL8SodLo0Q0rJc6OQdQez8mgaqbKz3LiePGF1mTkI4dxMOulKoIeR0A93Exc
iwBtAXM23VGdHms2Xe3Q5QCpB/etLlT8dJmr8tNFPKv7Nhf5ph8staPirBFhfIxVhxIxpGaii0xk
QQa8ms8Gk2Ll25iBJL7l15Xq2V/Vxz1MTAM5Cj1501VQ80UHdi5DlDgh53h5tjZ8x7c8J2euyMbO
tTUO5wevZLz9nidnf19bupUWA0/HpjRAs8IQo32wsORJtgS9682limkNUhsNTLUavkF8Ny0DU9Xa
U3N3+t8tZfn/mBD0uMTQZ1v7BoW88JzTlyI4hkLw8ui00SBUMTM3oQZHzYI/dCb+oK3rrNVo5B5I
UGSW6GlEWkCyUcllfmKjtwKb9AobOGgHzye3G9U8jawxUIKbMfPnlPWhqde3WL4z9/rmbGIL9g/e
dDlNWibA5cgB/6WSv88jfRzKIjwL9IgWBT7PLwXJU1oxvJxTTlSwh0Y0lMDkVOi5DIceoYEUkCaf
yUu2MbXvG9eb2wi6DMg6Q+UseGySGYcMSgKJ5VGxIrAkzFTtCjljcrx4UJ4IPGZLB+87ODLhprdS
ijrLHR9+yKHQYQTx7ylL9Vr0VmaIOCGDw2MpnN2Lh49KYat9Sdb3YDufv2r5IJQN9OAn/c8JfN7T
64mZYFpr/7E9GZPr7Vp5aTYJyngnjGQz31bLox5CzNZfCTk67D8/Yn1W6Qz1xbr4ThCNoZvsR3SK
pUTwwu733zv8zEQOXL1u2tYWB+/gboftYAcPjCscmFCi7p4RKNLLZlFs7oGPRA7b5zOOb/VQeewL
TY4ZRYIesWJk9rzAzZByqDqFycDy6DJwtmDpbzoST0yWpsbyhy293w54fKXjpnWPsDS0GPJuYbOK
GFMThirLAs+yd5PKGQQehxKvZv7etFy40ZSUhRcTxf6Jb+cKZB6OmHeGe7RfysE1zdlRsFcJyks1
q5VCptFl1hCBzL02D2m/OPHAHeWAG/2Ek48pO2+p2ZbglS2qJRVVYOq1a2ONQzapyXM6sFfvFitN
DGYaiAwLGIcm3HIcJ8SpqVzaP7pLb4hu+jcvvYPFE6TfCixfZoykVmfE0kYXAXMcwbYRfUaGsUC9
JDpY9dxZm1PCWSsgbLPervjcAjm/6YXm9OaC/AjgTIvpT77qQdvmRsP9kE7yKzwZkMwi0eCDJX4B
HDk37RhqTltmHHbSnUnWJ9O2n6KSOm1Bb0HziJNjCAqdkuMpgrhKBKfNk007VNbZRcxIa7vUK6i3
28RAP45x+e4gYiL5NDI1JKEe7f8a1C8A8OTeITLvMOkiii1qOs/7ABORZlhWE1jCaYtDm10hiHAK
NLkuGe2UNINyQw8bbOCWLjdGYqKbTgWca8AxLZfjHTPXCVrWy+8v5tggMmKtUyCneqTmXFFTzqkx
Q1NN4a5dkkW2fC+wKTkxNZGO9V6MSfoZC14GxumTu/ianQeuOfthSaibZDjgBEuAyUktyUXGDOXD
WXMSnuAz4RWxBMWdcth2Eq4jXjQzCLjGXWJEvwTMAy7fJ6LIynXvoEEP0BDQSl9WGA2Nem3+Ft9Z
J715wEeTUAgS5z8KwQbvCGastum+K4znKRr/Q4LUGvOT933e7N7VPUw90YlnmU2fS1T3ZbeDwBx6
hcGY9x4hAwINaG9vc9go4gN6mtf5Ke/JUMnFSS1+JhhZ9S86nxl41jE/69BqfI3GF78IitAfr+ad
ZqIErSqZ8Mw11d10s0IGCnlSXTkUuizcBfvc/yyzrUBwCwOzolbP9QXoUZtGWzjPSd40asL5ocnq
/eoaVnxTf6uV5zfeavASGfUnFB/+vgXd4uce7httME/yfJuBWVZ81c9CxCBuJGkHIWNc9WeILFDY
Fi30DXzKYZGHJQeP76g3DSLOq7gxLt6drTfG3lB/ZeUtMmqndPVf09PuIL7y/4qV027ShRJ2fY47
cCHi2r2EeQTv1+IetERoP59yGmcIeOvZWggWlj8kf9u8PDX0Bt8u20hCDltXPXuegGf7EMWexH4z
Y5F4FKcUD0+6fn8yzSINBY72920Doo4+W1dJIDgg0Mlnkqff/TGVaxyiwxOGgoc44xItuJxjRfef
iQBDCT4fbvoMMLJts8XRXW5QMleRxUfUwATTLwYHf0smvdAZpWbKPIPK7b1BJJfMZfsSZtG2ec9L
DrrxtnGyw8oBXv45bCvk7+KsNNdLZ6PlglM/SvyaDMqwRolPYhNirPAdWDHk0QF8eWJOFbiDjqkr
+ItBJCWji/082W1rr2ot/9/rsiwtvW6QK4mR9L3mCtAKReBcU84CdMv4euSZ8kcPSlglZWcg5LZZ
SQdCR3Af9TaHTquOJ0m3iv45Jx1EboX0PQ7U+O45WTRpIUwVN6uZymBPJ6LysDiP0Dqepx3d0Z5Y
cVOfzAYBhteXD6VuO2kx+tQtu1c0YZjoVk+ULVtWwgTp9nmn0o1MpXercni4gu7Q9j7UHp2IgoVJ
hJHw5JsQlauSgP1LARV+irCNklJWeu8Y6CeA6tqaqo41UNercjIlTx/cLPtA1hZHXZoMtOj7vR/c
O25SLHnKtVdaFKifmqIe9yDvlvItaqV4DeMvBKFPzW/WEuOsgH7Ltd7fudbz4vvel2Q1amHe6P2g
EX3X7q/rxeFKUAvqe9xGwwul4B+mYaKsIzdIyS43yX7f5mrRCy5eumnvHpbzLXucnniGOqX0dyWc
oFDEH/Tlg88YHkdm8Ineg3q3ShibKu2cu33/5LFVfd2FJbieiCevliwz0UgI1vKRWQPiXBMPCCCN
ZHo92bDVnjwRHO2F04vB5sb+BzYQ7RsoOtwtJxSWUI9phjf8X0/mnAWD0u0b/nQV1kgGuqBGnvj/
pLV7MhULr7/KeK8AyJLfWOUKBZR3CEkirMjDnrBsXSVElpkHWLwC/44UvIUixJq82fC4eqrkJboN
nrBYNhzY7fCdqW2CVIcELduxfKlRhLAL+j423gLtUxLZVoixatXVTypa3iRqOLF3gnU7+CHzrDU1
FEwUH6yQdA6Wiy4S4IBh/LL9bCAr1L+ab/ZJpYKgQprNcK7KjGYKcdmh5H9QbFH0/YrqIbUSNyJZ
VS/EPIleYJzH7qWFCJ7AZSXCC7GErmuv9Oqw92Ltahd95dwO9+Af568JOB+pYo79ifJ765ngzPev
p/eS4l8WTMuLPPSpSYaerYaA/gAmetfs36cYtBHi3O8xnkspthG7sNk9m8k+ffxoaNxxjpkHCuZf
+391xwyMtBjkpqIoiooANY31kR89M5Di6IPoxlx1lla8LM2F6e2R/nCHXFFdeMmNHkSDcpIubodt
epYH37hwRf1WDpjF2dbgUsCNDHA9PH1F3XX+jk9L4Cim9Uo7ZuyXRKI1qnUXVn9ZE5Gt3mwS2jGg
WCYiEqzUtJoSD/6RN8sJ8Z5mHTjp/hQVk8E6udQm+mxPfF8OXBy7nRluLrV8o/gB5lihnNwAKJaj
3XrTKkIJDubMCiEvavVmGFBgKkU/jQqX522TeAAws35Q4EaF0wiPoZdT6LDpFZs+H/MlHIVkQjwu
fI1qPgRYjzD3CxhSFWV3Riy4p6iMTlVIK2ivNBG7xJNV3dNGQHAzoBJi/6smXf5VbrlDJRLw4afy
ZU3b32/t90Ctg5Qt+SzBBm04bHKM5XGTItF9Qc1T6o7udhMdL8Dbn9TyQRrW/g+bZSYC6Qk42PjF
gXGqBwe5o7gfWc/m5GRw8SpDEUklNI/vm8cET8c0zMs2KgQJusmf7wySetEL2S0bRrg4kd0Cr2kh
VbdMt+Gq7TwOVaj+5e43WqFMFZ3Pe/2LoMvNYhJV7JqamETzO7/v6NFhJ5VmjCIDMBSnBe5nM/s1
+0jfJA5nakioM6Ta5spfhUWPdM2bitd56JLL8zn2jvxEHV/HOCDdYMFPrGhfsvwXEBlr/hkQ+x6m
7WBrmUiandl2KSntPsvgLV0AcFgqq09F5W1sgN0eM7r5d9ixNCx/1gv6cgBfo+9fP75M6/04/4mx
M2p7g4G3ebjXXmqhSbjxXoKwPKjyMrPRfDDb7hcUR+X2ilgpLMEQIhJlnv06I93rPiQoO20MDER2
tjmxLXWQS9wD7ELO/v4yKxWNmISk0IssAHecu+I1xBuif/oxd+uYVuhKEg3xgRbmyctqLCXEfiH8
5wDiDWWhvD96onXqTE7ut5uG37kszuVeZmuJr9IZfulxYtgw+Kfr2cy1w/oJyNStDytY6ScF6HJR
t4g1Cw1pyKkPwjnqaVi9amdQ1vQXALHbkv7Ycxoa2gOYXUvSNPcvlPSoJ8s8Ob+FZfZQUoTrza7E
W74JvG1Rcbt5MEagDzNy/J4npKUoYfVNKHqNQ6JPI/UkeF+34dlczp1hN72c6x11OAyzIUs55vLp
hB6Dln0r2jdqf9rjd61dogWvaZAj595cCO/M5ESCFX8zVIQw6Gd4yKr4ews27rezfIHSDx8/esCi
R928gwkic/SFK4Ndg+ZiFrAMonCZU1rWwbvbOKmv3ZbZRDtP1YhzufsQjbv0FdPu5Prqwgy1b826
35+o+q+E8yEDz2ESYs2EIQtr7XNg4eUUpeii4bkS2dzAh2Yd0MviRIbw/fH9Yc43lXY5SY5uhKKa
A7Siygh+0A0AzBg65KAlHbLm30o9q/NaK8QNyOynx2WARvLZKlVD/953cHh+arKkf9Jo1npI2uQl
eJDewSk+VSj9YKIvcNsSrDu7VeFvwjQHXcbyV9So8ics4spNlAGYmzaVCRnzE3qVGHvL9SdlKGg+
tnDQ03AGkzgcNQlyGgbXyDFXXDGLLs/ogimRQ7sX2V4DnSzE+kuixnywFyIlru31icKPsC1kX71v
mvJHZMa/VmslvA4OXxOD/vRy803RPySm33UnMKGI+nX+N7PPE7zUOPPd4ncSgXCdUVZN7UDEcTJh
9PY1uibPN+ry17ytoIgAjsN60I0qu76Ei+VZcQzF6a+RhTeCYT0BnpCybYlXmnF7109nE3BWU2s+
L7l90JTQDzrt2H3I3nKG56IJuitNz90hPNIGoyN6Sg9qnvZDr3NG75Qm/GPZRkSGeJUl+fZdJr5Q
V9baMHUpUu+sLlVtdMdWwHuqvnZi6fQd3HqFLiEYYWhjPwJSTJVZ/UtbOtVuii0p9VNS58GxEEgr
GEnA4Md3IrhKPtq7aKHMmzyXAG/DAmvni3hi5PO4qeaE1yyFjM0PvS9/A7o2agjuqzFivUovCbaZ
nScUXO3qafUFtvhmjtAi7mFc0h98z8/NoRBh9FH0EtN7DfD0oFMBXYCrkHSP7r5UV0vOTbBoEsp6
NY60HfOqgp0aCLa7ZIA1I95cbievxja91HQDiOgUsLfF5/lGOQl2GYaUJbcEv2xHsSiboXtKosK7
TVK380FK6au/oFKJf7/k2PhQ4eXPCOwhyyUr1zE1Rs6zY+7yo8DtLxw6ZBECj9iIKTUnuQP98He0
Cbl+bH5XRKsb6SZrbSYiNp/9k8qDbaf1rGHN5EEzN5sU/9M9igslvAPSJrc9oiyOFSI++jPNjw2D
JeVd7saK2/j6nNA2E4s2T26viGwy3WWa0M+n/CLUG/6iBeZcdHVvldJonm9WBP7psszEmVaiqu9N
q0JM/CthcVUAW54Tnx5Prvwbdx2ghr5wwGwu5Gxb/5UnMZUbJneKVhrxaL2Qa+XmPzeGvTAIeXNB
c7sOcFa0PFvrGZcFcrGQQQq5A18FqrBlbdxaZStpGLa2/SquJuWzPTbajx/H3DNLoGqRGF0/Eue2
YUFEvuHpL47CuwC0xEKYv0weZTCBYHJ9yTY6e910RNJqUtD1lETslpOFMLs+fVIssn9lmsLI7dcf
3Zcbyrqk2A3LA8z8VEsMvO7NKJcOjrBjm5ZhasklWVawcvBfD8wG9xXcQLqJG/YX5J0Vo7ImUUdD
k6yzIIvI7l/am/ay+I2MaNnG+2GzE4Z2+3OtImvcr3WO44mHBOzquv7pMDI9JCehT23TX5jsaqhn
MwHslRFtiDZV2Ext7kEjIqtXDLhpiBWp4ppiq0B9zlmzPidjD6hONKhu3XQI9K683v5gP/525qcx
InDIJcurVirNte+bJm5FV2DVsXV4IAdE7EeskQVaZi39w0yMwoDwSbukJbSgjQNeSupULe0L2I+c
/Ts+sFsEbTos+gfas0SSvjOMnEiTJHk9yKnD2WQ3IIB5RudC2UmDRgZeqKs3E/VyTWfjFb6GuYYS
pWSOzhaYfTs/vyxhZ3lSUMGmHggUaA8OnZLVlDQCmY8Bfu2gFabIa0p/oZW/mJDN8FdwMFts3UB/
sQiuT7sGTeqsGRfMZv7EbtHf0bhcans2BEkMKj/RRkfbcpPPQ3N+HYuSB6Q4HGehWodjgJEUv/Q9
Rf5z5eaWGgd7Ue5+ahq7goafaMMJ8yvS9+Xf7BPo3cGAWWDeltg58sw+MCib+cPeRp4BGHD9DJD9
wwG0bDjgfTWg/iifxLmxkthUtzjuWFarrev/iX/J/ybhqoNwRey96cc2Hq+YXarFMP9btXK7XRoQ
faqdURjOeA3f1fxZVVH0fM16IZb2FgJmEOG8l1qwY1iRK6vEApslw0zvESuXRfqnys6GDbfYLGsA
L2eLha1T65MPRmlE/yl7TBXCf+K3QyqYqitU9kNNvFoEYMjxl24bSVybsrnPh9HvBXKWZk3u88Np
EiEo4ahVUVxtEYzIEECWVYaQ6zWzvNG0NAdMNpJiZYAZWjVFN+V1bc4TQHIEZur25R9l7LBtbUR5
sRDzkNKfA1jE6pFfjtnvnywGpdIy0PfPt/IvBODDeJCtvTYJ0dchyaMdQPao9hO3S9kNyYYvZD/D
1EluOvrESla2hq2WGNS8Dqh9raZpYCunMV/I6pt/b5bom6WdJRuu2yB+RZ23Xevg+53UEfB2aE5F
Sort8RiYp4BLt0L/srQMCjCH/Ij3vo+aHbae5pbUP/VBOI6dCsO96QM+Na+7abvjb7TGTa6/QWFe
7XBTK8rYqWJIU0itOY+kAB54sf1gBGuFQcd/Yxt3dg68XehLIOB3Kweq7yIICJ7jRGp2+mqg2M/O
68Lnj78J0T62gPlMW1kp5yZ2hcnZ0hXJVVJo+93rwv7GpAYExT/Qeuq4RAWYhgEylrOKFMv9RVKC
duHUtBtsvFUN0Lfwry5lj5dM4kRAx2O5ZXBMjzqdInPRrlD+5y7AmL62FXiLblb+wn1QUR6KIfbD
KRdMuEBquQlyJskuWNo2OXf0U3aK7ZNQnsl6YLnptZkGf88V+WZI1kEcsZJYyqMmMrKRyGUY4Tji
/W9LYEIoDhNFnNV0EC/DvLYtdwHDc5U2Hadk1TKuZ2e4qcLnPEEHuTi+DvU7K8+/OWqaataGPelz
EVx0BGNZYMDmr7dB4zsKL0f4ZThIyiy7whjYTHNh3CNGweCGzqK5tlP2YlQbnQOXoP7jPxL3AVv/
jCuVnlyhkQZwPSMewbM4DbgxNS9A4+2W0MpLGrb3vmgb7fCzCo6vWvvQReYNF3AU/OKVn+98wOv/
OWzrVH2LY1c8aHnF2lxIVRVkwrz+A/RMlFDQO3wibdICO27K10PzYaKrpJu/yD1nzmEMo24LZtQd
m6nV1ilRZQLO2NhEfwsyqTgO96ZEDvUBjJYQUZE/U5jVUuVBLhI/ob3OPT/27zAgtSp7C0/BPqLx
Fw1Go4HD+7mlRi3/c+tQAnBEWxMTZ9lpmCmwKMoqucCK1cKwa+V6vM16Gdx6T1jWh4g/RlI/WzC9
pe4aXHMTJv6aoPzUy7TcUzmCOl3VEQN4L2pj1KnaGWUjveI3d550mvGd/25MAj7oznVZYxC9HK0k
t/O1hMK2uOtsA4nrMaCJgpmGBSa2qa5hJ0lQrxX3OsLBZLpT1Ykolfh7NVFA41Lub7JH6SAqeFcq
Blz0I5jZN2f2/KOcUSAj6yjMphTPV9vJyyZM3IWWBbjiJPPZE56GXgPy5jHpHvVYSoWQkKMhC6dP
J4b7sNizEEWIeyOLqRcOzhp658bvcDQw7r4htFUyIJ0PKazkDrYIVL/cuwTONZc2QfRMxGnngmLM
ZI/I+dICyQUmNM6uJImEOhCRUwGazZ7KwZh62jlSoDj7EunbrKKOQxP4BrPAdfoRGFhwRAUN7k+G
LSy0otlTkXEJzc1Dwk+o0ETIUUkL2fAtzSdKRMaJ8SVNp46d7JdNRXUvFUF2G71q0ZgfF6o4ZaYb
IMPGwHsYdRYJrfUlpCypID9gyJBa7Haq9SusBrdD2G9voECa6uD7RGyY/3uvMQZAqINh4oulHvI5
LL2ukby3BR/xQSRBByGn5aZgqkhwSdcuB9h616VVQDAIp5ilNV4vdaPBbgNTmW6PJLkmanqjQ5wt
Pxx2UQC9n50XTA3M3vTBvDulHDcnwVkMAqmIfnNi5tI7mYW8eZHTXks5L85vQXrk0SPnv5CcdLJZ
G7l15MNzp5pHTtzSPJYJ/dUSm8PXTNJjx7v3Z4FYqarkdxhFf3SIGYrKB2/rLnFrgs3LkNgKDz3x
bzLcij8Uo6LKhki1OfNtGmVsTgfuuIQaaRCLb1c80xOp5sctG8sV+/fzRnpMStf9x+Fe5er+5Xk7
6YwYpXyfgh7ZfLUtiuoCnA3lypTjFnA0ut5Y3PrNc8pEvx/KMX+lpqbGuM64bYze1gZ9Q70gM2gz
tKTkpSfVZEXv8IABsXoYdJBMpGW2fDYtPRR2QpcMhESVhZQEn8D1IztaJjwcBYQSNiDUnPwikp9h
sUUtmWHIPcwtkmxyuDiNaiQwgop3dh+88kUuDVE+soH4Vb9ZZFoRPlxKkRehrtqKu+fzv49lMIX/
vLjLq3uzeOivm8R1DGTwpEAspnoWuhQEym5qvbVOkCGb/tICQIVT6qlel7y0wPr8eqED/wC1pxaZ
6ArrjYtmiMkyz7EZApExCF23LRC8FIt5XwT55OPXjB17HG8FuMFxhhHdBkW77tKhJKyx399vJnAd
TipxVTkzWb1bhicgQ5ZdRB7LpTChoC+iG1zIhWFzUZo0SKbdULnHl9zBoVL/4KdFsBu8BtR+Qz9X
wqv1oD+WE6C0xTzmEBkD+NVTNGZqsfTUpcOSoM6ARyWgQqD+FdaQ7PXpciiTydcWccTywaVzvLrB
pK3+/qJRJ2mg1J7lIbZZWl9LSMwfJWcTH9o6LGzUWrRMoQztWLwhEINVsc/vm15DPRckzQx9mOxt
zHJf+1xl2PMSr6CXWm94ZRr79Y1yaSI2A2GepEny7f2jm00OmcK5MzKM9oABQdTGlGskBY47MU0a
DbByLscu65OWRXj396UF/nEum1rousU4K/Hju7iLZQesZV2/fswe132cbqVERB1Ng+uj+M7xRK9+
zUl0ioILLCUjftNETdgffGGrXv3lcBMIL8EfyUqW+NsJeao3/2t0r+nNT0eF2cwwXcgvc5j8wLq0
fvA9ayC6YYlCg+izpig9bfAq/i7hFAUSsA+zAoD6tZNSVg9VBb4jBFjllo0TIbVRBXcc1BEjpJzr
0utquZCp8pfw1BbFPicXLBR2fZlJ1xlf2N5kSGDD47pXn2BWUU8ZqLHOhsSLfapQsBkymzdOeGn6
85bdu8osbBTkPkVr3IHZpjT+SBGJ6wSiTn4bvJhJlW4Da4lhGQpUzNp4hIn774zKje80lKISN2u9
i8Ecc6NpBslgTwhu6K3nzpnDnxoYbTppa68IDviwuLAXDOdipDTcVR+yP77u9KRS/tH1YsC3e0x9
mbtVHLMO5tZvV1uqjux6wwXMq/spKmdQG7L69aIcZWLZIEaCjECh5XoSBlyqYBdJHgnti2BnVqZd
HXjZPS0CyMssvJ1cXTwNSQLQKfrNaHvzckZMEgzbq/OGBoL0dvU76EgUkVZ5ygFub63N/diR7jnI
geUokn1gAa0dnr2T2+MpqOWmL9AncS3jJuxZZ6Be3iKj3Rjp6c4wIOSRc8aadhIC6iXpk6bjCMDn
oDOKOx+zBhEJJIVXX5+B1hPe98WIlWbAD4skcXBkj3r3bCGgjuB4S/GymAt39biLACwqykA9g2uq
MAjBo+8hjPvYIjBsVSpPWrMfgVM9ZLsvkkPRVyadKvo9hEPzI3xtS8rkfUorvtOgDL90PR1fwq7A
yQO7pof12pFbNnBke/ENs2L5s5vwQks9inrgDvPSDr+KkX4P9lStJaKJrKDfP6+IKSUucxDwNXTO
qHPUL3ybVDehX3sV7GB4u8VbjFb8qx2X6KH+DBdChQaAF3Qsz/2HUZJniXQnO3e6QMqKEuT/0VlN
0e4RMns6phNdrfLNjFaFOVWzGQVDVuPDU9O4ppsU7VvLxvazQN4AjuFrH0RCeh/pHy1tRjADQ19h
6n+ijRSoR4A6fQSbR1XxU5eTD1RcRyUY0lidD7AQNNGzKO1YXgZzSa/W0aYM+Yc7AQ6b4PGzjao4
h0nKer+VqXfPhe7gkgZ5CviE60XOeRQKm6a/CT9BZznSbuOoKjq2gupU82Vr2KgOQPTcH8lWdYrp
PKoRZtphnd0YRNc2fpgmrIqkm/+93SpRlRS5/HerGnCoMeYFLjJ+R79GnEhOHkReBds5ixbqwmNK
BRMBdokL4uhAkzDSoRbd/KrXiGLn3cvAhBOR9D6KoT0B1fbl0QraPrIw9RhbMlWKgfi1eXENt2BN
J8NKtRkFZ+TWcMoDsFhgKy3IuiaVq0fUaLvFwGRccbHECB9bh6vybkF4VaiO32vrQZLLZpDUZm7I
dM9ZPNX8rIJ5OosTQPDR19WTpW7vltnO2nEgDrzxuOChnRiGAJtQmHaZIySXmhzPcn2eERL9IjJE
mZ0LVLCr2JYdTnTXF1j9MZWtRRCvXSr/gH9PebmE5Sj/PIZD3w+UwzugJNscp1mOgzHHe5vxOdxc
Nx+t5YfGrKB7wA34k4IWelHzwX25Bt3MLOqWYtk40kriRtYclpXF9Va4V/v6qYZ3NE15OzfzbV/I
KdPCuBIMzFGDJZ+omt7IszNYh9L3joz6S+gW87s/yBISfgonCuD2HfpnxLTK7hJDpzn/TVwanAGE
PdEvyJRmKK8xFxZoblRk2KI85IipVfKpSvzxV757AeW46CQ0ok0q/xWJqwDAzs4Bx29pnKNn+TPt
GqxaNGdDOzX+6NQh1+b6a/d1MzdbKUnpJ2Y6/JLQcv4p3VoO0I5A8k13Qi/zlgfH0zxi3er/PLS7
HJmcxpp8Pvzgj38qZG0pfOWNwYOzT3Qryltt3NrIx1xx9VYJCA70a4GgypjUR3YKzqajGOSeKHfK
rBROQBLf8jKsOMtYCb1V6a97gC30oZPLLUN05rrGvJY+rzCNd9/Snw8IoEi9vmvOX7qewSaBeeIc
xoP2gRktXuKqoK4lyB4mVf3L8X9sOyGwi8sTAeVLk3qHrR8UXFwdK0bFOV+6rRqM2AdQs09vJ/h0
iCNMYWU56cpFEFf86Ur/yeC+helZoA0KTckvgfFwDEPvO2UFU+OQoIDhrOIFysFj2+igvI34L5s7
Lwz5iyOVuSp5YCtvV7i5vkzQbKQr1XVgaMTPxhdNli50Yqd9od76S6dVuoH/uJDNJ+45nM/QJFhE
xSznuwHPUTTqjzIx2VXG0SZ3K2G83jeKVdnMax+3ulox8cpKN8QRNO4B2f3J6v2So+A/0u1OvaWD
M8xJwZXiLOrIQxDFmGKdgixAB8mFAgzaEuX2FJBhLcVh87KF6MK/v4sFVepCLfuCMJOVjnJP5dzL
spEuXQaDjbTX56bHfAlc3J0j5dNj9j5lj5qr4UVgWWQox16BKXpnXCiqzOgzCy0jYrXk1hdlwbyR
I+rTmXGdTcPcrqKGr2wUsbGN/1gXAQZT367w6lEAiNVLOgkRBSN6vWybgxKa2w1r6hOr+YfNSUPg
hO9TWCO+sut61BSfcNI87DN6BxfReLQf+w6KcLVRvJCSaGJ+ShVfwdRg3LEoLsWPC2V1Qq5hUBq8
uD9fk36SMoWUVKvY9H5/r8jYoUrbNwNSCDc60zCT7uiq0pOIs6Xo9p3qnPqGBVE4H9p+r59zpQ25
x0vxCHqfJ+WFWRU1coZwZLP0RkvmjEVjdPgUDpQKRw1chxs3XnQs1dOBlINeUiKtbzZamFGM1st9
VH27SSEKBizQlpmtlfOQeoVQ4u6HbOgtZPcGtMNnQsh/A8eJbQr/4RNls9JJETyXuh5rdgYSksp+
+h22/sH4UpVdJ/pDqF4T4kRHg7GChc9fThXsOOvJC6nhkOQOld0ArypYDG829iKgouMSZiJkUyI5
1H4JEJut8OLcX6MimeUj/Clg2QCD3IJ7bN5FiSTojoT8IO7vxIhAxLde0xTgCdWbt0IneXoaVz/q
cY4TfdrYQqEt3MYwSNFpiYGkbZWm4+di6/W9nk6AUxryG9YlBO9NxGcrthlMHepVPZ+cAVE8fDKu
CS5N+wQHagyn+Ihyd0lemuET+94c8LHJa5cbo0iOXfSe2Jkwtgy4bA9arowepA0dNJwSxaBdtOUa
ivW7xe4NeIGdGCd9jmpRQdB0N0Ufdl3JcAs38ALjwdiQI/0pKq3Q6VxvempRolv47Yv4eWhFXkYl
fOlcHAJuowIlvWHW7aky7F2Ht3Kc0DAIF1+3+tCQFI7KLK6tTQ2iXfI9JIJL51RZRs8grYXjajiR
qjG7G6n+5GGCQ10Rs9ciuupz6eIIe/bYMY+nAKNrWbN5DdzsTrwxUmYHKUDqYreXWxJ4UHH8Q3ZR
yT/BWKoIeFDYOEZyH4BqAaxRYefxY0F5zjmuj093R+OE5I3qFGlEbKgmfH1YR0uFWg9zPhaacU4o
y7kxKlvzmdMFJ6clwSk2i9/QZGzJyc5JElcVnGac8ThL77LHlqsbTlKSYIWvTdWWv/hUMACDSytk
rndmPZU1VPlnVB8s6wUoh1AWpIg3IbBvs1f6+emIwrgf+9e1X2Jd1e6vcX9Uy4JzhVyl2ntEcw2E
ifW9Pok0Tu6m+e2PlW7Rcglzth6tz3oYFySTBFET5JbfZJOej9KnhjD3kO9+p3uFysEhEBqw02uF
YwottdaTZUREaOvbNlk61tc5+vbZCjsD+QPDWsBIMHPjtwwEluFeRlzaQCpi2J6qXEiEgSegAXy/
a0HO8s3w2q26seLPNv5uTMRbf6NzhY26vEjim4lRcWsnpp0tI3y097UVm0j1vMGKtW7TE8rv3s+R
D5mPJE05CNuLZPSfgEqv4/E1anqHqfpRX8n8G1xZld5BPaFfITkl1XXcVKizU8jNoabeJUF4cL7v
LZNSWprhp6C5pbeiwN7iRWPDGykZDwyy7ZQT+eFL3r3MvN2W/psT1TKn05q6iOQT/7mUtGpgJL9X
3uEo/AlVUgzN9paGXiLLIq7laZpmn4xEskdU4faGGwwG90suNE+vJSSbX5eTQsGCDImcRK/hk60F
uUxUEKLA837lz8hyLwyXY4LA+TYXBMYnv3JShV6nnBrRuiFF++a4nUWBvVMuIaoc+RhfSPJX1doB
fEBCFttNto0u5bYotfs8ATrPMeMZIDr0L6tWzzfxuHr2GWqGz2sYONGjS0eHXzITiudz+jIHzKsC
9v37majo8qG/8NjhWba8N7n/P37LQ3bVsW871ptShaX6UMSgU1gNZ5cJVljY2OKQOq48ACFRbCu+
WTXfNVvWrF8TeaqLzyKc7xiRfU4QR/c8sGUcSK81hx66CGg8icRyPJ81CSdCtiXLYYjzMaYTDxrj
+kdS8LZ/IFS/8MHJuaFkxfKBEQcbi3RrLGWvdjNhsBcCuBTbpDQi4tr6qh7fmfIxrCIvJl7qAIhl
E1NrP8ZTB5ev4U9W3P0AqZiKWBkVE7zFLol27pGvUDsisuQV4KEQZ/rMNpIjrsPg5sThsicVo18L
Kpt+wM4RwZHkBOKX1uezQ4nDujjmPzFtLVaqk99Rlt44wcVl4WeDEHcpTo/oP8gWeJMXL4m06Odc
H0LKSpjzesSkkvR51dWnWksNDFPI6SRKrlN9OKoIl9WL+jXrM+EczFxiAOylJg9J21e317sPad5T
bxW34SMevz2Kk0aYIYjKxfs0WhjdI81KkYq1nao9lzxxP2muG0oiZ0tYTriyG+2fZawMu/U1d8zl
81qDz5mpEYvRTLRubjEmfMId7nflFIVPjA89VmNgudLFrlH4rsv15/3iuWdVtlvp792qTEYdf0JQ
BY7kGA72ey2NJ+pLpkeSCCedndF1fEibt8pWTiiVlyIcqFZOLnow6xGXlobXxzixxGX0Qp8+NzPW
BlmR1lOf/JP4LtcmGha37UlmK+LKv1Awj7Yy1Lad2R9LIQm+4C8paC0mOqsdzqppjK+Y1S/qggDQ
6rUXjLreHQcN+z/GswzKX/SeUAjGFygXk8FSwgJEse5KapcfDPSA0XJv5dtPyiwVLNWLY22w38L+
ieyqU5G8apRhzMA6zOg9PvarGQjbFalyV68hX1194SQYEIjpkTzAH/7ZSzzME3fO89wKj9+8ZXis
Bnw/JHFerpe7uVRKgqSGpPCA+kNKcqVCiPwYc9JZ+PhzaAFmaiESpZLSUUhhNGh+Dvw2dJ5ULQMK
H8XK95PjNKpMZjRJN4QO4Xy+1XjRwVO/oIDC/MJmaNyq5mVAo4lE6pnTqmRRkB9lRwHmOWL1EwNy
nyLMkXJzQcoFpr7YOO+NCeq2v2bUXGB3BHS8dN3ooL83coUJ9F/m4qraCBNV+V8dbbK8LJppZ4tp
kVMBzceorFaTe/R2beA9mDkx98aEz9E/smP3Ef4zF5RIaDlTwCaZ/06GVw8zTF+IgBJElkXNAifD
Yt40953fRaAzLHoCADttih1q8GxP3C8lxXqfwzeg7GBQ8YcX9cjAmMpKy4L+6mjBCyBtaARKA04r
F0swFK8IebZlApGc9Oo1rgRS4a2/D8KETeqVf4akNGIqMcuFPNlZsZMXFnGV/rWPCbhncJsTBOOq
9GfqsqzFRNAoLaOSXTVqWb41nY11yM4B0xi/RpCrXzagMzxqyo8W8LnzEJe21sPR23J4HojyFvJa
66DSdC8fhJK7x3vmw9Vxonp2yMYit5Oogbbz4zCyMNqWSAqPN0rnU9P8fYaptNwLfkEbfsXQL+2o
yP/A5jv5JKD8CmaybPpsOjlXfeJBJ9i4N05jOZOf+Z7XuPt0ftU8zWiQTyvLDDpQAi+nrZaD9ike
u+wxCslMfNfd0/P1QuOkqKoVHKxryKKE7fiRsmr21voQP1loIr+H00vMAEn7KEflbnhpi4o2fKHv
YCKgLE8gfEYKPL1MZdqDvIlzJTyZZQX7NscEWJOiLtoiE6tMnhPB0R94m5tQcidbO2feMThTFwd+
s3lNEjBQG5ArSLnw/Ar/QrZ/IN1LIYf5qjnhSiO777MjlHHWwB/H1lggNzDK8jq2JrLlmlJQ+dPk
/q02UFdZhmGRy8kEeUmdytNUW1pKs2pNbWkl7czD9E+K0zkaKPOmPrKv/G7frsBrO7IKr4EGf6AZ
ep8ZXBxS2Vos+KoS+dHBYcQHNJ1IUDrvWh4rLyt2Z1I1+v7QSzra8AoFw9S+OAcY7RHoMVK5jC1W
r+LKea8cSQ0kRX3UEPvKmwp+y/4FlgYjKbFVKqiX86NFeNnvwy6l0N36FBmqRtL3w45MLzRq5/i5
MxT1Tx2juJZjWyxNnaxNvIUtDIi4vY3SOl+lfHphvcg4JnZ4V64YOOlTUzsbUPj1vuFuTFGllyN2
68iuFIOdlhgt7AN3tdGYAuohONX8MPxDJrL2QnNKP8u8s39S20UZhMEQ50bV6u+xnUTmPBFq4PKO
S6b97ChXF/9YiDoXwjwBPjKDy1OKozEiTmx4ZrZqcWCQ0mJ0G3zc5tLDEg6YhtpV98Ro8VbWyE0J
wB5XGir6H/xZ7hSlPWJJAq1e/BmhR6buDT0bas60RcEDWnM8MMqMD7LJufmBu02iSCwwuOkhyLzG
v6OLKTepy0uXlZgaKGNIcn3Y6/4HrmCaayiukYa++X/zqfcOgK3Mazk56K8BuLvjo6+giEZayo0+
ePwNC5jI7WOm85y+ppgD4JUvXqx+PwzwAdhxEEH0BgygdlGnV0tY+nV8d7RTQR+vmJ5eqBl8v/UL
sFqSmgBuiiuXojmkYK/IYA9hs6GCq3QtRsX+IAwKE/a2znvpt+W4Yt+hnz6sw7b7QHhZxXdpyTkU
Ho6gD9cv0550I1vOIClJ/X6x8oFLZEJdVvyVuZWu2nNmMvwdoJcIKsQN39XPdq2oiGCsE2x/jexp
28CcJaxIovSwwaP6vYFarJYWvYQZotMZNfwJigsc2ILVS0qXa/l0wzqir3n4ZKUiXlHtRpFePzVG
n9kqDUJi/DtjXmWB+U+p9/3OrU1M1zVfxlcBONhoeR5wDVxqK95oj3C+9H8w6a4JeG4xBlUmUFfg
GIF1YDIevnKKYaOoWBFtQ+TYRjaCDR3slXOlaR7BMiYkNdFJsYZbY8u4AIKCGpthjrIAGNauKykb
W31e+z+jy0eyABaytOa5p2dmEA5YGkg3CUE/h7xWhVeGpsdBrxTPkfC23qdq8kdO+qjdJaCZ7Mf0
+0i/mi9yu20cbeGmbxtCdlx/3+CF0NmFM7CvumOZe8IVEBF2dxFOJ/aekCbZ7bK4fFC9Uh7I+b6J
DrX29w5ZKY0oypI4NNZyvIvNWpkDdF5MTUsMPnlS9e/i+dJ8AD6IFr3bCAER85YvRigGg0U8Ca/M
fWM7Fb80b/xzruIkhR07IB4fecM8YVWLNSrxhHAoCV9vy3/Wb18Pvdj54Po+1fLLIgSmVbOSDKsw
8XkoBX6AIig6WKZrGKpz7Fw52rNKKHnGHYJobLMHxuYbiG1/RjpWgB3IGwo85LDHFAvb7WEK0R06
nygUyImk5pDhTEkhMTNXPZa5bGuEiEnYV/dMrAWv/etvdpPaJ/ORaWygHypZ1cak5GTyd/81ewiz
fHT9IX6P4BbUMVCebzGgLIczRfeQW4+c+NwGFB+Azyl5ILcYH/I2WUAHidSW+1zE/sTV8YNG/Zon
i9eqVPkE9OkTxzhz2LU2JoG9oJpez0BCmJxXf9uqLrXvB5YRbIVP1R/WV/rkVflkM91pI8zaO//N
OOp5X2fVxXv/lVNCGyYGMQclauN0IcQ2Ul2j8IXFXDtQR5Tt5bI+LhEQ2/xbtupK3xgDMjv9dQdp
3wnWbTudVI5uGxsVJz8A5YpkjkRCu8eGvY93CqGQTyc6V51Enjr9YImgL1xXyVnJ/BhzCy8x5b8S
8bBQCoGrMyfYNVHzB190VqBg4rQpFCYyifXQMjaHqFMr2q/mpMmPVNpIYrSyTtxJdLj1ot7EA6KK
5xF+Sb3DqZbDaopM9EpOhKUnJj9b5f7QG0nHoCa9Y5vBY1y8foB/FZDVY/uqDVeNP2SjlbT0AQ5N
l61Jbh9X/RROZcicuYtbrYCVmjd8v6hye+KzNMLuZ7JHoO1ie/+ynHAcZi4ZSYbH1iM7gnbUeopP
ZPTwHh5m2gZts3DJjEfjj304KTkKKpdsMPH2vl6lPQg/vM48sNkSOaAJUmAFJ32ZPDVnPuEO6hBV
ewrRU15Ai45UR5g4X2VlqQ2Kc2x4us5NQfPEZ7F2QzR3P/RSq3+GAmOmxPKI+1x2MF3dsIv40sVT
Ub4yUjJauoc/0lYF+p2DgG1zqOUUyYmHPMN/Yp3cS8kYG3qiKMJtr4WU5WfpmGbGuLw6TzHJQH1p
08675YX+gBeTHZsYVPbahUUPkm07laEjDmLy0RruFGULIWVqULGtA4y6HwvnMbM5tSnb5C9ch1M2
4E7xgOhNw278pW7CN/uayC13kgCrZ3PGkbASJhWstXHUUjG4xuRTYlSWOah36emal/n6kAOX7l5k
bWHwes0qwVJFKvOeUQzHikBaI0pS2OHWwximZCaELzilYrzDeiE7TmbFc8b4Qy5gqxHJHIOgavrX
XbgchatF7UOu8lHnN+6lVhsTxf4O9EG68WntY5MGKVPuTu43dpH0Ur66UtLiZMoGqhOA1twFX2rA
RDdI9oqdVZNI0dWuvMe9rmAcBnLwz8x6VmNOYKUVbQuTSsVmiQBg6WG55WoL8voAWihI3ukI7c1F
bOn1qUu8ltxxeoVZ3LOMn5uUcZb2v6c7lfaEv+G1aIy0T0eWBWIDNotjCU9QSEt3vdtscJl/QO4n
2v5S4BogVKzihWh2MTHdudBiN4blzUmWVIZ5HDOWxoGJzhMFLWIdLZkTUp+Pm4+8p8XGYcsD8kXq
nE1k4pXwWuyB2GSYEEFBzwFB0E9OQyB2qc+ooiei1PRmVizpnA5VsuoGkKQO4L3/UN9kB1VMAjaK
wd6Kf+OgwkkvwoH7LAWH7b79W+bzsjK5lN9DKwPDWjj5rWZiKfH1pRYT+1d/4KcjJsPX9uUs8OSU
Bw1ClODHCwLr7a/0S7cEvLB8tmOvCu5jpI6JpEG1NFHwUxa4PBvB4FkgERRN/x9HLCysrVSJEp3A
WGePA5bFlfJA9RvadgP72/eehQkDH/4p7lckILom8M8q9z3CEJBoE3Ujn4zWPBB5G4rA8l6+nOcM
zlm3ofuHINtTWqVpgGro9UGSeS5RgAauF/SBMRvlSx5NmI24yEA9vdZ+owSHRPS+AFEyVex3zFbi
KOW/QjK+7gKoBh6F+Q7ejnSOJCIejF5hCgtcriLJsZCmupEfZWhqtrACk+wbx6pXQdkQt2FFUadx
OKbeV0+O5O7kouQayd44LABvZxHiZnuFLNdL5fPLsaZKk9TlPG/bPSiCyECAg95YjftOCcybpIRr
c6Y4AeEAwV2KCIc5vTDbY3K2Vc1Wq/RDS+EjDGZthpsRMjSJhpq7OkfKD0QLKL9vcsutMsrwN172
CcGMeqOvxzo6rZL9VEp3pB6wbtDtZbw8ztHs1qwikyyjV54iago3oOXyHGUJIVeurfTo28dgtxHV
Ll8U1z2fWAhTwKrT6MiJwIOPm8h3A7h4OLwIrF9YBllvU3tV2yGPMCeMibXrZfiNvLDYreRZ53xK
RIiErTuJVVdxOrv7LmuWBzxNmcxxTXy5GdTTidmByynY/hbdoQGP3DcefLqsBaS4U4uhrvGdhwOf
fn80gDoEmxKyXmFs9koIQkx641LDsCylY/g1yxTUkhRcbNsr6/XqmXe0p7yV6yAok1x59AH4wiMH
L+0HHpX7IRH9q0cTKeA5eLvVPjZlu3FpeHcx3COaE9WUZ5k+rYMN3Wxgv2XOldl2+1a7JHzjvdUt
PqkKRAV5VcEWwaRvr/QGNKz0qdReOSiihZWUA+gc60RiQEMugANdzbcXcaMpUS7YLwp0Nj+QtPUq
bvKCA+/FQHwu8ORszhsK08jQrWWkzJVDWQYrVK+2NTGqeXDP9Tm+XZp9+cUizjDX44/py+3XEuWe
0mPLmVtyO5N/29W12SWb1lmfUwA8BZQ8q8zm0oTmtQblTY2uXqfwpEBpPpso8cJA/1pB4YAtvM39
IZMxaDUf7D7wxrEJRLN7OTZxKcKDSTnqYCOanrAALfdQJwjgNePiTlHk2uRZanmZghIglGcujG4r
khqE5W1CZd+nfT8grpvZNNcxvXDGg2DyH+tx3NivWe2723ZXmN5LyxcNqgUMbB6J0lcf1IUieDMY
X9R7FMPmNAbg4v2zfPK2va0iVMWQKjmxPbv6c8Dei/R5VhAz3T6xPvUyk0Lg8VbHK1ncu6JHs/Bx
KQ5g+fMXb7CBRJDGmKfAkqBzLAO1b9Zm8vzkFqz0JjqdCAHV/dqEhbhOUSdBw3Hp1mxqeOVFcQdR
KaZpJxJUnYP2IH+lvb7Nn2KT5eU/x9c9N0Jmx8TfpN2zxz1IvJzbGpMjnzsP/LiIW8p/n+93YIOv
CuDvcKYXPa/zVFGkCYVJaVmVgRfC1x7NOp191YZbtPasM+SMW7w8yOqO0othjSNfam+TlY4LHaI3
PtzRX1jrPBjnBG9CRRSu/RDZ8TSeU+ptKTmaWq665ww01AKFL25XksGpaTBPmGnYmIIuJFsNo4r2
G2Xu74NTtRG7BbamWO+GUggSCdN0QVH1CzB4FZomjDNkDVnfSy63FS001C2jkdhsNWeA8ZiVG/1Z
2pAbS3W3mvbpEpCb1weNNEp6tMzJl06a4VvZNSLngOEGFL/if6L4R/KoTK6OwXKKa1oQWHwiqf9p
ZBtKVFnJxKrsgb31fPXq1ozAcgU5nZzK/gBLkjmPSoFb5vf3L65bdZuEixSAVmrIUpM6vctG/i9J
7sLhChMZ9q5uA+YnTtg4ELfYgTxk03zrNE6vYNfi2zNw/pP39MYU5miYpcJTrVfyGve4yq6k6f7x
4q9MblBT6wIneL18NIquI8PJqeb8yq+EIFkafAglsoceIa7ake7E/zYas9uqMj0zWaXhxixR2buR
piOsgso/j3VuxEkiEQz5sKdYDohgs+1E6uFS1sUu9NaYHEGbMbARtDJwZdV24iS4f6MvoANz4VHb
PZSVhGdAwlrI09xi803shvWOvn7+NY2snLAZgDq7kmwO++yHx7yIwYkFJWMNc3UIQPlJ7DX+0Mye
3agF//1+v/IQN7tO4islztXg1A25r8ZULbsQM7Ze0s1ceUiyGjJmH2vKJUUWk1vF6uAntI5CA5kf
lID5KZEiKqpHhKxRWQAaQI1SBaGnVUQAjMm0AL2mZTU4m3LG/bHnOxGtQoYe7dqptM8+l4htGS16
EhBBxApXxXKrozKQNAhZkBCSZt1aEpQ7iYW72ZPY+K1sjJnIztGi6YfSlzmZUh2Vvwj6C+JtFa60
RbLKyA6lFs9kz2U1aYV6/FSbU6GFZ4B5NQp26Z0Vx8WdGu/6KpKa1MTRhbiuaEI94w7Qz58uGL+j
YRGai9U7BLttYJjZ0t6Se/xrRfajnQfltBAxlg6RJebaCW2396ftJyyLy8xjAPDQVnDW9KJjRobv
Z9MR30vpyePGjSTck++y+WaeT8mftKn21UB9y8V3Gp9+HnlAWzLnD/gga2gqo4dAD9G9QGgrVsh+
Q0HMd4sD3vF4E/JK6joO8NlznIR8U3SictJKRyUUz+S5fpv60/VjnHz+6ILkUOsvn7FGrJlObNt0
lz4vlhpcDVZaCVuC17wcqPZXpV1R8tpBLJlOU/DOjhnABQBJYniX+v5WePo8FBK3r9eUVh35CChp
EiMANpluYLlyfesFt3Dw6iSsYfdZ4ipX9dAD1HaRcUtRLQ0JaNMCBE6D8+zI33AAJHS/K8v2qzTe
pGk5X1nFINHaI7t8ubPZCaYO9MCzJnemwFrlozLir7ruhTAY24U6DvEmItkzUQMS2AcGB2pFeslT
H+UjYM623Ep2E8AvoecF2yTt8+cHaMPN3F2p/RNvm2kHAA66BiKV0vP6dSu9pzBakU7+ome8GD8Y
sEPYtxAOXr+LAzuyo4BfFQbj3d8XdK+OK6bV8zaHqttDn5aBcjVPZRfl0vubtIZxoTotFT5PfrlZ
sxO0VXNC/U5ZRZ1BckRYOliog/9fOJAr1vfZMzl4J5vdgtRqeukiDGvHYzdbIRj9hrMsHAnqGQtY
fVkOmWwmJTPkyhr3dWH1ZIaGOGsKDMJnh2+F1CScS6jPal+HbC/+RynLUETyb/Kkxg4MqqodgH9i
9dMSX5YGnfy8gSwaCGQWWHX8HI4rZlKmnn1U3JN7sOJXmv1IdZU6TlJMneOvDZ7raqwQOClAfo44
IULiKX2Aob0J+JkJjfgN82CeqiBdMKnJciIsD0Dxl1t3uEGwDaeqMiLPsrc3DkhJIA3b/6snSvSm
jmkkL89f9ApBT4Hq2k33ceEmKPi+sYKQImfNEYvWQ3jDVjQ70+FjYK3zb8+2yfSPJWnzsAdzjDAe
a6o3vSgvDvNx78w4b8ikNZxxkFPxJzXO8IeUkLtYzVXcbiyiBdA1dxdkNUPJB0VTf3xQPRxu59DD
htIiYvwgCDSxvtWJyH9RnWjS8GocAxjbVHaoIqVeSUPmvjAafZBwAkQKUwnimAjExSi6jhqPAvr0
mVKrDP+A5VNFMvSnNVLAVFkylhsHB/VhweVau/MX4XfFdLiL/KYRatG/yRBTvnjojqQ3ejKwYPyy
9eNN1s/NjRqDsebXvzGvDAvodre+KP3dHC9h/n/jCg7Z4rSnEPsMrxJ88S/RKKZ6BIySpMMWmhkL
gpTS3nCxgqVqDBMcw1zEP5pHANXonH70O4bGhqSwb0uMN7vUB7qcGAAT++riP39i9Az/sDpqA5oV
uXDH+6BTq0voJ7UOei+vIr/8zz7eZubELnvjpNAjiVroNw79Q6ruq69tG/pk2vkeKOYDq7h9grRp
2Hc3qjI+ke3b8HHcTIYix0hO+t4bxCI8kPaBks3iiISrXq1F1hgieRAGvjhlruCtpvHWYw8rLc8D
IxW6wW74l/HOmnhEArAdXxZx6SKjkGSYvuBBsc26zS2/I0VkI3iCYnt0rRXUNmCNcgvHLFNsemJp
jIqPauqz8Kh6XUbjUFv88rgXywAd+AP+PZpcx/Gl1gfHtLn8xbyD6nJhfevkuoKdYuLJrzKmJhr0
d3dInCO+a0p3QROIYSIJDRulnHMI4nFfwzsmxGX7pAFHA/l5IxRm5C1LZwN6s2ZVkJHkVSIoNUqI
tPgx7X8PZhYd3yi3dQ4YKLHAOZD77GzYNZOBrNlaMxQj2DSyxBvQpIYUIPQRABindG+7zbcWMNoA
8fo0Vo2A/ki5GV/KySZRbxR3VgV9Gu9Zt+6g5En6u+8R4TBMdoIlP3cLR0s1QLTPREM0qIA4AhHo
fGHJcQzwA+9BJf6uNIPbEOnE4Eye7wtuFP6KLCxa/6vUnieatfvKm1u1KUOhqDghaP6NT5ispkr8
iALxD8VPa9dvKgm2bRgfDFmrMpWoHm7PRYpqJktd5C07oLoyKdH4NAUQtrweIeV98j+2rK78bf1F
YeijFtjk5WQva9w8pF3YMhZGVpINCnEJoebjyvglMQxjMkq5E93AsC5vt3w+UdfbYe3/3WmWFdUa
dHSjG1rJCAkaZ8M2bx4KK1652Oqxq4+y1RRUi2zknKacdwiL0ozdcYSWOsng2S7lJTbxl2o8v94c
xfBfjw4UovXjKbo1KAuMJRfpZx71+VgojTYtQmybWaXqTgvSDbjSOM3BngsR4vBUGd4E8iXkCm+6
EcXP09jJUcjkWqX3faZlLM0oQwtVHiSkMJxAGyyZvshXCZrK4fhJZMWcU+Yij9rCc3UPfKVtrr4G
QkdLZSwfVdr9ZdQNKAVSdbtMdmoaun3L9gTiJGutm80lOtoboZvv6MGh/m4o6i851Q+lIDGJlGSH
UxYMzMX/I8AJlTUXfK72siTEt7c9061ZMs4qrAuiIAWT35+ADS4HU2SrQ3JvRYzih6OJNqpod8FM
XxvE/jZOEYOZvaUIjjUMubH4D6jI+qvf+3j/2vlfyTDrtrqEmA1jBxiV5flZ5vlkCjo7Qb/DZmh8
B2rej7ASGFX5VhU5W30Nf3cGWZ4yjkOTEyH8KJzVnCZj+UUaEIuDuiV7mzi4EIUWK8aeyXxm+g5r
vc3D7LvoG/9ehq2F7KEtzbkJrhkUf+FZYIrgMabL4mbbx2hfzQhoNnYG79Tm/87dGSbsNu2XcabH
nxyk71xTf8kMcm49OQoVSr2trLukF2vrWbKD/CvP73aBv88za22BT6X8j6jOlq6jXVca1LMaHArh
69FmUDU0IJA75l8mgSySQx3Zqceqsxpe+6l3wc7ptRRgZG3alYEKA7ymrjpR/yLwQm5vSm13x8ox
kkGgxMOFV1hZz67nnESyOHqlPr/tFTKVJdhsNoxsLjTVesuauS5Oc1vncDeUvm8irUU7C/lHTc6m
LEAl4wk4W444fCm48RipIWYRqzVSpNnCeBlzif2zyoUnMKOtxvcHPn2XtlqZ2iW1zGyC1gl3EqW1
Wz6gCtayxgcZ5qDsQEcn8A+N0wTwEouRCWcBAThqJ3NZtCdNB76PebJ30kA7osOuNj0IzaZ8QHCZ
hoeiuftlbrVQjgPdf/EojO/Y+oMR+/atzkuNFDU9S+7qSAapfX3Q/MbOKqg5YJPYBF/c5AqbnTyy
IiAzYMfzqQiJwp/QADaKalPs4SfJtzriJFWcaIIWP5BlZEo85dAtIgdPFc3T8pUlXf6Wbn3YTKcA
QVOshFLSjsAmMEWIda9PPUf+wLKn1xHCkTK4xuBvtj9FzgDVmwcxOTHriuh/5BbXKIVqX7CxArY6
Eg1tXoo+NRlH2oZ8LdFfxKZL8Ac7TkxejUK9fJbVooaE+SjaRUf/hk/aigC8jkzvDc+xDsZNfm27
h6qmbDugNHwThuBM0D2HfO3fClc11StcQd4z1CvaQ/nV92alt0Eml5+x6LYPvz6yovJrVLzQtH8+
IICo7yxH7c8cYofTj/OFCSd4EuaWLONbtI4PslPkQ2Q1JPIeG90+oQxjN7QaD+BJOURUJK8RiRSb
d3WsDNVuhntiSb4u1a1EpV0r3nUhu698JEfKXeJq0NTFaxU512vmIXnrSlegQDP4HZgc/Ku+Aja5
vdu1+gsYNWoXILDbX2ij0hhw+jDMglG/XaP1DdJX+GOylgZAihPr+ZpbHxPNRaF3oio1+ZynVW21
vI0H/PzhxopfDB63eHDDbB1lzvYmlpNJGmtym1r6RGlH92wk5Z4ng6esSdfn8RTDf/02vuROuq3w
IYXmdwhWSOZDZOE09wV619UWG59LEbBppmsKwEOGwf5LHxaf3pf7yezhzsMe+uSat5S66IL2ujJG
WehyuxKWfx/gin9VewJsB/HlZx+h+u69U0CfXavXsFcjfbbsDwH7WKk/TWZsuIqcZdzTBB9CTmbv
WIgNSPanEiwWW37J6ezBqZw8DL3H57qbip+zCmqqRUkgQuOfgYhSoWar204+L+e2aMnAX1clQslx
BsUH5GwiixNWUVPwVvaE1wEf5l6k904Du7k5LRJzlGLrbZoOHvnOJMzPMEXnoHGd5O+X405gKfPN
8H7VPVDjxBouJPQeiv71GUwbDZBD3KB79+l5gawKdMymLlSOkLfMlBfri7Yk8Lf5RLpEDxxKMHwf
zgfO/v/zOxxlqzPYgE+blW8RswT3Sa4ogBtaE6uQelLUKANjC6YZczeE/UcZp9eAWYXpkUKq1cRb
V9BK3kRS9psCbK7ytuJj7KwNL/SXFXvmRoYIQjKZRnWIZtV12Px17f6k+8yFXXa/1WOhGFr9IJaJ
65vh7N/rwWo+4WUslEBzn9ZnfBmkQuV14+1CoANHab0wzxZCRk4n2bVbmjrLzuQoWnWmVGhBZg4T
JutcUcPfbxUT4CVSyTkAIIyI3TiJfZSIVz15IofzI0vIt4u+JcxX+KiK7oTC1gsYat5XrvI+oryO
TU1D2VbvKj9ZZ6fklOMa7LJ2PfItfa4V1hWVOkTkvoIV3X/P9bZvMob1v8rHImA+Ga+Xln2zN5Mc
2ceAKB+kHsAUQQu71rLq1K17DBqPBBdGu4SnxUlpp+gUwtvnwGPcc2TbUtn9RhW+eo0BfEyK2l6d
STONmU1Z90e2R9Q75Yc0hw7giE6qcZtnPTJSYO39s1N7TE7Auo9u3DGXw9yLFovqsxYNn7MgC2Mp
PCWwOnvFNO7mbdr//bb9M33TVWPob2LIDO33KTk8C4J2FgOinOfvp/0Cgj9YexxTz2nxByhiChrz
0CzHOLFp/gQSylJBkEtx2M1Hu1Madj6u/Um9uei0eZVjHuYvwnOPsqspo+Ca/Xoe7JysWnb0v5Ho
y8Ku6l63QdJEPH8TYk/fV+lIrjMm0QD5+Pmd15yhdmmZ3IUzmXp8aHozcreCYSBS+ZjjMRF23gAS
KgiM8Har+zMfLpmmqSzF378d7XHfK3Hh7QcUJ3sjeP+qTsfOzsDeIrzapRHGFgwljzxpn9bfwfk3
RRE+YEMcy/cvrU03DeH/pZMRzFKK6Ssbgg1To3guF2dkrxwA/aWsZPATD5Codj3V4+4xOZ31VPkO
IBWS6+NeDt71JCwzgCsBzrEP2y0yyN+kgBAiqfHdj9enPAXyVZB/m28bolVbkWkBqRzOTfFyIqdt
OjbROr1GZJCiC+nnedk22xaHG721G6QTu/Zua4WykZGIz+UR3+YQcMYFGoTjwDko3JfajRATBrCW
0LJcixj0320ieYXSK6msxXWA67le+BWdMEABxkjjG32YifHXTAdOdBJnYPGZKhay3J7F8wFdEf7c
PKtj4ayRY9ucwtupzGi1CZrRCaYEjSJm4b2pQg92LO0WK0lmH09tG7tSKaKXpU39hw3wdHDZDVez
esTH4NNrBPVSDObJ1KGfEVoSuGFrm62ePxXkSz4YG398QpDCTv2St40Uw14DimnoYchuJRctuiYq
U6GStQw7VmgvhhqWTEIMkhSM2FBG7i6P313G7ggkZKykrtgHHn3UX9o0foFulxjpLHgo2ZEit4RT
ln++CP8myVCTsSX9TOLd+8zyJawhppuivf+NV4WdmSKvuitUpfTds0IgUBKRMQpB4kIcYggxGOIx
9dI1oS23ym1cktUGpU7y/4a5mKKkVWy42joYFlStJmHzwWJVY5YhvjHggGrLzYz4QBokfz0b4+eb
l4le3AmpEEOYubRCOOHKTQE3kQIPbIOiQts3Jtrcq8WWzePdlZE63G6evhjbSbngsvzwEUqxZGCR
BFd9SkkzjprWdgVZiIFM/6soCiur+5zhSbc6xswLgzRCZxwdLDDIPJLuFKh71TbiL8VMbxJog1Dv
15jEvaFsiCzMrAimdSAJram4y04STwHPGEtGZXC6m5NYjAIQPbdvipdC7inp4zRjtCagujB0LYhr
FfiSzK3CeRRsjxB+TNSAsnCZ0a8Y0YFAIMx/iROXq/e+MxD6IDWAchPsynLFpOCBdJMekRFenpCr
eemygdEFWFZQAYK+tnvH92AdZcpYoyNIYUegWExXLbu3T0iRlGIgBhjASUsCzFIr9xzKYojk5NDv
PkM00l86NhTPgrnvXbA7WWxP5GxwLjJ8CSmPGpsZb0BB4H5nF6dvJbHeeA0p6dcpstAhhe0+s82g
XXuJurAKgZ4IY3SFyeKlsKqjef4krdszuENBTTSKpYuPeflOr2jXnlpZT303FzdFbo8PGBSVAiwv
46AWoaR00iTLYGUnk+23YUhyIB49p8UU/DCojmoDZyeGtqGWOrSYNUp8a/SBj2xejav91LYjHdTc
EN3yUnoUu8dw85U/1C7hwfcopaZL/o2qT7uvUWMn1PAFYLAP3XBsHyahyl+9XVKkxQKj1GAVvecq
9tjibXfO3JSl2Z2spdkMYLrGy3XWbh75Mi7w7+GZouHE8ANRYCdTKeELo5wO/3eCpQD8BqiuXT5g
GB51AG0+U6h6k4bBSV9FaNqkjgbR9Hj4ORWXnvkZTcdd4qzyBEsoezCX450awvE/OoerpPgfgmMd
8/nsOEhxaVCm38eT/IzdICy/QJjJLYSUuslMjAbvPMuqVGKQd/jTyS5ykGxB6WrbulCrfE6hHu5U
C61cVv3MWdxfD4PV4PMq/OMDWE7zZN5eiNHpuD1c9hrJfRpCwBMGfE7JEdbkoMn/McjJjryAJ2cS
HtGyFfXzMK3TRw6LQXCAmvG0MoxKq0gBi1aX/uK2VrbvWMXb7K+OFymF6aCB7Mba+YrR6qC1m8Ya
+KKGUXNF9qH547uA3iXJX/ztXG862Jf9Uj2M7iDU0J7qfKStCKAKjft8BrX7JkIS0FrOX5Zt8l0o
87RI1AkdA7LFWCCeRlUPiG3WTNvr1VtptLCmvcFJ4qLYvjnOXXNbkbDKkhmW2/CGhbz9loHN0o8y
wj4Qc0HDlucZGyP0ofRlWBjf+Bf98kRsn5UYounW7Ngt6+cqcW3JSj4iM2yxxtOh5cphfAxp7Rv5
namsMs+JcPDewoLbEQjd9exT8cFoh2KUCu1OZ+lUnO8bUmlcKK3MMQVVNO3HpMhCYaHlahv9GTSQ
RyllkM5J+m0zgDBlJFQ9CjJyhbFLspTFoR+/+o7BwY1TtwyOm7mooCVBGi6qBmmq1iYBbk99LCSD
YsL5nOLT3lwMM251vYUodTL+CMuet4eF/qS+ccu0ElE4SAqBeMSfucmRhPVUqSS6J+1mXso/yRsy
ATBZXqNSKO0QrWSd/eG2n8UnS12aFxUYyCe2WwPRTzTV6FB5QdF86XGW4STALuPwSFbcUBa2cOJa
J9Vw36fewkxtEUbQxXy7d29IxHFLj1zq91zVqodl4SQNAeFJPT6PsEXS/OEDccbhYHeSw2Ha2/ml
NapUeUGQREBMZOc7OHUKHePn51DG1bJmljC36MvKSxEpHrxpVHmPzvNuV5748MgVI+ZnjYa1XVS5
OL28cV9yaa+dJRNsGAZ2ZcKJ2vmvI6cq6BwdlYmjoZL6+SeKQwfiglMsyo2VU5cG6AVJ/8iVZQ1t
sbE2pOud4/p9VnnExduvabmzT9GvMAlHg+Hz7V2slgVHy4bSC4kfuxufjh31P6Tzh1uoU5lzSFvc
CCSGXlejvxaVDLmKqB0Bo6Z5sibFP9hgVIbFd4axwwZhH5ytCKNaUFj5V3/WP0TA/sRVg0l5RW5/
Azvza21pLuXb7+5BNGQXre1C8TbltL2yXrEXUmf5Ik/fZtCQbBpPHiPUjL81G1AdmbxkTOyrlxvX
GXOCdEa1M2ILMYFdbftvbN/869P6NCgVWrB4+21qiPJodEtthtdhJCtgqQcqgqcnMk6PFGkwxcAi
pt6vIKYtm/2uVGFcKriRujk99jjUHEJeaGz92usXPC5NdfNyqxDraleMDDmn8WHCj7ZgljhafBPZ
NtLo1Yheoz04bXABuXoDnjFjjvPww7VdMpO2jN9v4g75ugRKISmCDzo5IoLi9DHocNDsXCLERKAz
/iErDJqr7v4l11mohTQRGEufgeOpVVJcvGWuzi70TIbmEkt58EeSvpSyNnitQDuWY2o70X9iW3sw
Fy2CVE3+GEcwm1oKngUlatt36gVpLIqHrqLQmFUX5LfpvWmzP7/xEqDlYuEYSyFnp4Zr9abul3+g
KNebe/qt/aBLD+UYhQHesmmekllarlHKt37n5bvBzEA+mOBR/VXvK7AdPTSWuPA7hJoIBKio98zp
Lv6U87X6+ks6E2EjTiqLPEWOp1myPnFWaI87A00g+Cs05HcMpMibVQD8DAd9zCLFjlVRt6U+k4nK
C8a1UZAm8QCVUOO1gZBPluf1D1illCElryJpuChexGP8hHSFSYIs6U0vyrbuZgdUoqZhS4Ha34j/
63BEjCMPPjzKnyDTvAJyJnuReLJ/cNyIF82oo2BD6nTiZPEQkdkmBakza25OvIC+WQGM/ZskNbAJ
7YqdAAJ3lfbskjXCdadMArGJNS0/tfvEBdgcnbjEZ90JgDMGBAxdk2mLNSChvgFxZamQBJEu33aX
O9ozpqCNeExFXO8vHZSeBPZJb6CYzu1i4HGl7mOQmx0YG8nJ7TDW3HsbJplDGkvjH8Iz5eC1osOn
C53Fsuts+TzVM9gIBOmN3CKPm0+O5OYB0I9NeefOduiKuxcnLPmBN1tpEDkiMAbwqkzOh6DWdEm8
gFqvcJ4eGU+BtEL0YzSNuGZPOCjea578EwHUWVR6E6kgLjXpx6y0dtd66eZnDaBcVQLW0FR+2OG0
OmZaQeo7fHGhiFVefrJHnjowL9bzM3pK2MKO0Z2tPar4i0/2w+yGCoagqxNrS109ZBTeUyKE5bfo
1cQbvshYLSoNcIrNJepY7JQBIqbeSV9RF3wC2oaIkycx6dYVZZw6PYRPkVur+0vHDu/rVQJ4Ygaz
RSWf01vwTio1lQnIVQuy1qpodF30jI4WpNKUjEDlDaS7oAEYlXZn6Is8RxfNNtzPPWt73lahmqDY
UEGCtZ8YkYHrQSPS8OQvtCSUAsoBzDX0qpboS0WYxuXqQW/1s1z6OVM27rCbopRpyUJpMNluovdH
1WolclMc0rcy0lpaee/DoD4tchQRe1006aXf13OUhgP2osxoTxZs+rXcZOtFqtiMDyzXOPpv2KsE
0arkZHjOYsRXJerpf6BpJ+ugCNqqUrufuQqgyog8MxROzFzY1nhGqmoXkGu4sweRGDro00kvkRbi
aekq1+pXEXVi8dLpBx6wjhj01DpivafShZibIw5zWlMcKqHMkZNHCz8uKqUZnWh89q7ljPKTQHDW
/yBP5TKZ7rtkmfaPib3Kg//W52Lyw7ipE4/qsrdoR+7j9B5BgL6bDHlrbkW8jDYaYNLxJ4X65CFl
GqjiSQwvVn4zG2DGbUkzcfnBjlpOmIrHZdaFJcWwV3ynbsrIHmeAe11Wox0DhYnBdvXKALzmgY/t
qV+tgspucs2YVle5+3r2ZvQpUVmWsTVDiEf+5H7Kn6R/c9vsp7T/S1jS1yDhxN8PLSu0FJ+jJamh
EmrcVrrPdG5Z1RqJsnWwYD8mnnFgpYyuzcw1DVdkcqogH8ottdVcMdeaPPFOPTn1B8f7I9b6wGYQ
2EMpHVki30U83nb4LqBdeX3cloOx5hk6yunvLRfVNzB2XfO69WM2UOLXMbovEVc1Gf8oP8l2R1uJ
YZ+SkiVOQ2+02/4Zm5h6/7ezmG8/KOKILz6CYRCgUvPfl3I1CSRg/5Y0XKcTQ+1mxe+PbLSrICrQ
TWCy4DDbkjy3dAWUI9MeqmALTmfNiG9eT2o5ckyBtOaNz5F0EC+S4gHjEYGgq/tf+MJ4fkWOoISk
uulVzQbojjREp4gEGfe3BVzxzEiJQo3GvAlC+gVYbHfE6ON47dnb/f+9qHjOUL7/EWwoiWVPt8Aq
uOxSse2eqCsIfPp54JfA+zsijfvX8mQ69pRAI2kk/2UqTaCD5m3f3LYtnrpvDIZXJquAWF49s0jr
b+Zj/WRpmInmE+79ScIFKIBVbEo3kA6OpHN0U9rH8L1RVZJMJvmQVi4mDO4pJsy8PwYl8rrzQ11/
kkUt5hxIyl3vkHYWcaKOzB4XJPt5teGKTn5PhZxN2vTyWvbsX8Eywz5UBMYEp2UAyD66X3f40ABL
dBgknB3Tp9kMorC5jSTRkUDNLNsdogiNscKMyfVnwbad8qQC8fcV5YN8e0OJwLI2Jn1A/mHRWfNm
/krd2RlBcT5ftTMt1Wgba3Ao/i+UjHF3uDZYIHkmZAjPfxN1+2CJ9SOEmqiiOPDBhXSU2qUaXkTd
ZbgevrccZERMT1+HYy8P45YvZRqq2MKYpp14F4S7yBVL2/NAeuPK5nQRY0lDiaYBEnsOTLYvVFir
RvVeiI+EpjGQFZoAnvQGz/m/s/XQrKJIkQ0x942h91fyMzUQKi+eKM9Lk3hIuaaSbbCosdpfwQZZ
hSwDFLcil8R8ngl1Yb+sOC2OIRLb38XqPu9Hn4ZVp/Y40O37Qd8UQjx3WeNP9UOIBF++9JNFlPfp
Jeqm1UztgobC8MS+Gkhjjq/aPoeRhDdoB9RbvPrRXYY+r1UHt0bKxvNqo8a0jjbjE1x4RflPR70p
xo+b++IgWLisOdt45bJ/Ck3oI6VWjqL7VSoPSvsZ/9OCzMMO3xyJD7hrsAAMfyw6DG6hujwq1/Pu
CtU6hFnV0Sk5T8uUGLv5JCWa859zj+xDjkLjJnJPbd6bG7UyEuoUOWvZCrCOjASjtTlQG00N92nS
iISJfvpNoLt8pI7QvktoClcxZ4D+MzO/d5RFgVAaPscVNb+39Qv1ICPS9DiITFi8tK/pK3hhPVs7
+zHMWl0uiPYJNb+ZTZIg+h+gHxMeRrd5b7RSBYwRz46qi1mjOSW0vag7EGlmsCyLhFiPT9u3WsTl
YRqVKdFhIbvo5lUuQtvAC10JEmZdX7iLIw1WAjTYffS6R3sTsN3kI+h4vA6339UM95Mt9mP0WYiQ
0FTs3JJLyBflu9vsNaN1qdBeCV48w6E0HEmG4n5zFCCaxRM7gN5Meb+cLVByOMOX1SyxHwH9wb8Z
Qpk0/GRMRLg5fxsnV9U0W9KO+JRWHvUYsv29oX1JMzEFcymy70HOR76WxZMkElbl72NzIaDnMDgQ
b1g+yNOq8+pTHCyt2de28E3UpeaO2K7ub0p8m4rp3hqiD0gI5WdJ5VfnEjvL/fY3lF8JzbyCiXzn
2/JUhdHDiMJVe5s3MtOmpqfi9hNubpyLm4/lY8/auklVEp04z+5LSL2d0lYda+mWEojN8jGEEgYD
4R28iFaxGpnzy25/swagalQPsZ7Q6QLUae2a9Qe6vY2u5RyWAEm3BuFwLBoRCgEw23Ip4RwXbtli
y9M4dN7N21o3rstnrg05vSC/i6YxpDg2VP0VI6UBg/EJ9KoM51fL24Z6kJM+TkBnZw1QZzhqM989
jZPH+Z5I6PZiAcgHbrJrv8Kj8o/72Hi8pst38bbux6nNHJ00hdwsdPnOnou7CDi4msvA3u5XdRrK
e5Aswld/IqZ6kL+GTxCytCtbIMUfUPMcAYHI/qmPVDBMFHx446ctyzqELFk0N1c0I//S9CqNSo4F
17GDjNxmb0FpbX3t50RYj9Vjjw8yJ7w4Pz5WMgQ+D9F6gSy+gzLLpCD+0QMJpjYmIzEItyLAnoWR
qnbexZiSFXQ2BH/+TC27GlMWf3paaYtwNKeNZD87a8lC8+mApJ2LudhK+tNKJmmWOdNeOsNm0Y7K
U7IRWDD1hJ+jNz2Tvj91SieFrazkMhbN1YRUPfFKqzQ93e4Wg08b4bgb2TlIHGLnDn9MeSitszAX
Yy4Myu5/lFya6bi7osvJm0AfsOMfIEXDPMI9gFOiNMRKkrjdJnJ6WZTBAsBDqEyOO7CgBrNRFez3
tLj8PuQjH6yfASLHZK8dumyt9qjgbalC1uNl0ky5ruKXNrGODFu85Q0oFA41CYE4xAjx0kMGI978
uPqbpgPZi4zfX+AzB3txXMLYmrBuqKiGaep4h9RFQAYlXKpk51gr4lSjY1yYwa0BkFpS3KVuCyMb
aChzSvX1x1NPuB2SVeIUhtiaYjo3lvDHrkxebUw10h2hv9rfEBOQFmBSWXOE8EYHV0ljQBh5ykDx
NVefanLiQKbXYuJGKnx72G5sTdXEpmXKWfU23tiNbIOE/e0AlcoVXNfoydQ6Dvl8ugbOi2/70hUv
DWBqsSvGCnQMIkkTOn5l0x+WURuroC864MIu3jgiwjONlH4SNDLq6f9i8zSXevciKvjh/OHlZEl6
3t/bIDTDt13KQfwzDSp2kEtT/k9AEQl93+eoQ2ItxyM6wjxIBy86EKQF2oPXbsXT5fpMkFIwqLY5
gubftOLI6l0JIAW5EEHHONOwrUpUEGi7HjhTlGGzyvGQwEDmvmrqrfjouI3Ds8KCuffLEQ9hBICH
Hqo9ZEOethF0MtnW8YGRU+JkE6DW6Gkh8xRLKJcpXaPMfSu43XfPwVMjS+S0/jt7RewOZm5EndXT
vBvp6Se/yz5kh8O6h3/x6+vaRr3QyKhW45JkJ27PnJc3oL74YwumhLY/R8NKKYAaeyu3XD63ebO5
H+l9f4qseV0/0BngcjrfbE4AEXcHSR9sK6DE4Coa3oPVE4S5bK+UY02VYpIcjLvDDWdCIyKtRkH4
H0lj7JVuLEZ7UCvurWrv1wSUYaRSo9WW3YlhuJlA7eA4yEKN1dOrVXq60u5X/bcSaTCws86MoiP1
4HN0MoIXDlk9tQjdcC5Xvii5zO6Ddmk4Ya/CLL6VYJ0IGLeqHBT4JGkwHJTTD7q81xCqt5UUjUsI
NOLpfePeCJuZUTjgxDUEhUdmNLgVPt0rnskzAhQWrkOS90jX9M4wzw4nqH4G2imRRnjVvYfFuKbW
MstVCQCpNWhGcWn/xXR+LuxQ239jl3M4+2p40BEVU/TQ9ij+ZL0adHJkI0ukTnen/ljHXznbZskx
fZ+8lZdNCYcs6gdYOuiM15d4EbizoeiqicUnu1qI4gRXUwGmkqEAhNv5QXTMdUvOip5hYz0pzi+B
ZfH3nviUJa64qN0N6cl0i5NqiS/Nl+jEBL62fzsKQvFIg9ylxYZNaeJqyDnW3eAwj4KjmHbb2gSW
csgmCaX2jmmDuZZM2n1ERieNH1kL8tfH2gC2BVIMKuW+zyWzvWsAn/yD2/xKxBYkmsTOHCWgnDkF
zyFQS381e7Ra2M0/Zd2VWXb5Ior9+ImrQwtqC9jx5lsxpoPve3StSODda+vKYs1vMz6bbqn+0+x7
R9X0IOujTyokl78wT4fCD3C7EtDrOcfrarN5n0UOaDVp3OMKbpW6Cegbsu8mRcGtk82B6OkNjtLS
VvK0bR1lCQ8ZSom/8OnSN7+RLilsOR4FU66b6giUJgeLQwqr5i5wWFDFhQudwYxHJ8oyBaUpse3d
eA/EWcHTiBh6WrVvQYENusU//fbPfGGoHletQ1lanKbvFmP4vSS7rQiaHAVZpLqyPyf7dCD80yQQ
ESklv3dAznidgALUcISC0dEowmgTbBbaq0VIEY/laBnOA2qIEhpeVUYOuO+FTaxeNaSVvbOti+yX
eyWdKe1qVIEnXxSyPWyyv/ow9gQpBcIqWptfSXX8sxtMkgW9RZiygvNpH8nirXIt3sEZekNsoty0
AGHpNdPC3MEcT2HbmvxMuu0YLJu+ylmzpvEFSrYKWkf8SVjmIIsqi7QtyMdkmZUlIyQdicsajUVO
3gKfUkaOYv+oY7ngst0cZdjbnkDZTta0DuCtPyud5EPjPfhgz3kM1m358b0OxgMWXyuM6zVZ0/Yy
JpbTOeGqIwybtdLXMs41+mespmhQV5UMq6ZEg+/DlE+wV5Lii0i1MjQIPvBKqYmQMM8fN7+QSdLB
zV3rsUPk9jWW4Mjo+yR/XociGTg4LKWHJZYXdQbaigunzXnxnWmvis4DY2eb8cxCZLNeRWeyuUcQ
v2bk0TWapoFKGNDkObIwTfmCao9GUYClPKGSBPja94WuPjJvRFBDp3I6U+EXQOJkzby1R1+lKzUz
M2E4JyNoJr+Ba4yGk4meLWcy0pXaXe70t0ozEHJQXAoFa2LH6bGw9VHE/YJpsV7nKRe1RKPIGq9L
DDAkZBLGV4pu7v91yw7XGgTtdGP/WEoWQW7KzraJATvqerrO0bannOZfEvx3QySAjGHsFEbeUvKo
y5Iny8Q25Q3055k6uWK3/9NCS5Dy7x+2ZTDOM2XQKAUUlvcSMrtCyNmvubTKRAsaPiRo6PQJlglq
+94houX+rpNhY8TZH2ebaZAea8OQLB7zW/iPek/Og2FrOyqd7if0TdzBpaYRJwhQn1Bjq3jtc/pX
UgWes1D7trxOUySRcnP6rC03v2dPLBN0Z3r7SLxxsOZr4VU+60+SXWGCD0xujdG+vWrgKY368Pn0
sC7zsjTYKIMnX4rVESd4vtyYqkd/HE7lSBsxSUlZpKlCGb1ClZTQFPQK58ItV74y4o8ZPNu7ltRr
vwoh00ZLrLgEW5rlSqMXqOraoGDo6DJhyLf5O/NqY2MSNFLr2Ng6ydtpcdlbLUMELYDaxNdfnRzU
snXgke9uZy7kN/zsdXgh4YQjuSskpC4/vHt2u6oQ6O4XVqScTgIwZK6whHyi06eY5osKho/kGAw/
FciDFaFJ+M9Rgj0hg4CaPnFtAcKHi07UvWu8cxJDVe6teEPhaqeH4vTKIS0G7ncoGawld0csiL4J
NinfoDPC6rsZL83jAHtdgOPXJUsG7MRk1SdyUXQSZ+2QaRAOQYertNGwYbCsuc3jEgUAgE751owZ
RydaXC57alMZ34V7ML0NK2bo5+Ev7IxcLhtqoUFkpxx3GHOAZSmQqzHrVjSMdu8KtDhVMuRoyUsN
vIyC2wULI1H+8CVr9DgqzjJErDSirdoBbc+qVClW9huqexlNdEDfLAxxu5hH1JOgUZRsvqX2mB28
6WCAS5VhYjpJSBTKhNQXqn9h8bUaHtSNHIFQAx/T4+4cO1dqs/S/NPyOF0XAerbjDi6YrO8TlWMJ
yG0qQ+4Ekt4HeDJzV/bL6cLNz7TIvlhENMVbb13HSz+UwVgxbMcO/y7fDzKBKs8z05mBW+34rqzX
2+Dvo1SsZ0P695JSXLcPqsD34z8tME8WTgkzlVjbvVVCPp6b9Xrj6Nn44KxMA/RRRBAyNuh06rAS
pKq5hX4cYNFe5fq0gzgnzllF25acexL8CDMqaxMbporPjk73ZNJ/xgQJ0KtmfHkoXxax1NAwEprE
Vwu+Mi/cnawJ4LBMCfSwIl4GNxG4QVzxE9gzQBUK/b23l5jS3iIiaaIxFUgB7FG9H47NQvFDrUb8
HsJaz8jUTGfZyk3m2gDF4b6cZKb7b2nt9TGms2G7979Y5OgVrUO+j7M264NrfjBzB3CDxs8+lufA
8d/I/xW5Ddon459pK9uZ5EwlP1lXI5Bd+VJoqLF7f49coJGMts0lj3T94FZmvexZhWAo/U/N3pkb
V5DEGE44CQywefovmyQKaJpIgwlomMAcGvz/EIpuO28ON8aGLFuw+KJuqj0gna1y0+TK9NzncRil
wQwPjiKTj1iKFcOctUVkXsPC6QfNNjXh8AgnV3AvEMMC017CEriGztGf7B38hTCE5/9CKzi6swiK
BgKJynsPlPbWEeDXgyeONAEyHoI4pC4L152/kLn5d7s1vPeaHc5io9HF683+P3sooKw2f0PgdrXQ
6v5CvVXrpgiuhJhSTEAe7HXGfxcTkOEdU3aZLc5CQh5AbvuNxFA1eQF7OAdoPdV5kwTS14WK1Px9
aenHOJOttoWXbFNcwe57jSqkcLu16oEQAqMT70D6uiRXYA4PAiz9ZUpERsWkoB9IVKAG96BMTFzt
LwDybmVoJVP9hHbqKL4ne1QJi7GlPfkMLxKfXWcvr56msmZ6i1B+SgJQ+vAFqamMLHBcfFWpXMNg
YSQqCpXFMc0SfEI6lxdRfP7qbIqCsih29bfOoijI4tH2z1D8eCfQOOzdxGIJy0cMWhwaLWseIVL1
egBpfxcButbNEZmgOoTHhK/jvWgP/K+gMcEtr1cpXfQkDvqugL9KJHjRgAJ+IMy9EyW5fEPT2CJ5
JI2MRZMDEOjBfw1qCnc1wxkXFKR2Gne/fHCGeWJAVSTI7WXm/hNGNO8R39H3Ra4S969DsqV96/l2
nLBInm9OaLCf3Uw/0+cFnsFgUHIzYC2ZpbiO920spuqe5u6Bs2UUejx2gNdr6xdiDy1WFug3tvaa
1jbSnYzVQfTk0YGaBWzKhIlZhuH1eH9jI6dSu5SyB++7fO9BVCrB6ayHF79x8SfwyLy86cOUu2Cl
ZZlyXO1HNb3khPBnSbyuZXd/jiiV113EgZOlcs4ikJaDBiDoQKsGxBfu/TFMR9cQ2q0bAqSYy96E
2xgMi3Cqgw/oUVWOeb42sfXJH+sNWzhYCvAqAl71zqCPf2pUP3kONFqZaiuToQKgeVgCpsWyjnnS
OmrcrTGXJYwVMoEhic1e1BNWMuB7aI+gVCxsX1OPT46MgHIWZ5SyygKb0ulQadz1GdK3cz+r+axP
O06aUAzis9kfI7LKNKTs4fs/vHd86tezfsnSMywgKFsMsHhV3kGwuvU49w2m0NYTaSUeZLpTjg2N
/6YkqIg1WP+0nZ4NU3pyc8xmOZ7DSDCP3qE08TdMh/EWfsMMFadmLXvTyNVx136A+IiIUGfeEomd
jOGeeIMZdvFU6vVxHVUEzgDgSfEsy+Ns0vtptCh/48JGfbRUroDUNVtLzMrBnV7xm6Oo1iaymHEG
jPAI7tYLGpDdla1omq9CycptpjNi2R10o+C6WMMsIf65GdNk0yEfcI/sUXSwWdSEknSK1ekYL2S8
SMwgDedEiph2Ude3Wq83tW+DVuTj3Cshu3FUDSeWlrHCReDrCTYmjAPfFXW5ED3MrmRIiKmrAvU0
+dLMyCkzvKglIRZlCDNR2Et6KKLIShz9vkD760hu2fZw4qoQzNnrvBkf6Wb/Aokb7aWQ56EPYr0R
MTrLrMNlYJtvpng5oZzhTYFujeFobMOwwH3/Cnyh3MOzylopAYv9KjegM2qYbv6+ekttObNtoLLk
gqIlJCu2/EGZjzH+/trqbs4pQP6NuNSwta79KZiNMlPV+s0ybg3iTZ+puCwIS1SEKwA6auqe4Hp+
BPMENFZmQglnq1UQuBy21UhBpKsjiMLCsfcTDJpEtXXBFERmnuD05W94CzCkzICnJ4zDp8gr8DNL
kUvgdiLdvAtjheESwC9h5v7ie85kgGGdLaxE5hcGkj0GkvaPoSswh8v1Fq/HwOZ2nhwLpMtQk1Ra
cfyQ6X6LPqNMGp+SBdtCGHz/4yAFDiUXjegQVZaNCb6MbOs9J5vsPXiSOhZ+xyIWH9FWpYH/k9o3
iEcRBLyW9kvmGc81wS4qFyIkglv6Kaa5o0oy12zQJPBuOqFHbUTr7NIr5vuyq7ZlAokwSv0jSlau
jg2l4I18dnQldUuuZMHasIx2V0RDX0KuI3IuqzVHKhaN+LIx3nsrweuSSC6GIBINtL7F0yqZm5dQ
rAQP1wdCd0w0Jz58QFRm2Ptwl7oE2rl8gI0AQhPx9gBCz13DJrTaKRicP/miDlARgvoLYRSlVKpg
Ezac49Q5J/KhbniJXBHlrWULTnN5bNIXaZoecm5gSvUitJsKO4RO6rHsoJj3JiF07Wge7sGtIYSX
Z9UOvinLjEiTETsDCTXGKPF5u6gxDxBx7elyy8+cATdu+gC3mHxhEWqJRqw+fcbxk5jaXzBs3pGt
y+hdo1Q6ZNoG9agN7k3xDV6bFj1btGaKPpRfx9uGYjiAl79Tn7fVPPAaaI+47afx4askyJRWafVD
StsC0qoPDVYE9ZVUkBdwEAJLkJ8ZhlXrMcYGmUVOK5pGkHFx6Ilv5rH98OHWb/tJjeC0UjrGG//N
mK6OOeI17ZRDT1HkTjWCSYTN0avJ+MeRoVBXKi6Tkg95Ri6knXBnq1/IzpiTCFTjPOE53ACz2Yyk
nHc0qreCvEJxBGELHKEaFIUBorW3CX+USaypcqqto/lDPfNqUmSGDNPTzhqK0BU+mrWTn5NGgGKf
etPDD2EfbYkU+QABZGYLQwDzuWAaEWf7lDWrlK3HfU8GB0OZ3S7ZGKQCdrAI29b99ZU8dctpkwAt
9AmQ7fIC6UK65ws1NJIT1kA6xJ2Qext1WOo+ApouIC3lCPPBaMsWUAZQaALK265jfXxYEh0rM4fi
YaXn+1G4cQhNxeKh7mSuKajAVrBywA/PmhxWwTvA39xEbh0abM09Dm+Np82Botlu+JWFDalPeUWE
BqCG2uFbJcGZH+bHoHBendRh51uCO7QJQ5PNa9IgeFE3ADeZwXhARbNBwgX0clbw4Y4NG1VclGF/
cLrmXyjskCDLFdTGRIiPyQZqVEypc9h6SltiNIko8DQRftBEzx5S7aFzuSXFoYRZFANiPAMLTBvA
uXSgHqnMMDUH1r7D3mCQfobouob9mGmqsRtCYnw9vM9kD0UKUsSBoJnSjGMcbs8sHSkDfe9xGaak
o127Oqf1WUnv9R7KmN2Zxra6HuXyYqtfXEta58+xjrbrIkavpY1Ut24pqQIn9VJnPMTNF/6WobMi
65ssJuas2pbvBnLF08KAksZA8QeJJXqq/zmRZ1xctuYSIfO2FqOY9j2M7QgArExhX2K1QpM5OHiz
UKX9bVCUmnw1jxy7LlDJ0LyuFqQ4qKaSUs2CZ4qm/eNYHVQxUDdV4k0e6B308jiXjma1usu6eV+2
5dY0iiwchd+sYRFoSNU57ZaRaB/xO24UnGP60mdMUP1FlCSGg9S0IbX9T4aIxVDyFnNRwSOx8a++
OyyTH3fqoG6aX9aDidZRPvcYKvdNCqPIf8ucCP9lIGnlNSrgYDCjAUd11DbZc7Fskx1iXUrTePrJ
f1wLVYYNP6qbbsHr9x75ZhL+zzDip20vS30/F8iU+S7n/QOFnnUJemfX7OvBaLbfeQzcghlpZVJ6
3llutSVQDWq3riimqsVx/rM3olCQ+5Lp8RO53OHqqWRJex2ZQ8dPrVaw1em9vURffJg4PPCOpqt8
xWkm+i7sc8M3yahjL/xco9hUIjTE56budRLIrMyR7jFlogTs4UAggR6Zvlx5vq2OsRRa/e9lcHtL
h8v51bbXsVBS8md5qwd0C4tBHdLlVIG7gEIqwwV0gHljc4HeJgwEB4EUr5p51bGbDGFWPTyB3rEJ
WzWc6V7d2JtBqlLyi3AXhLffyo22vyUiCq8jg1R9msZM1jrblS5V75VCIAk2Kvf9onLCrswTz9/I
50Y7K2q7tESh/Imd4BqYJnz3hNUhucZMu2mwKomHjHabJyYCQT6q3HKmqverFTSI0SyBH4nzTqwG
MbbKaIexuXOhzjQTl4iddqJ3MkGjSjdZ5zEK6b+z/MIQQah+SKxmYj1dOFvq8FVWdpBtnJKmqpg7
qJ3FemlTOXlbrgDavNMnEe48Nt4h+VW+VBwVk6uxCCA7k/Gb1BfhVHUsy5XYTGbiLsq3i28d0uF/
O1gXtkPyL3OIz6Yo4s6JgYnCz9M36MgdA9FGe7yVL0xtRosKrSOOnde5P1FKTQpZxGdHoDaTlInk
hHWnu/2kawhdJ75vlV/s4EEpf/vgfQgS5jiItbts/x2b/g9UcSucS2JNhbYc0dsgnBcUOTqElq3P
Rd7aJGvnocsvbNwd5hiwupjNl6oNLD51bdHcvwT3NGVhTizok/O9Gn0Y5tpVqncQeeKu5E6xIj+w
rZhW/tckwRybasa77O5kd278UhlqR03bTkwWOxOtjb3xYKaLF3vuZTXXROTdbWPZS/mSRnkpKBDs
JJD3IixN6WtBYl+D+6IBNddrvEfDRtm3996QQjtUVneS4mf8s/RkhhTlNB9S71JF7E3pBUpzipkz
EEwgS/Kqd2foFNMYpcDe4vj/k7iitRt0EY3R7hfuacxzxRZvKck8pj+llgd77jXQ/UEljDGPtfH5
u8OzRiCNaO+X4eVtpqKJWUq+symbPEX3TX2oFlmHZJNK06DW0QrxZ/GEZW4iQwA66ybQzVP4f6TM
NtJKrtJ9iDF/ELe7YTbjCW0QkoK3YFahViWJ084p0MvY1V+5H/y6MYDcb2eDudWb/RbJXoBug5EI
dGR/mzYqfGPoJhCCaZdXxHyDyXVOqkG3UlFjcgQuGbByWcFlcQxjNjZEBqkuoUjBgjstRQmoyqOe
e0J8pptDeOAjgoLbbSD7qfvqdSN2LH0QgiLVNNu+wslmUh7+YXc85monNmi4/bvJ+lIKX5YkqTk1
9TgrVjqRU/OTcrnxdWsvbdKUMkOCTqgUk5N5PYpNU6hGM2SEasKME1648audgC3Vdb22XdmmGIGB
1Ee+CCLkbdF3yrqCd/U9eozmNgSHwCQquZFKsmx1ezxGZtr5nStjMvHVWRGKxtelB55sxqSAGOH9
vPPeb62gHI3dP2AgiMvG39keBSZMrrMJUtwfxCQx74SfA7TjM2uhzA/DSc3eOSubhFMHgLOPBWMD
b+XKqg6HZWOr80XL1MLTFXwIfjzqZgLZ9ymlFEpMv+c82HwZ56kEG9HbjnFw2/X33A14Wu4i5F59
fyzMFsQQN8CviJTv4gSljGKmLfyZXk7p3044FRSJN+VDTKLnrmDGf1uV9djddttk5Mn0ydo6eQLa
x3s6zkRJSvlAh5Fb5KNanKNZpHgturgnc8ZDnLVA0quu3E1011Lh6jzR+HA7530RYhzHS7SGsa9Z
MKa3qWQ2gCvolwlN0viZctIoTkLBwe4XkhqbQYm9xq6ipH7PahtJ/4/QOIM1bvEE1/8WHGNWbx0S
D36QNa4QRTymYr/T1c5VdHwP3W85HMhoPEQ0VAB1jLPXC7S0hqn7Hw2Aicq+Jxh/aSg4t+FeQgoh
hZK+XM6zzXgeRpK3w02sZ/9emfGBqYXNSqYfwoZJhN6LRwpeXvaPSGjzycooBYYpkoa9jHHXQWgg
1duCHCvziScla923Zcip6q18Yf3cYMWBcNtTMd/a2FC5S0iJhFnrFa/Wk2HrTnmtdmZCTuKYXZ1M
OHpbZUDdmtkbvPP47juTzSPtCsKrkEeaB4tn9z0OzRkGTuJbEV0sigBxUaYundJpTLvsmrHlIRVu
APLKt7TueH1HrpzE7r4MOTah+LzT+XGTDalZpxUL73BxcxART5rn0uGXHkn+nzi7G4RXgjKbSHzh
gkWDMvAwozHfSiIXtzpFbsDV6aE+P8M2fcn12KcnrImhsCT1mcPPhQJIYJQELUpfQXkELk9P+aAo
wt4U0nBPOCzj/6uqZSum3gqF9va5/64iSW277LnbN3cZedRYq6NEzH/lTd0AdLUioJvxtCFsv4c9
luS59wyUd+s1MNGsgOryzoTn7wCMPMmEmMs3YsAAcLOHREcbNmDm/dpFFzVddb1PWBeJoKtgLKX0
eZtxsVdMh/6L/HQmikQv0OVQboQRWxICD2IDqI1+uwiaNMW7o0MIOQyni9vsku4i9gQgX8AgpDT6
97TXMDDafxKdjnG6Lg2JBianOLImm//SGxCYFDM8b8DD7X+l2jWBOJVFqaivRzDV+ZlUrC2SzUG3
bsZynaweNzowsqWIeCNyzyjHDy68gLGTy4w5zF1Vjn6mIbkLCQ1nzMo8cMUHwONwyw3D96sg3S+M
opB/n2BOBND9AFLYYoLemf3A3GRDaYwXrUC7VAlqC8NfRIMox/dBCMJ7xEfglkgSGKemJCMu3fm/
7rfApqtquqDt+0FF+fNSf0P4TaOS3by+QCoPTF9Xewi4ivpO4Tc1cwArhfcSRYzMU+lzMaJs5LS5
D8CoClRHpnyMTo2S8zTN0UHi5PhwpMZ/INsjij/VVoUZmNDMsE/pFTu+xt/exTKLW39c0WKaDVxy
+Xq+WUh/QCpjH+0GqMoUYxGpww8xBEyu6c+AjGwb1ft+TblHZVY5aBybPYu+4e55nHBWkufvcRH4
r+sRQ2knTRHet89xAwSLIhofWdj55w9E3X1vsO1lG+y9nxcq75Jn3TZhzHnbKvHeAbvSnm8JPi8H
YG4zBvNeMPGHckPUSVSYMp45G5hAGYiiU+ms89MU6m8l2gBrmILe5fktzE868MHR1l1yjeIjUI6n
jzDUeEdK9EoJ+0GhvFkXGWZlBYbHBTDhym4/pXJ2TvAEFS9l2l9QL4Q7Ln3BzQAQJNPPMaxU3KMq
R3QRu7HGE9iri9nttj8zUs53nIE8icJ7KIJByYgcSloYr0Pw2CXEhrAxOvf6uwg1dzAO2dYFACzr
heT03MG2W4L2YwLB5KCbZz/yHRxSJGVMHw1UPElKfjFUsvs7HqW2h2QrvhurJaycLzBEYvGieskd
QejZpHFs4Snjq9J7LBNGzVlUzTEMvy+Id64qNgn6rfKhGt/IDBGJSiMivyKaGuLOqGYTZ+D+pLPz
qqNbnMUGVY4RP8yIpF9kKEgcdLRuqZyTszxPXTuV0HpUBGK8Vn2icjhRxjsSwvWSvJVZamXCVuPo
gXzjch9mzOH36quX1KIo8QytqA5c1lLEhzTqa+2I/2fd+Z/kZ7wSBVtRGyN5sBdwdD4m/hu+9poE
bA/UpuhUW0Vn+MkEgX4zvLOJl5hZ5MPCNhH7Ijs/lw6EsN5XKy/Y1VDa7aOtZ3hzgt26dNCp3QEp
/z4SwX9qTYdllbXWzLhWc3jssLJL+zo28R/o6wfVWpBHm1jKj1Oh/jqBFAXyM8TyQJpaHZx951ZD
Gg3cYsB8DsJS92pOwH0KJu1ELbyZO3n5kkA9tMeEM2sx18InZKDJ5tJNwrznlRs5bbOURsUxEb36
FJgQM4RX+zYCYWi6NYSZ+s9fhb5yNS07A/IG1PoHJBY8ClCDXjFtJ5rSdWbOHsngQIvhLWLe8xR4
M7S0gqBJbB0lkDUMulEe25NodOvdzFjswqEYnRwkIbnogf+OKPeMJBRGyJYFLRhtfDLB3ipRPLjv
ksf7kBavXlHOITS7Hs9ogoXKJcxxqezHkMsS1cHFyMHcDhD1luCYN4UYxmkMEQiluCwr3GEpGmqt
txjKIhl+9x2GXO/HZvp8DG+0WvkMGTiWA24FQhFOEceWsvurimqLIi6r2NkQ7kQbt8oWXU5kF584
/CxugGHUq6o8w/Awe6YPbq5btTApyTX9DKK+uaR25mfTN3RqPzYzzJocf2p0GlllF3Cy9MVQVliN
/zlSfk31Dvo6g73dRlCKdIEORBOPUsQXjq1XlkLs2wZk1bJLW40z5Kf3Y0g4mYuYL+D6SDtBpPqQ
BFrA3wTqGM03w8EcjGcJ+W7kfVr0+mpEgEEc7lNIL7VpjFZdI6kkpDXAe16ZYM8eDLhtrKA8Fd42
sPqDIX8eW3RI1UV0/znkM6xrHjbdRuOoujUZqM0pZZfgYKk4PCEQKhCItZiDfWk/kfUFUMHFgWX1
GDcW5J63IKs0HLtPpVlWe5Q7QWQyr4dGsznFD58vWExCnxXXMstdDmWuegecgra8Lich+DulK6cx
HmYIMtzpivZPS3A3+MxH6h5S2G47tcbIWnsGNHiIH9ZxZTK4OdYq/a61hMucldxAFFgMT0Lf1oHZ
QTxqu4pb0baY5eyARWu6vip1WBbVG70iJIFS1KDL6EWzTa67+EoWd6YhQ7E6VYe7CeAn7h9b9dBW
jlDwJcTui1f8V9XYtDs+WPl+somGG7lEpPCMbHzuLwZXO+Tgt/BYwOB4pmz/WJaB4Ddvrbt5yWrZ
44w3UnsXqIi14W96jw8KdxXFM9gd4oZFCFQ3DFunb5BaUO9ma3vqiyehe69C0CDbpasqJ4fXeGoJ
1MI6HDKy/gdadoluKBMbxbzAs9ln2av3HtPispChz4pR1il62LtssquKCi7dRaLYiUuGNfH42bJZ
T8wx+Y7D4mwMPkBdQOQIHczsqV3jZ+A/ZnO1Yj9Oh01iIAs0ZPZrG+PClbLDM5rWvvHbtKb0Iovd
BGzh2FFzC5KjTspO2UqDAp5R8zRHempGnni0ycFnKjFxkiFU5rDndVU/CgGWI2RCa148XMe1P6WI
4HLhQHP0xu9rxPSHuJoWQg4Av2LhHrM1m9jz+ifwN/xHwmwcTYu2W39EmpYHvLeKImFszbAziZdO
B1yvryEfyZUPICaRh8BNjSGxYWKwleHO9enKF177btcUvV2vjMVruRuXsVyJa06J/2jrbdFCdr+s
FWX2/7532sNw9C9nJvcFWZdtQvatj7/ieCNH9z4kEjEjGX3vUGFooXMUEyaquPf9KV3wLQqSjkTn
jRqvTDQEafswrckiA3MRFFmG0VMGhVXp9t6SpB0f0FXppUblTLZAk/x6V7nB9g/IOvLqdFlZH++L
nyyJguS/u61ftKhss+vuP+6qW0WEIsIrBaaEDSgirF0ypH3mwJ6q9gjx9Bevc2WSGigmXB064KXR
zG/jZdFqP3mJIfNNSm3TQ7NUkPgRzZ3GE4nyVIbOMpyMEfRYL1t0hxec6jxIPLD16IdLlbuTih9S
fPEVOD99x2HcxxMrqgO9NjCJc09/TeauyFXdhIPelA34UxzT2YUylyM2wswa28KYkMHNnVm2WrbG
PcviNHjhysiwuqGw8hRvQKmCj1iLmsJ/jJOxDVdzrpifLi/me0cZauk8Zwua/gPmQuhbSwiYCLqO
bSqaLHNI0w3oIN1k01NZXbu2CL3hVH2zNIDGkvid1ANE1G4LWKnRVM1qJcYIiqVYhVt8sbxSuq9W
UM0z2jQeAdffW+xTXyXXFgHKg3apZ+WGQt0Tv62RaQBGz8k7qfVBZH0zCF9Hq80dOBPX6OzdAKNe
YqJFLSalz1ifJOch8/BbnwrgFZqpDLQglUALWwdiE9qG1A0n6xxqQDbILdUiPcPjZQ90+oLVZazd
b0Zr3IN8k3RfZ9D6BTY6AINsOx6ZBZAIZgdksp8iJQeuTAy14padrf6HEsNusHdMdVZOtQOTmEml
nIv33/HInhgc0/bhNazMwTKmEkhgzwZ2hA2F2tMDi6b7o730+Jt08Ca4suI8vp+At0HDHZTSob47
WiiXckZQyq0ahjZ8JwMrz5tjXrOl4YCLOOjqyP6UvU40be3H4E4uMDy/J+NNXTqjPLI40QALJBni
n33Lx7jWICJrJ4Wu/qO4ZdxhsgJr7CG1zJGopkqGgCT9cP8Ygz4CJGU43X9fCs6ccfwCl6Fp8Ahr
5NlKRWkmnk+axl7svrn8Joh0VHkZnk5KSY2fGatIvbfwLljsegPXDg4wQBRrwvBy8HGQQaFxARDO
V/5IaQ+0cjUpXl8WePrH0EQ+JSLGMpNlwDQN1N49LOv5WCr+yylUl5ujEcD6AUvLB1bs2FwePPAl
hw++fzFYYj/ryUZaq/2jRYzboMuZ2m2oMNURNIBWQs3dp7Fh94yuC7TTiLnyysKIGQUKnziQqhqZ
VSPfV98BgxlV843A+hWjGeVRyA/njff13y//sITNzMVgy4kUgfUmHyvk32mXMDBV4f5ZiGVpkCvV
qJhECroNjaPEHI786tLzYf7VFtcQVMOgeK9ovkr5OvPbhVdvei/4E0K+2TaW1pIMRmrkmvponTp8
Y1TtNeRI0jI9Ni/7qTpKpd3UOTfkVQ88YBiEaKfvms7B3bgTcZiEC1RxmjdPNCr7vDfsoJfyErgy
HVQUiEcbQ4od0NEUmL3+Y3r17G0Uf2qFfQnWYwLcTpXqANRYJG9rrqN5epUgSqIprbJutC1MbQB+
Bc0ZqXCiXqxqZWP5KRGlOma/VB2I+dlEOgIMKKnLwUlrh6iZWMgRThbjnGaRm/31o8zfIEyLQqrs
lQl0P5shPiLUGwi2BZ7pMpmjfqpunGzOXP4bwGf6Qcvqeqyii7DVdZ2pi/Q4n09J1GcIagff0ZNX
+pC8EY9bq5v5pGFtnxxLFLD/ckbuZidXiEzsFx4/0FDxz4YA9MX6akrvN52zx/XTmNpZ45k/qg+1
t91RBGZvx7uHfeF3OeQ0i+SSoBEd4WgXKIvkU4KgDX3koFfqmJSUi1yPRcyaAQ/SFWe/A1NroZ3e
lYq1BqzIANgXjPJM/3tvI3TIJHKqAYIFLZMoD+/Hco/Lm4u02wwZZP/w9kbUg9RcPh5hhiShc1vC
iQviZmljfuOnSiY5+C4EzEvMwCfNW19lO00Cr0QgHqMoFhS9vI0P6NIWG1zlC4kRTj6Z5w+HSQXT
qg1ZMpLHX1iAG0OfH/ohWLpb7iXk2aAJZ9SrCKr7OLzwdo9luNmx/qxogEtnx5qylCiHvsu62RjR
CtLiDzny+Y5ZvAUqvnMONXt+rnkBY9YWyIkmHJhkdd6brjR5lpB7Nkr3xTIv4QbjZabrpTrHwmtt
PF05teQMM3DqMPyYyTH4Vwaj30+hMxyNN9J99Krqs7czBqA+YcpQ+1g3JN3v4efTpOJ41elXpU9J
v4zoQOkaG5nmA9iXD8sTYx8GG4sGxzNFUtUTVKOth4IfTXo0rxTLxCApdDP7nxH4YeUVNUzyVGCk
LF5HARShVHzczUPEwMut2S7LdPsRSyyvDYf7GDmNu99vWw6uKNdInyUQklUh2nlkWOdFO8pGHkdE
N9bxufNdtmnR1Gc4JNPBf36VVfo2FLSEeIeTEZ1FneMRkfXzdPjRFUR98e6fJ01xZ3NQWCu9Gf7L
j34vnYY++w9154SXetsBarVOIoHh/u3NArZJMUxTMRLArJ3DWT/Ae5PgYetbr0Pebpy+qFToEEUs
xu75v+7aHcsMTPFyStu5pIgADYYr/RZnZJzU2EZBrDKVWiRl5gIDggXoVBcUVeUvppBijojQO3lC
h1C7wTh9niNMuFVmXk3Mi/BiO62eg/1BEeuluDs90tbonKVULTvc+5NFX6Lbdks3g83bptctWqoU
HFiqE6H2BoL1odDx/fjXcmKd4W1jqu5Ebp2fx4oQcPJSSuC8X+DeuIb3SpEb9sv+8/eA0eToyGtS
hJIaW0wRULPaWmWZWsZrmQp9BXj2wMR+Bx91EekSUc7NO+1mGAYR0M0NPJSMvvQHcwjaCp1DZA1c
3sXNN8frP7iGEnr+3MyYsUsmYE21Md0OK1o908P0+e/crw+14YxbDFjHp8Dpn15uuEtk6H5zK1pJ
Nsj4u4SFkiwRF2+99dp8+fkTFj98PdrIbV+jUd8Jtd+jnFtesD3iqw6UGKXx9PuIRhZq6dQoQ90c
AmAVgphgVdqGO64i3BYTKWNs1T0yE0O24W/TG86oAYDhO+2AVNldH2YK1Ay4AWHDxW3cevwO+1MH
XNWNh9GBZAXd4SLRkvNookqY9rQjSUrle1QomahP2+ndUzeXYjmJ9TyaOUE1HOX98Twj+tT95W8G
b/7HC/ieqihfY3p64tQQp4kMThCpk/V3CM/avZmowLPRDDl3su0Z34UqAhNq0F1PNIcP2qnG75Jn
3vhjWkEtPDuAMKWAT1XRKW4LW5UPvIUk7tGiyr2CxbWNDdgpoxG6sfOUepaajleCPRdxOvhdI8Fo
BqdbHKNRfZ7ehCRtfFOCDRpj+HQ665gRPOhysoZ8CDgrLebQM24t9/GXJl17wBIndFJuh0j1EfBW
GTonk2rBHmAZ5ZpPPFt7eDHDOv8xiWXUojWKMHO61CPRgGQ2yCsc3GhpzFkevopjoW7QZclGmJ9p
pRn5M73TiUMUCgf3vGYBXqvbsZZ+yP8UMV1SlSFjHzt03Rgf/MJR/Bnm51r94bmJOJXIC1G7BCPi
mrtoUw8tm+ifbL/tF42LJUS5k1HzEn6V0/RKWZIgVgioyp69DNUlwdorsyxCqs4svMgmpCfsfMoK
gHMaVDL4WrnZilFrZ1BEA+RYdN0cQEonski8DYtDUiFGQ+9WBuKOjZsrJ80G4miVcomoA9hq1Zp/
5kEcWyYzHfFvSqmq8xNtPjqahs+yV1N+v+IdYncHUH9yaSZw4r4jqXQd0AhWSklhsOPCyTNMAl/w
3WrmbMjq4wnNEvFdxkXRvwk4U+cIOSLpk42R7XZ9YeeIyQTfadoHop5eNE13rCGjKGhZ6nJUpiDE
pyC3i6AnNhkZDoTlwWnNpmLNZ4mEIqTr/yBIxneDtWWhe4LEiei9c7ud220GATsm9F0mg536lnpg
tIqYOMAL6WxYRz6YspbJREZaqHaTi1noIxZPRRttapPqQtb9jPEwbFI4ZU3pKlG7QFvyRAC3Qc4N
OLmyRu1Filh2B87JpFujH9pZV13bHHmX5gpIVhdB11N9o+xpS15i8GtW5S6EUs3rs6z+tBggd903
Bgmm+zqv60Sm1Lc5dPv+0RXViAboAB3STKmvfm5ZGbr/3wbLLfPR6kjFFN13cqT0pAyhpRcrGQ4E
fBYMp049b6v85o5iy88pU55qtntByirUB2o37sdNdZBKs9cEqGiHBT10Mbpa1zXLj1J9e9T6mBc/
zt4DJgq5k5oR2qfmOhfawv+RieRM2Ufnu5EMdtSYvS7cZJV5qO4IbrYK9Hv6lVqrgT7pWF2vu3C7
I9Bi6SvMqsJ9Sdk8F5KTuUvmsYIlCLNB0DZqhZ8eWBAx2v7SdXViqUQvh+6jw7ApFok5wADroi2x
RN4Dc+mXP4uxelZM7wHyzhAcJ9sCTGbWC7+Z3z0cZyWN+gIRfuzAZK6Y1QEpHZMdwS+5WJ80Oivi
jHI5kskhTomj+foWHMws9HpN06YnhRaKZ+4guliMPM3RetZUXWEtkiKHoRiRnOnx4pnzEIhGbOVs
xwlV+9HJoKn9+VGWpNYq2DELXvUF8794/q7Rl1lrWWlziknuz75wUmKTj8hpGIdodphno8spftba
Yt713nq0TKt5fshrtfz7WLnX/LXHP1eYmW5jzMp0EgvR1mjpEQx1k4vUf6XmSe0LKPP3zppXljNP
Z/EMMAfbTIqR6qQHuDrOTwTrhuQP+S8nMYxuTEolT27cUqncBjw7A56mXnJSjm4aZpzdrBFBLMrs
0lNnkTIXq66OnVZFhxmJxqYtYK9b6F3bjGVz0aeAC5gjv6piQKMSSfDHKkQTLb4z6sKFwZpNsiPk
ecHitRHdIVxQrzZPcjJvvxM0BWjiYWAl6vAfiZkDzEhWdCVQrisnCJB8UXF5VITXcOnhpzJEQA7j
GzY1W4nRhz7Ykzhkd3XxAkB6jM1lzXzIgjQul1y4fet2UbHdG0Fe52H5EoOVR18KgBTZGWZSH4te
9pU3pXqCBwJ6wpuGVai6lRXyi6rw6ZwgezmGqnjza6MqSEadgPevRtbaqlxVkDJ1lJaOAYbdfZ6k
aXZp5cU7Wrgp9Au+MhTDTp5jvtmjou9JaMz15y5b/LkPmyW/YV8Y1juaeFOkDi9xm37JEcFRZSSR
73YvyYriQVsVtDOIFKz4jLVhGDsecNDePRzVV81iwTPALflUm/tCcYY8NyxHBi+bkrt6p1PrY52P
x9RBlCIFPTQpq5P0vNkuipJ5ALcex0kdU2KQT9UDDImhiNGjLHeONMMNvTNabc2Z/Vd1LiFf9pI6
/bCaoeVN9Wfo6p98N9aaXCOy5PF2SH8YY4GwwIQQ6poKag1dsw13YC4T/s5DCcmAH9BGCesreVkI
km1q5xrHBZLnJdeRr+4HOKVxhmS2ubp9qMPYzdnMEzCg77X+bXELx5K4txDVUK8bOeFr8y2YuuvR
HfUIemmnCMS+UXh4LCOUgQPKgrorE5QxDKT2Xm0cA5X80YA/WFu6bdjEEvYr4SMQhKCCM4G/DBhc
+UrTvnKYf9OlpOp0e26JuF3BuXwUDu8lTNREY1dS6fuFl+BXeJwQ2Fwe3QiK80eYGZDx0EyxOZhq
y2QZP2YRvGoJrPl+stq2BGC8GisvJ1/cZZeDVQw+cySBRA6sZXokMeqejmNwceq+mMUXxg2UvTcR
TjBeexdIu7RJZV1JgiGBYCiUA3+dM4SHCToauyPaqWJSLCuB4OuxUyz2FBS0QuS2VyYaQfX5qiUV
GImsMwO+W2WHYLzUbkzIVd5qicTojc064uXaIVUsSRh14JY6KdJqQxThbde/BXQaEhOFx7wIZwlh
pMngGKECaekPjiPChMbAvIRTH9jIg3TLi3nJV6pyy22Xwh1QgEmKcfh2QXwyYGOkMf/PJwRH6LAe
KsDaEImTb/U41JMVs0OrF6OOHY665Td5gADrPRnvPTZB4Q+9Pk8dubpP/5hCjZ9CmUzkhinup35/
Mh/PXnVp8/9+uNUn1L7e5r7Av+bCBAZ/Egl3DvELBp6xoMsromuaYZGzr+ZxFlftd0/MVeMvqnxn
DK+Z7+D/ubAJFi3SHgxap8+hSsCDHvZifgGIg+K1F6Ahx+WtV4xOETwuJgblZWad0q2KidEbyS5x
hcMIPCYBJlMSf6JZcVqt/uxwFmtiWH42akac9cap5QL5YGV/N2rsbP+IHzvpJNbVk8H6cMlmjrlj
HcTtEZjPfYRKRIJj+PZsmelK3JdcIVDr57VwKL0gJnA5wxqL6kFWilUhDgyKaZK5twyleS8s/wb4
Qx5I+HvEhr8t+o7a+W2i+n0aZSpYjLnqQ6dQ1CCeW7pvnIko82qsEi+WcNtaBtgpRo/fLgYnnKFP
y/85UrUOBZO6qCEJ4eh7Lr+vJbOaXQk12w3pMF5qL5z9llIGL2JTlelcne8NkxjFcwp4HnNEEitc
Tbdw/GAFiMQEuZheUEuvfqaxhcwawS5QMqwfoU+EJY2bYrg6TJnInR6ehXe44LRayfBM8n/Vcjql
AKwMJHHtRlQOuz1AgX40i6MKcIIg3hNGo865WZCVgXSjJO3MN7P7utWSNpt0+vurVPZ/QVB+qPtp
TjD3que30tmw0xQEIODfHaHHGvjbr5nEvJJmfW5bPZwspfG/7cz4Dm7Z6jN5yydkzOxX85tN7apy
WuQQrEevfKWpjHWTfOPIE+VZBaxw2ZTRWAAsXpMmt3vomhzm8HF7twscaP94+9c3PXV+PRzHwm+m
nbzNw3Vlspu8nuWdVsC1cgIM4tCJexC/bJQjOUobhSEPxDxejljK+5KOVuqYckmoexflu1GpOKyb
B7XM5urpiR1K+d6gpr9rrpTrd7jitK4IRgJmAehDmq8jAxsq/jPT+Rd/NVHZg9LwQVBhizGAy1BD
d9XFWIJxGbtu6k6xxe4y5QIpm5FPBrPpxlnnW1iF5vFBg2mRnvMEqo1P77bAL5YDd1qv6ntL9nsq
7ZztyS9AjLP7K41R0hxRkVQgURZ6nYOPvg+rKq6j+mVnrI//cFl7Q1DJBdsH0GAo16dWiMbrfr7L
JaHqLJlXSk/3vmY8UYuvZ1gnVbWGyh1ZVRdkIaSQpDXWnXUNLbNlMEwYwqywXzoTT+wqiy5/2VYE
QVzkLWHeBbSCJU65B0SvIQR1nQj2ImXNxREIXb2CrXWZ9L/vU3rA1mUPnHv5D76Atprgc6X94C78
UDPoOHIPldrpyejrLenXpXxtuivSQR+YN0/2epVzf1q7LYCVOokLBDN8Y8pJwvKASQSlHVksV7KD
K2PoW9OuuLWiX2ulQ0lt7hgJ9ATrPOQX3AW8twLV26CsWbsxwfzFwKbtxRTXJdKJzUfGk/Slj95R
rQvmqTjSc3fu0Wcqdnjw+ZVDUl6ons8h35bLkL70YVKlT3+fV851mCenuC2Z+9wUMR9L4/S1oxBn
8ppxM/5VxsOXulErmtYNEpwOyM+dGu7Tc4NZi6ed4OYYgHt1fRLYDx5Ou5FkQ8aCxqD8JXoVDbdf
caR1lSGFU9jRevIr7F7fFyZvOAxNyOyANVud8hqgT57b2dSMrEb3WLR7p+aDGuRcn6jlGc68Ifa+
Et8XhYdb4xsAW83HSThpsHD6xm0umeB1IsPEZefjNtXs5mVy0kVFmuD+2XRYEBRmLO/C5n41WKHW
VW7J/EFamJzl5DxCa2UjiOSHOWizszUcMxoMHsrag5Iq+W7CziNDoiKKbqo2wSBRFhXupwUqi6Uc
66yqwatYqfD3BBhkaAgTPNW9YfKeKHzeuLzNX1d61wVKraUUsdkgYr0MbGdoWD5m3zbULTnUST9D
lmklRB+dhHrZ/G+7fP9384Bo+xvwaN4Wl4GWmj3+K5tdIrKckrpJYxdODPWcJ6kyqI8ASPSWsW5f
BKPYyutWFeKstbsEFYfmDq8dreEPTjh+MJv7YUiBFYXwHv5NWUoPXywj8ArJc7wbQ40P1bBbh7n/
SqjUdm7TgxO8WhXf0V8MOk8M3C0quN2YsDVDDKZq4Mb6I/v3nVvCWTiKt9iZf7JqSh/72vi9pqkC
O8zBHpEO7e+rUddtrUp8BoyW85BBmZy7yAkEfvCGM9B9JOpv6hl14h6frUR+zkiDk7cimKjzYVt2
rLaIm7a5/aF9tLCg2M0Sh2SpS4dBARUSHD/moBVQAkAQMAW0nERmAzVcYZr7+2RmsEAuCE0t+XNO
OPMkJgjyHZqCozx543njEiDysJDtadmDXrc+LRQE2OE2ais48vo8XARTqIvjghmstQvBP0K8l0iN
Gi0uluNeBdJcyx61CRhDsekgWNnXlpHwLhct6yY8hvFUZ1EDpkRmVGMlPHxnY2Qw13m2pJIdEklR
WaWRTUhQIWpSWKqUIciASXBkYxAUn3iP8VSqACUUCTMrpRpCgnHvX2G0GCMdwI++r8EEoQK7H13S
IwieaPA0FZ9Pg1vI2vHaMeb5pvrcMRCZ8z3kQOmXTn3Wzk6Duaf+tQ/eJjfQ3Y53r4GX78qv0QUK
4L/0QLt3nXJtEDnaE9easf64S0UXUgEmfeKw9X3p2zYA4VCDtZLjGi3GWG/4BKCLDZeAo2O7Cabj
DZX3AYusgRZSAp/+aONj8vF/obAT5WKz36R0scLRslsnFtPMJgjBfpDdHWZbWAD5lWsaQRVDVhbb
W8F929IXJPwklIM1KnYhYsO3PJZpl0Xn6LwL4Vm/xULlWVVv+LuzIGApamf+VUEk9Co/Hu39WJj5
Uny9l+sjoA4+Gb1mgNfRb6Swg3GSNOvxefVo+nQq9yugt6MlMSvB2qiY580CcJEJKYRFXrqg1RDF
PRe0BeaKbc6OChpjXTyFc392Ac2yVuN0u5pB/r8+JdGQOvZlHiha9+A07G+eQkWZ6C+6UkA9+fM0
pQI/bUnai4O2LQ30YrdVSs1DFzJTumVDNskO6c2g93eDoxdIQRoyQ1le++NFCTkZ/2HExdp6DhPk
VDXwDds5m+C0L7qetznsxdqD+aiMwmsybBCiqGz8tDan7iO1gOBp8ZHzMc17+wIBXL6BeCyybnHn
V+YHrPI/V8LAzSna4fVRmP4b6mAZUppzONzBZWgaDNTJY0CakyDgmvfbXgC6bFZNB+fsY3qCO9tR
tLwWdAL8vejW1VBcqcnDrOPv39bf2j+8LJhP+4ETmDbtUxsT1Y7GOnqlB99jrXmZQdBw3WxDIz4U
RbTEH+7SXmdRNGqoUn4PhuyUhGUa6VwAEcZTH62qEXjzuC7pls71YU7ZlQKuJIzRURnO0YaEAnGC
PjeqK/9ZzhHk5UKQMBb8jdPBC8QAwGuxxzv1KfWtWXcLPp9pwjgb/l6grllNlU7fnX7HkT9bUU4u
DB4wQxQ/KY7xrQcvsOO4iBa/xIrIQ5+buHvfcsBrc3t7+RWkW1eSioxIwmvJt/AXZOFwguW0PHGp
Dku4o2y9HtVj9UyzTH5jY3K7E+0O972+33eML1SM0699LhzMSvm/e7iKGc/LNuEwDBSQpuruhct0
8d+Ms5tMWWDcYiv2smJKr85NBLUz8xnphaLaz3nNQD/yw5rODDSlEGFQT6wGcP6Mr7UBg3akrvcQ
UsQj1q42JVa5bU1KU+rGCdnasdaBGXRCGnvi54SeeooB6ULGHd1ov7GxGslcBzNs8psxn1gZokM/
GrZBrFUiLI/GxLjSCqZ+4FRO94kp9cXY/fHRjjwrHlhK26/piYyz2RK+t1jAKJLnDgaoXwZ0BrMw
EAG7ifb6C3KS3ysQbwagQB73RqkzfI7+ePd1mutvZx3gFz6pdU+hnI4m9XGlM2WebmaPOpnHdU75
mBw1XgWLiYclSwY8usd3iEfq3bPTMYMVckvqMYefRmrtmG1qF1nGBfp7edPkpZ56j2HyJNAv8v4B
gFjlTXe3qmv5zty5V53uNYeRTysKJ9HgiPZsRydEtKhUkpbLUqUjvRDfH8Kkq9BnO8keG75QSv6J
Nau1IWoQXvca0PNm6Ti9mWDUzzzRRDIIkeTGJDu6pHNc8ZTEnmZ/lXYB3JezvhM0LWgJpHLcuC+4
dnX0stZPhgQePZoTtrhgnoR2gbwsZkaB+zd2ndgnodtKJXxJMPhh3X85r9ubF2U2L8wdguyF6fVj
mcIdsuItIcRfEngPR9+RilewTk80wgcrYIBf4n6ZZxIqBsQ9P/5tAwUUvnVoqijzcmSsKPZ5ik5g
vidHJfe7mnDryMDxs4csNdOByZCjFQ6zTArhIN6lQ784oV7Tp/oUCS8J+bBLxw2xGNxhXGo3Lbqj
RDb86EXKlL20VdDqaLeI/l17V5IB4scRDBu/1NA/yabrqaLA00XHeKEfUAlDVcv6c6n5YZ4L6Bzw
UK4ZnCczfz7T32/Eo7vYKOjURSChhCT/0NDYIWCCijhy3c5uRLzaAgIGeu3e5BBw8WAru9M8k8pX
tBoyUBSuTZDMIrvjvYGFE2QeWjFDCH2hIzI3S4nhP99JgAKSjJsXIOHqgZXW17A5VUhPcv4OtGMH
RaLwda3Cau8CUg6MPStIFjzLW0l6Zxg40dlNrYHjZLWgXwAFY1wprawnQnxpDUjmJIaKnp2bPxbP
Kp/r2aBuVU8p9KzlsA2od12Bz09/3lnsxWG4/wYDZRsAWQ4vDD+/kFHCuXNcHjyTDoaUB9cDZJN8
mafDy6ikMLKZkwW1GEBF6c/eD43ppMnBPaTgSqdW7QRjH7C7yk4ACAFrIkGlLVAfI3yK7nlAnvYI
AWNlUK9xNYC+gqM8vqMCunjDWF2H/cdoWoXPxXH6gxBIvhRI5DTV9SDRj0kZncogDpiimJhJm37a
mqHT1KzrOR41GdzlCkAZDDAHLk687b8BDQLlvrC4y9YpPvxwNlhw5koBnG96gtxmLGzp8F0dXNTq
aQLwHYFYwZZsriol11HUaVVKb7t81N5ECQLzupGBTlU7iG6MhkgRakl91rNkFnBcRe9Phe/rgf8F
Ok9BNJormS/Dt++IOD/w1Se+SdF0t1HcXv6UfD7WYUGxkeiB1m1NShH9/iAJNSGG2SfM5bQ/1vPk
OORcwUYqiOIPeZqpxNn3tDI1Eqed3rIA5mXNy/HJb6sDbq4PITCm6JsowAO730b7bUQvmUkRqEws
7JDJ4gOdLktnA1YFl9bgSZ5SP/EaKKkumVcHVk5mSem5xxtIdwMX4vbGbhRdkujTf2Wz0aoS+rHr
ZZU9K6HLwzEsSb3TMC0EWWdVCZQUPHiJmvsFNc6wH3z35RtLy5lPpdMxk2uhYmDUe58q28EO4GiT
MaY2nb5Tl6tNDhMLPUeI12Vtq1tHRHFCWMiWnsvg29SjJiYsvb5pNa6wNvgglnL1/tMRYLiAZGI9
yBGgrMn4TEfzYpS/vQKrZyr6W4e+wVTvTD12DbRKYtk2zucMvqfBbIDzDLdWnOFhXwt9IxFqFHqQ
HV5sEriicdtsniTiOT/oo4XZyQ3ZU7TJgL7W81nBlEeAkpdzEmn5wKsdF2Q97Ucvgd1mzijVmC49
eOIszlAJ1pPFC4ae0QyVEkjrhfWvQGDVwmIJrRT6MXiwiHpKoOu3F6YnQmyBXmuaGxoT7+vdrdED
295FBx3oQ6erdnV7ucVg6pJI1pysalGMf4czHpZ7WjuMXu5bUuA9IZAmvoOwHOhwxn9juTkBaKNl
zEIZ7Ji0GvAyKZI8DeIvHJPB0pCx+l3oaKwUrNSO0KA5tuJ27cTQ1XbSBuPGUrNTWFtI3drz33l0
UOArPoh0JmtMKWYIKpIILqdmYI1KDjo4EeDqHd2vHeISYvA6KbGtb+nVhWq2hauBteMn2Y2mKP4y
JkSYoMNaw7MpmIB+TOekkXTQ7g96qQw1AEFzXKfNPqBJgUFhc/Gike05IsL04wtcDe/ZT6xcVyoU
V9FqQ7Fk3FoRqLOYMmLzSvmGugnKYTlJG2nADVvR+qAPdMOIUmYP+ysnvHX9fZ1zXbEwtcONAWfF
t8TFkB8iO9fevcOoET5RjloxqN32mEzKL8Z9sYDrTiS2Kcfz8z1y4z9sEGMjJdEd91yhAoPaDRCf
COjUL9K8YAjIOQHgkLTvrkMW1vSHhMzYNt9w0kZRfwv4prpR+CSR3dy2p+3Hxh8EUawjk7E5OOD+
wvBR8MNfDYTK+uBQxxeR+OeSUr6Y69YzMO/WO9VIwF1Rd1T7G9NmsCj6w4vaA8Oqrk2MclT9WQfL
sv/gmZs9pJlfSbFic/1SCwm878AZHCAYmvAQaGLcr7WUI18MUx4eAMkXARChpmDBJHNfNr6jpEoH
QNmRe3bLYE4ZZP1JNrMaKzi6wUed/qoVMX3KcV1Sj5/j3mpfqfUAlVcxcW+kZQg/rUox/A+P5B5i
8kFRZyViMRsiYO0yZRWmclaoQ3/0XGpJ68nyg7lF5QrWLrwjIA+HqswHyKMUaDPnUKZ5NWdykh1M
AmRk4mRmOwKnT6NAd+lMl9ohVPesmAdElZbvSsdB8Xur+dIf6IuDrGbbHPMw+cgFppnnJmX4gOu4
y1IU9QT9bPeOST2Oy+mUZ5c9wSJqMkpjxDoi+Iy1YxGWOXqkFsKj7/xsYDDnRCj3RaZIU0d7d1J/
ptEfCPeuwIevNWRP0txicV5DzCwa8Dct0Wbfd9DwZe61y4TkPiPsJ/wxhLUJeuGFGMcRaM0VYD7R
EhefHWfh3hGfncg40Acod3bMeyD9lPkt2cD6mdg79K90fyCoTrhgjJGvWvNyzd0PKnkV1SgCok/Y
O0SJvmvMbxXl0Tq0rfzMP5I+8YUb27C73M+CKh2Tm6ZyGLiZAYUGGEZTjEfw8cvPP4X0v22jMkaN
mDutrrFLgY9AXOYbc1FFQTRuCsNSsYyNIGnStpOHhPHJzYOhyKTXbTMl8ecI18hXHPbeSxCk8c4T
Ne8hXqT6WtU9nSZlRisFcxVdfsh7wxu8QLvgTSQpgbMYD0lxRSlLBpM9hPAu+MqibGUiP6ce4r/l
FT/m+slfpdB1YxA//IwfiUHUVcSBwN71nR3AyWfLEWKE3RULfd/t4Qpg45GW7UyfHcoyT1CS72Oh
hx2tTRo0ab2sTftFvpgKrVCjVe0hve9MTrhu8D836ayyLc1+1uOYIw0uixFcaVma8Oy+iaVif4f8
wIkdRGcby/d0wxlkI9lbsLF4/toOlFJr6LL7cNqpC2AQM1zn2NmBWMt+vhVg0Pz+1s2q4zdAmydt
JLsMXsK7REhS+ps778HfHkCVRrOfZhsy3SgGCEIHMFk9jNO/zayrmfKraYbV0gjIVSQtylPDU9p9
ykeRh92X1nyqceQt1PCwMUZG4FkgUecmUya3Zwpo4GvGlv4jHjsmhUsT7i/h/Y2rxIRj9X8Urzdi
1ec5Z9UzTVnBBOXIVF95tBRahgiAZpUKbGMOMpDEsZIps85e+v+qFJLs6aaxrP2VkyciShZtkmOX
DJDw7wd88j1amvZOlfo2/Nubx8iQeUSZlNaeb+s6m6NFNr12baBo7dEGz/WA+V6kjlpX7nkmwVCU
LioqmkSbgBw1rwEbnSuP1vYAYX/Yyl+NYPjIqPtI3BPbTt3zmlBmCtFS7vjKxSOu3QogdpazmfaC
FfkdmAe48Hl6dmVaJZTBGv0QtGXZ7DXcrZkJy1Wvb3dD2GPzIDGb5BsxpTJJU5j8PUq3Hkgg3WtJ
a8oLbg8kFcTkg6UkUQyzcMW5/VpBTBYFHaGjXgF4ru6UropGMhdfiHWBvDdBj5uY9AiW0Au9OQV8
JAEfhPeDG0yCZFGVgbPE4Ygxw85qEOxTqQjbXQCcCpybvALQH4AkU6J1RD4wwfDVjTPW5wFKspHN
JD+qSpJFQKZRozB6X22v/ZHSdbXOd4TjCpTAUxhff2laRBNhVp/k2R/dDu7Yt/M+meQKfXIR3CG7
c8UV5YnLoEwjK0oh8B3zsfeL1d6nmbt/ZO0HuN5tHDJ+UzSUD4DlVSPEYYoFR5emGqeUD7VtJ2/Q
81dREPemLiKLRO7RsUUKx4Vv/HJ9sDq/+Cf/WBLGwxb1VAHaCI74AcBUrGwqpNbHYo0axMv8ildY
dKeCDBiFMkKPB3x9Qa3c9YL/8TeEG2d4iN1v8FZ0jBzkKbUocsx6FKS7yLNQDpBewHIplts+4ykH
LiSiKHjQzw0ddmwMf5W5KuIhLPg3QJZlY/OmcsC53Qrb+29Pisav/3aRK1PuLKzDC6/caJxXQMVf
pY74QSc/7H+c9Z69P9YreoQMk9t6oxcgh6w7hEI0Vssf1JZHjqBPoQRzrUXEXLZ6zchJFEy4Uml3
XKTZb/KYt/64swB6udH2vl6foqbf/0dJOkd87aYLh9BrxEfsP6DKueFBl5TEsX4xNRjjWoXcUyKC
C/y1ik40bDNZn289y5G2oPV+rfGKy1cfNEdsVGEdRWjv0d1+LqqqHAU1MGMvYahbABONhkFMo+fg
eEgE+eATd6sGiEJTCX+M9bdb7N9B5/JiM/81g3eZLxOq0z1sBUarPSUJ3lNBWfXA0+h5qoeOR2Pb
7YK94QyqYbsdXYzTlY+b4sgCLhsRnWQ3YJAcC4Rcyw1IP97sTLmKYEi7eIGntSeXA0kPdabbJi0d
XnATB3eJGge0vlCAcQgfhHD2QcJQmdNIuFFYAv99DcALeZ5PdiO57E+KIgjkO2stUv3veLhPfqOT
+2f111jSnMywVePPds2dpuYChc2deSMN3Frg27xQHxI32c4KUhLprhekkWTTmnigdKEjS2/HAr7X
RgGAgFY9DLU9OJKwKDq3nTja93px0bI0JeqUNgSNVgXiHQs5MeIB+A3Cr/l1YWq2k+MWDIRjD1pV
pamwRy+0BUvJDWPfHyfvVOUWfQNeoSmZ74zGnBGabVX76cln5RUix+qSMHHmCg5eHh2bolOIt0lG
iQU/VP7CIazfi2qOodcXaQF1k/2bdeZaT8daLB04IKI6c9ElAs2kPvnMDl/woYlr7NyWWeOaA6Jb
sWbvg2YOmx5CNP4mESLAZCQDdlsdu4ABqe4rfw0amvuBiSrormZLI8lw7zzGdzyf9KGqBLL+H2gI
fYBdDE7qXClEm3T9NxnCy9EGRr2GCKJ5zGoN1FnWpaqVEAX7ijxfHZ9tbv/481YB4Df0/vLfa3s5
KVz822ElwMRMmpkYBd1WVie/BCmNb4I+xppfgfaEoL4R7UyitvhrTLGQwcslpA8sNIFrDmoamPWI
AgO/U2fnG4YMBq+mxQUHCvvgdaMfPjg3a4XKPlMrq7qO63754MfEBTcBk3+Mq9f9DcdHoDfL4Ltm
m2YBae0zr1K9ZexCHMCR1dmbPeST57CEKCJ7uU5oDI83V0AwwDOBxOEYFDlhPLMY6+ruxK/wS2OK
NYpJ3ZKy4k224CVgoodj5CSljwgqEQZz7hlHkVJlBsXuh59HnJmUvWhE12vC2LRZxaVW9cZVJvwj
syFnO8142B/1FG/RrAMi2NlKcIsRwphoCmCy1uTn1VwpJ9U6RrZOUvdseYbnczJ35OJsKi8NEkQR
jlRhBIH/p7H8tt4fPoUT8j5JIeqRxVpa3oyFSReLBQwbp4KRfjkp8XH9tEDXkH7yIyd+xfM7S3YR
wAdwg7OVehPYfHZ/OXB2jC8mK68290FFzfP7mOdbrHl+g6XGdGZYAR27PpsnP1iljmiHu4CeUO5K
3oL496bXZWERCNV/Uq0FCxnY/uC0xeT1y6+Ua+vaMx35By+FEjIbKiqvSioe+ge0tY4NpxtmzuoD
8RKjQUYHcp/RSw82F/yjcFspiiFw6mzppwtNcKMACoh4i6PiBjHOF855Adt1plqiA6Iqc0ty8ISW
PzqpMyl6b/kHx0hiXTzN3+qRwjGW7qyRIOL+HPOGjyv3w+nXdL21SKwX8VFMmKvX5w4qySi0Ca4y
5cv/CEqQ6i7qSw3RczIu4dBoB0jOddo9SpKYISjhJ+c8BzESJYoCnKrDMNk7WOxSP0qFaNxH8gFQ
Wx8EYLr32KUzNL9VdqFOuxq5/erjZfMWLRzeqhu371IRUrWyZ9AByX/DnJuytTDuQSHxFTntjxVl
eweVmYvexGFZlmN0NRZoEXJMD+lSzXRHRwifGTX8whCPdxciaOqu3bMrz47N0ZnC40N+ou23eARx
futoQFHY5x0+Z5zgDYRuNWg7xONpoq9lEmp4SgMjaoxd+6GBTvUNdc9ZEOIek7hbrE6JVr+NKhJa
Sw/vuHPGIQVDCbm5RELppOpcVb1kqCHP4bx0+WKGqmRVoHFmulnp2ByRsdusjZ3d+TEncTAr9746
F/d1LbHH9X8xfNQ8hBiZ5kn77U3IcbQikcpiyfS+DVCuwXKABBvan7zO7E39TbrRnDlf3cXGEieJ
scwUmlz9gtK98FZF56wrAbO160/0kD00iyUKGgW6hhS6/Gp76HtJOKhyBrkgzZK1/Um5PJwINQH/
Hqt/JkWv1pYKW1wN4+DOuwuzgJLNfG1eIxjFf4E5D+5e/raO5eJY/P3vNgQqahG5GKwQFrcLM44w
Ap+LSwcaxK0NE2ngvqbIUaJxOPCsB4p0HPHVlLwBi2flSyK4ejcJPWNYkDgdc7g/z4E2EX91G/6D
ZbGtTb/B5aLT9LzRQoM7TXSXsL8n+2JXRYrAP/HBB9xg3B6dFOG0kKp6Ff6ZFJgGVLC2Nt+Ms7Yu
oeJBjEAtTtG4Fw1h6MpalkK0OHWZwPY70DBEBj0GRDsqDRg2QcOvmKv53jlbqEkM1tD5TNCn0+wQ
VOF+SMjqzI5orvLP/wvdGf3OqRlYDi5jVfrq/f+URX84ksG0uUwY6N2zm1206Ws7OFe3sSvYF7PI
Llnb2TXbFzCDJnkLpUtYJ+MPNkfuaE1Sn/KwGZU/evauNSN0WAOMuB7CwdwcRy/4YYOGTW84LMco
0O+ncPq0PZv9BE92sq9+E7iEiJt4LUuKvzlh0b7mceJ7veyB0WZuwJ6NOBMjbPetrGpxYVZwxk5m
+s5X0uK8VlDH6/46fUZIPjgYCRaJUvZEzLKoqKTQim6mSNmg7KRBK5uzZjxDBlhH5k8+c3hB5f60
hDCUkPwULYR0DojinWQTEG5ruKGcT6edHCbV1VT6Zto2PDC2pGJdodEahrYhVfBvvYnDCquDTwD7
ugoKX1XxBchW8eQlVM74MQgQ3Qaa07ytGItrDZSjfg9mxjOsGU0AOYLuoQuLDauUnCsGepnl+XJb
8Xf95BwqzlPDr7DOJuMKhvJ150vlD2yoBtEx7qAw5X34GBue4XNbvwIKJz4FbNpP3hufPX7SQKIb
OIFqF7mg8l81vJ3EdWrSkZyale8QXJCz/1J95hGBwAGUWtDBKlhqe7UJzhraJPfTdBACnOFcpuPQ
xnit2H4sQd2x7YMLCdtc5HYXmfp+8Z2mOS5HK90x/99kTzOn5ctDNyESTNgPB6TS+NKUkUKsrQb8
gQGZJ6Xs+7zcInDlohvzEXB+kYEW4mO/yH7i8Ps2VwzBOPRoM6IP0p8/VNsRp+Om3XZi46Oor1pi
9+QXlpc+U150QedBZDMmEK+nVR+HAPkpaAPNqcwHIMw/A0nKFn/Kbi8MEABgE4wz3ZXf1yBzmVbf
UUp+jVU0kc5mgemkpEFogji2QvOufr8nxN4AwfjIRlNG7rrP2sRTBBsXlE9FzDXJBzHdBgAsubUP
UW0Bj6rkUcUM4gYTJOYMTQwUq1p1vjsdQJ2p2DcisTyWF++QGdH7HZp+NDV9j/Ah5IEKGNX+TYll
YXFLv7aHjCh8oA5IjiGU+XEbLPUHQDWHm0BjvHC0L7YEbFwmeQEixkwkTuEpdWXqJ6dNzWr3X20d
qPT4l9dLV6wdQvW/X/NgbPPFONdwaMSnf+iqtHIUIt6/vJMrZfnZxYJJ0gPpn5TKvkiWH8iTJ4ev
UJ0g5yUfAGqtS+nmQLCFlLEOm7c8HwtxF6GpwKhWijjiGbu+iiKTKchWOFFC7f6oK1VX6lwrs+4V
HkAfgsaYm0StWFegGikQ6NILmHZQmhgktj/NwiN/8jxh+nWfIOHa6KkPD1sq/isSxYdR56zczRzE
xaH7bniQEkWyq2+DrOg48aXsfZYL3zlZwjK1SF/j92dUOjqHDKYB4ihfv5AIoU7th1UvIzD1XBp4
doLILjo3aNNAcwaG4CjA10kAuyzJdhWUPLsIg0m+IMUSVVXtl8/hRFDwB5rmrq+gt6/X6AyB+1/u
00qFBgaRICgPL4yn6rYyY5AJsmnvwxQPDoUOOF4oeyQDxf6rcteFIGhegAQuCsEAV/6OiTAamgyI
1icmOk08qAIHJ7VCKJ6MvKdmlyR+k2c3X/W5bAWPlg9Bcfsc430XSOQWV+uttSAsjG/3G70gmt0W
LUnV3OnJYccLpw6qDRsDCwnXm2XHsewJRnnAwfjkbYaI7kgMj1t3LJhRmYYFI78H14AVszojQoH3
yLUNeh0LQwLICX5ozXG4R4lz7X4C3jwxmz8dnOMBvSF73rrJQ3aWe2i/vvAfGACg+GtA8BgFbrFb
dgnCrgSUCJlC4HJJ4uDQ7BhZ3DdBicEoVHp3JfYI4PCFrfuv/yXknKksJIBYU3GOfQP+ux1YAtnU
mj4uKwoAlx7UlJudMPIDA6RE011dHtkDAT/p8gY4EgGH+3aHSspOEoGiNQUE992dnlx12R5o+/gK
4amIK6tw7RHqMTNaggNLZm+vxF+lKT76o+zhAi2+IxFNii3SkchhBl+w1BI8QXvQOgqLVYfQPckq
rxjHQEvG3pJP5bkDU2QjiMhaaKm3mHXQEWb8MK6Awfvdy01qJNFlQrArf2mYGryGYzRxkXAWmOPE
ZRvL+9Tm5x+QGdbuaqfADZ3Q6nwjM/j1TjOeNMyf4Hqj9c/Qxga06uNPx4J/CbGkGHz3DLZmEqsw
7myeczC3/3a6i5SYJJ01LJA88WQKUCv9X3k1IpHnwLURE/ZfDK7W/yw9vXp4jEwczlfuV8S7iBCY
ai3FBovqIeGS5moP/55qO7wHyAyJU7jUYE/yB+rRsAPejOwqWSGQV5RHFK1DukK5tfnslfSrd1P7
JMirLMkxNG0qSMEag3Tw7dy+wxqipfmIKAZIB6Vdy25uGDb2HhFBD5s0e6rgYBSh9nfYqRii/nsI
EfDY32lcpKlkgx/nFGUc1kqdZLvoPOFp/LoHVpDiMZy1mMWkZIAyhf4yZMt0zzg/5ieeU01+gTJe
mkYDURpsSK/cRHrk+RObixMeDo+2zkF/Apf9jCfY4ElZ1ooH8XSitojA42Wc09OhrJ/WkTsRb7S5
tEe928W0VEl+madN0Lvsgwmw0plLbwrGJzKj6+fgZvQcnmTD/5l4jTzHQ0dnoqS9KUiFA0jVVx4A
PBkyfFxZFDTq1S9GaQvsZs2BFyplew1udL0KG9zT8dQe7GDSPrJqgoPU24T+dOVHsujk0Vehy+8F
hYeSxa/OVNcwq/TWKv8CG/PkhX5qDr28z/PD9rxoPn5E1XiPTVPas/ENL1jErZQBbvcGFWmK8hlT
P/Sl8uDUTAE+Yh74oInVCtGKmErj7S4/xxc/2shbyj+QgNY1Eb2dq7s6SrOWs44Js/FMVqqJy27/
V3L7rNu+5U1A7qqfAPyBYyVHKgfdT1HYZBGLXEuQ/odepiyXwd1aAQgr7783QayawYSLyy33gbnc
+wULg/bTiIuaIdlDdakXA1c9iD+TrtwosK7r1P2HT0yEa9EfkwN8nqUp3RsInziYOwi79koTemLQ
wPxBGVh8KPxS7RJkhf7HOmN2y+xd6Ll5wIXxj1Mc5sFzAIwtNyyiX0zct+7D1DLAhxUbs4UvFw78
ODGLsLHmHXIArZpWJ9gqjKTueeRP1rztSZxj1YD5U/DHbK3AX9cEP7rKkOASSaH4D3Mf7O2LW9sy
g0z+TsD1ODoPVJTvkI8vnSVp4q6iXSVibgT2BsMCOTGscnD6sT4t51XY+OWmu9aBCAI6YK3S+v6B
0JW2yUAKJMZccH7K+9icz1egHjSq4gbejWDeYnbkHK6UbqRRP8LKVsFxYR1VyfTSW2+QHtbkFISr
sHCkuy8uDgNygEQyG4o89yjTJSpIcclmwq/UQ0M5M5go2eCwxF49e08lfakjxZ189pd1QqsvTlxX
znz4+NOljm61CgXd/RFxEfRsRENSRstZknLLY4pafeBt9KrloxyBHdvc5VrR1mobwMaFssyX8jpG
Tuy81wONQjw5zlXm78/+EblkXfhb3AhSymx8CNSSC6I0Or4a2fvdrsowp1JO6ZRXcZ9H3WRKMTOu
TlCuiR7QRF1kQs0+PLJPmmBJg5POfVw5pkZKouYH9Y/YC34JGdCRwytcs/C6si3ejXeHYBJkLtoz
eaJyYSCZyyPMTEn/ekxMCH0lz4tev/WLSqh95rBRZqx5t6HebVub4Q8E08pZEy6jwzbU8KXD071V
UnxeZ1Bnc14IV0aL5O/hX5l086N+xDuX+gZcw+Eel8UWEOq1In1JexTUD4/9+NJAs7oHNH6uZbGm
EL1QbUTRtPkt1PMTjssnWptviS23ZlQP9QZ3GaKOs1phutvyPXtGTt8eKxCvOKm7ZhyGGAsXXlJ0
D9cYCNDLAXZlCw3BIl/pX5G9nBZLRIVtaazqZ53H1rHGh8xJ0xK6j0gTu12NnO4QO90NXNMvfuDY
FDlnNR90UBM9jkcsc0wKTFMD7931ip7w6Vx9gKsOGeMMr9MvXbas44hyatAPFMqHQ+31aM9D5rhf
QHsFEXmYJC06cu9Zhc/shaM6AoGgTmK9Lk2JxoNUWaw7mxlq3yh6lcjZBNEQtUrIcQ05jXvxiEIa
TXlLHo8rp1PD5vUWHoonGiJ2XZ7LJHc7EdkKLjPWkASxy7lsvxEIYobCLhiE7r4tVEaV6nwBSkeR
6uoN/FfF+Bvx3Bvg493bWJb6opwCr3kyOGFH/8ooPsrAnobhi9NEJ3uW7wXxxM/VLPYbgZbf8bL6
3KC8Din2zocZ4L/AD8X/BBW+oiUkwuWeyhTvvrecxoP0rmGBd2+/iRfVrHcaDqqZ65Bm6YgMoKwG
hcJ9XZMvNi0HVi8oX5wIy4mqnU3sulyE3KEIB8tC0PZipYcjMfP3GR186j8EWNw9YFfgXL2Xdk7i
mLhLTXJNTmz1jJRapprMo8Dyiv8kOnuni+Yi/LBjjf7kLMjM5Ro9Yt6TskQg6DIarFU4EaQ0C4N1
G02hyWMegEWRud5+oLzsdiE1G7tvM94xM+JG+djtvY/4Ieff7mfUNQ7nAUCQBNS/rZEHIj0Yciam
e/70IxiBWLOQJGWBpbNB9UPr/MiOk0Jg3vQzjUyg5GpxoLjX10MVcE5ZhmSpgN3I0cYJ30vKrxDv
tZGJqzJ4PysMm8e6vqx0czqc5n7rF3gEEz9yHVqj/1kXrXE93lKNqD4zNAfZUcDM1uKwiDWmSF/1
ebbeImvexV9UGafRildOuOMy46sC+cGf1vs/AS8ZbUyx+poLb1RgoX6EuimDzvZkt+YmkenHF8QH
Gk6i32PMVfzmquuIe4eOMkt7bqef3ePirCwEsU6kOR1/gzeUM+QwWFf5NGeBJeR3Xv+Rb6fiR0aQ
A2TwGG3jmDhPGNCuI9W1iH7I0dUW3ToNV5llQgS5W2jfzOT5GPEkFm2Q6S3F2rC5G3BytHmDNg1C
hcCfL1r3VSeHYpLOPXEtoz4dTiOgOXtTnypjyrcNyoWqLgwYWB84dJmJCyN94yjqQEzubhFUw+hn
rc9JoKOHDJbWKc9kq+DoNLMWobtldiyQrtR63s8aIpPpAgH///0p7SANVwyZgGio/6yqgu9rM9US
c2oQ1PF6kJlU7W1SesDfO9KC+c8qvMgCbFnmkbg94ify6THXZKiXJGCeumYla3xHH4C9xnnj2ptZ
2vDpWMcOxdUHaA3HtM1MPQVzYgT4lLl2/PI8X1SBca39kU1IYMdF4nU2HCrKD0fWWDO8ONO7L24t
w9f45Aov6nEShm7H1BRDdwRF2t1XRhrFtc6Cy0P9K5G1HVdZyvEgj96SUxsND0YH85B4ekdFySbW
PIJXGyaRALSsgnSMWlLA6UaxZEdar+3tXySyjk+4vQ7414Q7WJQqC4HCXO1G4xbuiiIZr46zY/QZ
+dDu+W5/npJWoJlM2CRdH8UtnBeDcbaizrV+ZYvdTgfMMDMkGgWX5sOCaXl4rnI9YzPIUjeIMcBh
ieCg1HVBIuoMokqTaVOKVpmYD/50UF8106dJy6nDUKsnOM7S/H7+bEn5xm7Lt/qK8snT9n42hW10
frTeyET88pTuQepmYCqMWV8JHr5HCC6AqSonsdphrZ03bsQqAclTdReMdjruZFLHH/LxrZRUE7E7
UtGoSUvlPb8xXFKm77G36gz8ZGVofceF9QdnQKxV92tC343e1O+43U+wr39SeTg8o8G7KyHb7U3R
Tqwr28Yd6rt9DtZOOSWqB85nTF7/PmEXlUgmKb1JbmzdsXNn2NCyn6xlaJETdZuCgicAYV4KeSq1
OuqcdJePPLjrFHMxnAzI/NHjnaUPK8gvUzpt7+qTUD7ik8YOZOjjXvo3Nfxj/2yqSKVFtvwSWqM8
j6FSJQJu+jSkh2yImV1gySbvItR8Qa3RNbvdVDHqWUIgw2qfkpqt3D3OazgcqpVhXdpSFvF6ez3T
4zXcgxf1GPT92M6MvzyjMiTohn0L+c+HI1n3u7Jjo4Mo/mMq5zYw0IJcXhzCol8oCaIomuJtkZ3a
RTaklBho5UykFFN+ZZDscVN6KIc4cprvkfdbsDnScrtMkrEZspKLslJlEbxqyAwZacOdEURPzWBU
khv+CXgWdUf2FkAA1LedG8BTt1FMj5skBBM4Gu5vfWRmVzgPu68Q8uLBUCSJ/bwkd2sOn8FjlYAA
lMP+5pkiKXDrP85RDoRtIkXy3dlgOu6FfhlYIogmYhWdOtRkmDI/lsqM35QLlOtJCzxa04KUuLQI
ebCbt0WIuHpasV7wYoXig+y4P/PdNbW+z7zANrUpKQLY+ArAaFSFmzKB1bTuctCvFZOzl0rrf7iP
rvquMZDww4MkZPJ9OLrV61O59X3WcNz67ltD4wqcxVProXMd873ad2WXvRQJ4NsQdntoY2n1babF
uxpeTt7qXnOmBWjDkxT/gsWHkcPhJuh9rfTI7oMIARx0v0qveYUZl32qKjmo6cjbgMs0qGXFzHtb
ktbR5fwJUuNO9K30BUGICGoL3gd92cws/N9nLaD8fEkeCurKKA1FvJrct/YwmGCRgsLRxug6LRMB
ypSDlNC76+LtQXLk3rjV6sskk4mBiCZDDzs5dvgCBzq8BVb3xjV0Y1CCQO1y+/UHrEYbBY72fHRx
SsBAbx/fa4PDcwpLYWjLRV+rqaWafPWplRqVSrXVlibOkopLKOr/tDugzc4+tKvb6T4m9cTlbmyE
vIXnzUCL7Ta1CAj6b3wDl69lqilyiHY+KTWPG7aDhl+/F99OmI834SF2EuAZxLbkWpjvVeNrk/XX
k1c+icEfEafXS6u46/Z8ErVYfgNnZnPeIok8N60JR6AQ4RY+KWXKwwIlU99EDMCMqdvp2OEoOdPC
Rx8LnjXzAiiWOxvPllh2Nf7AxKhr2eZN/E7fhqMkS173O7cBjee3pIjQmoDR1z5Z3YZQ/l2wAABp
KwG85p5y9v9GlLUbwNbBnHMGWayAy3lG2Eto2zB3KXQmUsF5NXlbFn1o1ZAFrXyGY5+hKcgfTAnZ
/crk5eqPoMwFOZAFNnjvvGLHA/zbj2/Oug93sOsZ0x77WX2b41XqNcLK/NLTtNcjB3sp7g0JLRst
qPPhYd2XLJMLNru7SuPtYCc5phOpnsk8rWksjsFeddodu4+GBYTX/dmVl4AM0Dil3Y7hCO4eLJZ9
i2/xaaCAoTv4Ji8e5DXJJspTbY1oznbBwz4Qos8eSWFlzFmulTzapDbvPeBH0W+sc+eZQAigL84F
32WbrV/rsy7TH6BUO2ix/E8DvH+KAYjK0bTQdmghmXeZFwANCclunV6dfyfubq3nkzhnAIi7In8d
1gw/HRgPRp+P3DnRIDi5USpo2cy9VC1cEG+HpyuebZ639iFT0OmXmoSg9qf5Y1YmoFU00EcmIpPP
cX6hX0O4LqiH9gWkYLAc7sWDenUuwKiVIMqXmhGCXODZtEF1pWilgQXQFxpEasfD31LB22NKO3A9
EQEMcsZPRbNJFzM5ZYkvfgsIcHEicrZDrI0GUfFg6V5i4vRn8flHVe1ol2YJD6wjUDRYCF4pUu+J
CaZP/EdloWhIurO29eJrY4H9r2KdgcSX345CPHYC/OMg8XwyvzYlKScEetVBRF78KiEVc7Jo6eRZ
KNvKQvGr6ZO50wmE0vEM+MPVzJRHfsXQGvWiRtweSkzFBZfigOJADlBkrwMTACm7cc8vgNbAopvC
H0neejE727oMvCufChcggb98kaN6AngTFizyHqMtctG94CPkVE5KNZLjBBzyHnLRAwkZtUYFWn2X
xeJRGcGkJ951cNaDpWQwQAUGZM2362QiCvU9IFP2+A3pG5sj8AlSyCTqLRFTuP4+c1a5Fas7Fy6q
Oe2qeE7mlHn3iCcDCPK19mtrhdh7n+QMsGrbaZNQ+S2EKnPpkWxu5/pxzyG7h6m6FRaIh/lklo5F
GUwqQrVF8S85h+PXJQ9rUFllhvK0bDDWl0c4gM0vZyEve/ypaUY0ToNacQgXWlxp4+CLTw6vZcEP
Nkvsd3/GcjwlDswHsbDY9bIbivnGi/LhfWavidbSyCg4HncKlRdgifiXlYjs7L2UFshZg+dichCQ
bPmac2XohE2iNTK9D+4dEB0SHuNHpmW7HW2B+BDIuNhoWIKRYKdG6u1Cn9g7n/lvVwq28EexkHwv
Ue/tiUVMXdjBPMjSYgMymA3zNMztEhwUgtikdGKqiR4I6CCbB0hwvboUQYKD1JsNmzCzgqHvwa4B
17vssfFgba/r2mxYRkL4FUZJXX+/M1NCD0OSXzv0JUVJv43cSbyBfQPebrZ1qkLvAn5tbMTWRSHY
2LGXAk47GRfZIfwpd5YVAok3cFH97yMFqM/orZRSAgTF4wYfnyznJ2YUrVVpt44aLSyp73DdVcJj
vZxZfTCAZYwAeGswLyXmlVSEJTj9SdoL14vt1rrG/iZmgj92bzGeV094/IoH+Zv5Hvj5ijX6uRAk
7b7jU9BvnJV3M8QurDXk6px1EkLWDymCucVjO/j6DmHlAMgUSaDUK7/RmfrJcjvg01mc4rVaqAi6
8sD0AqwrociQh1LcepEpLIJCcpYLiRhqLzzlMvd/CKSW62cmnD0gJ7KxKAp6Un4DFlIJPOW9dz5s
MX4bNcI/3DZESjiu5j6DidT3liMC2MjocLL9UxDjtv6SsbLbAjYSTmdc7GKJMUS2wrtfuC9kejX/
LdcLr4cRlCs8rNDzr177+iAjxfs+P6H5bNelqzU3TT6RrkMTcACKem9ughmENNc7tB7wmtQEE5O4
q9MXknDS/EQfyWO7GkSuQHJ+hQZy6RXWY72X7uH1yzRttEy1N/KghcqhxFDDlc8q2HDWQg+SEI8Q
eIsfny72c6OwZ1C6jBqlfAXtT/fa9vdr3elLWOaM6FrZM7vcV8JkrV81HJfMoNeiKyx+DtYgWuoM
qu2ToEEhIF7dvKDdtDy7O72sNcQ6MU/YCb6kmj5ftAQo3AaNQkTvzwxv75TRFCU2qlioSuk3g9t5
ny3u/e+WlNm0IwN4S+7TvdkxYf2mx4t+pkb3pv+d9zNf8b7FttwvMZblENk38a2A37s9mOBzEJyv
BtiAkOyZT3Y+HlEakRTTh7CwTjPZHabJ1X7vgpuvCZcfv2DVdgOnxUJOC30S+ROPcFDoewdPE6lL
rTqaAB5JbrCiwwPVLmda8TzAiv4Y5OH5w4cQh7cPo++XhNWwkcLf7yAjmrhd8Aagnz1ft4KwR7at
iZ0kR25iC5zWNPJBj6YzF4xVa8ItRJQYK9DkIQaMGwfJgYPLy00OXzA5HDfB9pnIiTZ8avVYVhfd
LVKaW8Igj4L8/KYz6T1ns60/Puy8a698qrdzhIgwjebE2QQNSaQMM2T9nbTh4CXAm0+NrhDafceb
SOKtBDvTZ/W3rzZdynGg0fTK8bJSQYoTjZtsCOd1y/fXXKzR2QzTvjWe35urpw2COeSI8HfpSePI
mUeYy7oEpLTh//YSVvK9CA1Xs60gS83X8pE5hlbCd/zEUOhImVr8wkxuK2r6D3Nq7jncxHU7YwKb
lno1GmvBBz6gd7trQDr2EuUgGdLNRXw3QxGcVdbMZ/rSquZeeMMFZVdo7bnQ7Y05P1I0eACqaQ0e
EScj2RMk8bAJFiZqhrW2DaY9btxL0qj6NfYhtDrHPgEpzdvxnsQQa8kH1Nwf7LeJgPS1WCxCh7mW
n9aKDbauynJnPIJNC4s+Nv6U+iovRgZkIxoN4ScH4GUAxlLybg2CmfPCZRwKNPF+JqF9LVznDnPW
oZPvjYIvuOLXoJPBp3X926hpd0xP33C3JYOLmU+YYciuJYz+0F057yn247X89udeEGY/U05m1yEk
97ZSRMzo1CRH/3I5/+7eNHmA/+BbWBHZySG12hXfEwsWIXKeun6H1fuG5pTPd7P2WtNXr3yhm12X
x+oxAxkl0hJVZzPxe1u6/ju4EjlZS2vBRBNjCw6gJPN65VCIj7Yg9bOo77FMJbn0EV7bZi3NpqJ8
2w4HdnFg4VQ6QLo4vB85V7NjGQ65MpH+jzHzdchl0tBYGfjmwWflyMtLBWWtts1sBF/8CfuEYMG1
oqEb7WY7X/hVEl0xXg53ooY4R4555r8ZZyN6H+if9TGVhGuiiwLNO3In6KdjtwZa6F1M1s8qW8HA
8x0YtBulgvNG8O4QRNFOv9igfHluy6rldi1QLSnttGScIu79ERPGv03Ec+zViqfqNOPpTmBnpIP+
eFBiFzH3IwIYzjXJ4Te4gd508CK1zCIkGhtanhv7H4CIYK75m4D4X1aEB01RxwFFgLSRCxxuu51k
3PeGi5zeJyaSi6kXWWr+H/pJedxJRX5HokZtL+Ms5x8W5kOB2RJ4hN/3RFwOry7vOKGIQ1yuc0LU
6ALw4QVTvh/kdhDf/KqYs/GBb5FBr1gvvyAwxOHyEZczg+AxVuJNGd+yP2XA5dIxjrYI93Ap8WJ/
VfLakTzNLugeao6zPUsMKC2QQhqlKVipZAaNp93B8/V94MLDpLtPYNuk2tDEGbg2C0CvzqDfinRB
QmQoJNeVFdnc649gprXZTxrFaOpp1w4YK8i5yeQrpRL3CwQby2Btf5ajX90mquBeD1116kEjRsvl
oxsNf+8JriwxkdXwNI3ssRDNgkv9gKvMHGwIfHsBWkQpUnml7ylBQNZUntInDYAqH6IQ+T0KQ62w
q1XSesHJK3HDWkYUilIPfJNBm5m7vgFPNu8i4sTe2ik6eS0hFxKNNsUWoGYJCaWY+dh3FaiYyi0V
SWn5pV6TQjljbfmee23+8EZuLq3mYoggWk/hNtHqjLHX21VtoZDpnxjJ9KhaW2Osa1gBGHs/BCEe
ZwllGuSYlJGBSoDJti5NI5rhZUyrAQ7zYJrCXJZBBQ/rDjmT3B/caPgokyaleMnf+tkJ1eTVfvnn
uQ1NTHlILrHolgHdV9YumpnkUOYGxfqtY+GMRu03RE80GqljZpX4qXNVLfR5TbW5ZIvePJXLnQ0p
DFX9nsWB8ENkEhYlPS1qwD3wsQ7QXyIqjl7pWl3UrkrskxcigdpUMlwQ0uTYgY0fqNK9Wpl7wyN2
crjmTOpqy5pyOcMkfOtLodCZDFIZovJgioxm5EhIBcGq373QPvyLUjlW10lxpZEMMqsxSf2M8p7c
rnPtIFj5JMDlryw/5MhaHM2ovgDRBI7tOo6NaOUBQEHF59lhnbhoHKqD2hDKPURQ3uIpmg/PRlaK
s+hfxIoDON2slT0+n+Zmz/vnFXoTcNQRGx/OP/pCssx6sDHNNhuCV2xin4+BMyZI1yRdZAAdcBR5
Hy/3/clXWJZX+r5qOQHkj9f7ZGKdhwF+oHxwl7Mi8NU+iR7OI+ctpO92oksjn6l6zU5o2/rReyK0
BezfhCJKAb0hX/gKdfuW3P5d5MU7ojAYMbC+/ihtzFq0EfpQ2+TK3yJIdB7XBVE98ovFcvxYxH2z
vjngNpkea3XdM7D6iqYl0PoCsNo8kzyaDtLA0khH+V+jDSEGSLDIw60sdjPAum91YWIY7KnXO7W8
SSobfL8XmKbKnZ2rNm5Uac00T1B0iYWSeVCbnii47IPWdTyHyM9No3/sxRk9qaRLezCtDnp2Btum
amWW/ozd4L+E7/U8BWZ2ulCl8DGukqpqxDeC5zbOPKJVZpzif/JDBjKTKe7Ky8Q4DcivkJC3adlh
200jKXm2jjcMziSefNW1LrjYNFXl3bpJKEOr3yUM34+lkTKQvPnxzY2GbeqEEiK6avyG2gwZT+LO
KWOa5qE8hlalG9DQWvPlJ63Y4SkB+Zi21U9unZWIyA6bUtGh1Z9ZdCTkM2GIh2gAKMOWlvR89I6z
yP2U0i5SbHAwKQqrsYdwnF5JvLoDRsZruSca20UP51sQvTJ/DIAjuVCuZVqYMRMUu1yvWCivrRD9
wDvu0Mna2xr2LMtkv+wdCo0NBtGe4ik6pvwSXsZ+RThPL8Rf6bwpu6UljvTsfjQFFuNc/JLx9t44
sCVzorskyvLg+pbeyeW+cABsFn+pu6Q0qLYcx2wbm3zb5vLiezAm2I5vwSP7kGcidbD4KU/1fxuh
hAKYZj7zK264C9lr6aIM5iLkOQKkCT3cT81hGlF8YmXV+V5+pnszBCyE/zEekDk4VX4cPb0tgR0W
9Pl+ursCJyIuViE+eiiYNHtUm9/6icjhuy+6SeqO0OfbNaDy239bCAljhirkOgaefV95Xyex7gT9
lLPCqz5o/NUOSIe30OItanzOxQ6vHSk1c1b3Sp7BOVMYzEMqdwh8agQlDpSHQUuzX8Q07Qb7kqlU
KGTzVhBrwS54xdlpBzH8HmRAehVX45NLygbV5fHnCo8fopF9jmlDaAiHNlfrSjoXlTey2gJa1AiT
m3y789NqMhrRui4mdo2Sks4b5Hens6AjhhPILYuWJ26QXquGMvGXHQ6AU6jbwPBvqFuiZQ5U6Dm1
zGPFBwYI0zYa6pDuXKQeQhgzQRj79DYmt4yzmDEsXDSsPLzU0xCw452Wzn84RzBJpT7TAHnjHx0N
da+zhwtBLAZ/lF/YIoF18qTmeGJE8TL+fy7MXACtJTjpcGBOXpJ62CyC+V6Udw3evaCL1pVxbavn
0sLYVvUgFP7W65bbC7s8UtslvE3hdGH1CHm/QIOjymDdISpd0BdJb8hAv2mByttbK+8ZyFXl3gPp
gaeGsr3SeTvd8GVIEUM59ODQ2TtWW/oeTQ7vRyNB1BA/lm5OISJDx0wEQmjy/Qf4oTRPj51F62bk
6IA+yNNgulNlkXIdZ3HccceaFerorP5BPnnBnXDw5FDjHXlB7vruhugwh2tzsIVgBDPrw8IopPbh
s1EiMMkT4g27PH2dU3OOY2AlNruP9aWilQTcJrVkpFjH8Y96Hb8gEO6EBkoVsx3/7EG+SIKJ7EML
yOzTwlhHIRAi3zqE08Ukg+dyDJsoiFxVauXY6iRSylFRSJDMgJPgkBZWwQ+klfnu6Hgua8qvjd4z
OQ1jp3/8tyhhZmFNkKkdh7PppUgjtJUyYaoAKoUVir7BEN3Mz5peLevw1yRp8ohmgoo93Sp5J2FG
8wNyqwS3sWSs3sDiPG+nFtNYDxCNnuw4vgS2H4kAUMLzL+BUnO8TiUOMLU361l5TTNMaYCZASkrE
GoBsOrYbiXcKvv1rlhp9TcBC6sowMLHton2ZC/zuP6kQboBN2TXyy2rPlYCCKW9RYehDNOCCfirC
/ohh9wxY/3Dl+usAsJ256ogLM0lM3HwMEvmAlygibPgViyOBjRyaOp7ceaNrqyK64zf/883sM05B
r2YFh6f3SpJncTrRew/G1sSimbiwJ1c2PO2O4ZfTJjh/9xxnvidrak5V5zgi6qWN5yHaaOXxtaiA
zfsbJW7GDccePquhxjsagq9ZT803jiHlj3WUE9f6Es2Dy4uOxjEKkqYi5rAIzJzDF19GU1XKHGJO
R/Ur8o1pFn8AiSm6/5f/5G9kmt6S+wCZdlzyCgBQQ+deMyp345W/nviP/sWqejeXIF2NqQBrWeyV
zisvdzobGS8YP5NAz4hplj30LgTuUOQbQB0GjbvKQHFrjAMrc872X5jhJxd6979u9UyulkFM2g6q
D4/4VJZCyozq/cmBun3PJIvXD8tiybRS3oF8WEEjvdFljMGy/e5iLf6ez46A0gkk2Ojj72CEjLYW
EsYB4TN8w8LPJZpnX9q+m8pU1mM88wvtIRlIzjtlCnkTAw51PwsSCIja8lH1+v555qostGy/sdod
xjLfnUimNYlXrtcqqSkUfkjMGPOXRxM0kizWnuSFUfkjb3Sogk15eLweIAt/h3Jo5wV/9X41MatH
iP9Wvxq/H4/tLtbro11+ohQ2toI44qxx0HXKADiFKowH5epbPUo1QGkwRrh0y+DXqNDl2NCPBwdh
fFRMM4It7epYV+OWNLV3SGYoElqJITjOD/SEykyxFRdWuwdhF1+Fs1IKe74EopATeZ6LSJViPWS2
nLB8SfdKdG0lPWP3mKuOg+AvSNDziepX+C//4lRkWA+PHYkoiSxL9CJDai2ZlmaU2RRRGiYtRwgs
hocrndA92dTCKXPrTep0YkkRzPjOlhQKdabnbJym4+ddZVFWB34jSHSkWqD2IU9Hdv+fSYi25L9X
lOSlgCfavr8sTBef8yuKccZFcjDRF1q46ZnoEHtf2cvHQm3PqTxStPzKntHumvOJ1ef1i0PnIQpo
sNYJkeVs/JmVHEO6VlY8RFUJE2F9M01ARsch8R32rSkwpObhtwPCVldtJe1EEV1PLfZWQlbuR6A2
ge3VEekYn3tzR8YcenQmjG2L2JcOw+qrs/YQROg2YtPJOI3GC5EmIjdO+006k6od5GeENPFhYnct
Bdq4YgNXo891LSxtOvkkWmWSCrjXfmlKcGCLYIW33M7R3YzXVBwDAQLwE3aJhsgIgYSl7ASkDtj1
T5v1sos5UC2qsqVHGrfc0qbwIJW94qykUR0qcVUQNRvktbTfPdOIoDxL/F8M13CVSiO6cjZwlblY
3jmNQ2JEZ7YBBePdS4UgzLuonJNNZSsQg9S7Jo4bHWzf/GWX1rlbMdiwVhRYthYzEDwktC7gfgOm
taYU8PMkWFU8wicNTLQEdNQLjcz4Szz/RF5ZOeW3RBcuBJeuVC7tOmbS8RtWwD9wv1gBh94L7Ppr
mA2IypDYw9zARdkWl17EIVC5iff/QbZtl8TmygzXcy38Dj+N5kAPYumR24o/SgIk6VwDlJVzcZSW
5v4tkmvENh8umLK1TCb6Z1+TqUjqiljwLEL4EF7aISPiTJpk5n8/rOmz+p+FFxfjvH4Bt1kFPEdl
AN2XQJMb4r1f4ni6GeUNJO9CWVoxxGyT3BQjmgY0lE8X5OZOUZd1juUjh3ggH1S0hK7O+NhbRuaF
rgQ6SunDHL4AbDWp59WJuOIz0AjWqem9UepGmV17jnC8ltNhGP/R7rlWZNRrHyU3Du2wAvUhI6GW
HD2n2Suyo2LrcmiJGamnPhzlpnxhzPxbr2mOL+uzXw+yKzu9O2brAy7rrSLCoQIxW5ZWOJfMYgvB
JrjSjGkiKhF+dt0GBiYMrWNFQViz5+E3pKSvdYekfCYrL2Zc735k/V72z+V09Vk3ik2XYaBHbxhm
45aTxJsxlTJqqi9VzgGuFYTaEJwyAetNabAL/VgoWJvAbvrb7H1WZycMGjL5vO3v6AQnMOEW/OG0
T5fRTGuN4jkH8xA/BxIPAoNwh77os0Prcrh8s8zDJ+OyYNR/x6MyXa5Rc/nAiy6i+o6/uIJnPENa
EunG4auzt3fJeFasvHnw8sgwvnqlR3DW3S6Rf3lNp2BpihCFH4/Ski3FecC7i9aNDd4x89bmMRmf
HAyK3ro7TtC9VJkmSuG/poVGphEh6ZbhmT8MYH2fECY6fv0WxAJy6xrVhVOlc9N2ptNchad6Urfe
OsCPVk+gz3d/baQbkMyor2pB533DKM47u5P1Ri9IOOWZmsessrxtbJR/dTgW0Yt+SETXnuUB2L/o
EeA+VrJePlQSznqeHYEzL6Pyeh3q1gLklOvujvgH326kXyzsba0DuRZRoDkT5gMeMVeppZJgLfxg
k80upvF6ySB5HUqp59/x2Kl8sgPGaaemuip03qNePOs0tP58i3ldaLpzPQOcGSKjEbA7ADFAuJGc
561HH80BQZ+9l8vYMmSjRZPUF2pFxoaOXTjCQbUXj8v0CnhLF5stvEppx3EloSCnfaUC9I5N7+fA
8DqcR/olz7nCNOV5ICOLHMJ6NYyxDyVjZtKls1Wby1nLvG32tLalKkZ/rmozwijTLXoU4M6sc9Zo
uv0wDugKxwzeq1Pj41h77b4GA2s03lNQgPG2Xf81VKtisr1NZTOaAWB+LMDYZBjL8vAa2/28IRqg
rrHoUTlgH+zTgek/jK/mnvRwq05GhyDLR1VgdfQIJIgLd+jZiwt5CFRjbiQyi3UfvT7sKZj76bye
snAW8wkPnQjI5lh0AdRVB40titR5wu02I+tC7ln9wtiPyeXAdl8l6YIjacvvtwZymD3p6KLlJaCV
olI5yJkJrQi9ZdDcVenRNL8mGNsSyDULaxmJbvL8grh09as88XK1d7CWgYj7ZfK37q0DgYMx7JWR
pSieQAYTsCaLfFsW2GtQ6snuMXv+bGfX6Q5+GMMyVPnj7f4UliLCeYEA7NzdS3UO7LThMiy1KXKO
MfDlSOE/Xe65fHm3VOVgD28KhAA7UMeBofrTaXmC9ZAvXy6IupvWgthcf64pLr7impmVkA12YsPn
Hzm1ywVZ0Uh7I4j5Bjfhub5qzMV5ZQRFOI+7cO5i1hzgdEPmD1Y5ROAZxuIJcy3spbw9SDUbLIdo
2tczsjvyZ7C4X0hNP5r5q34NCjj5fQSQMpnjG+6wo8yE2i0FY+gujg8uaRLxF9FXZQgbvPGUZ6YO
O1XDRORi37xyXaGLUaIs1P9PDQ1FuiDsq6+vzAFHJs1QJmMGm6p0YbdJDHo7Q6rs/aelAMt+gu5d
MZomTAL9ZiOdwGOSz1SuHiz4Ha6TQq0tSf6nrZqbSb5obHVSgcWtx2LE1M7xXG1M10BmfgQIDWa7
Pn6WrymeG1HuGh3C8rW+iVN3Sm4K7dR6Ugnim/KRhfpMH7HLHRtPCM0q+sZE3pkv9o3URRVvD95m
hrW/Ksdarunl9ut+Kmj5iMujUk7IJLv9VJN11EjJQv4GCwexrc1mY7IIxN3SVoAffXD4GbaZVIcX
ZDE1UsQqP6e9QgLM/uxcw8VPtw3U3fwp51wwdFkBrQKfexUOLnEj+2YCwTnqtEapsm8wVV0zhEy/
IMQehtSLy9zDpZagYz5+OAzo8IIQE4pUluA4bZt+xzAwD/MgBRi93zwDIuUfff0oTPsMbqmNh0GH
8d0O2RxzuJhQMaJKd09rONcAZDhVZQy3r2IRJEC+6P7tkyi8+vwYoMFbPhr1aygDH1vDnccBKSxX
IkmXEwojY/uPb8aqzpyu9xWTVfgadnt6LQ/uE2/1jN31e1sGcLYQUMZOebJ2rnbDoYG3rYUHT5fP
YjjxGeV1LYGiBobMgo3XrQ4v2o0zJwKjB9X8AwQu3PkGmbmbEC/u91QM5Bn6HyQJTv/qTEYsEDzb
h/GfiCPimkiPLG//tvzoIvuAChHHAnLJ7zESNfoA5MrvHsOnN2AqyL5+XsJyth3o66fSQCl8j+jB
J6B01m3+DoBAONdvyrA+p4EMJBHAVzo1ZuKqFbpWzrdBEu/1NCXphgRQw10nF5LhCXUammtJ3QV9
8pC+vPouOx1V+cC+hV8/4HVR3p+QJ00/anND9D5QY/iHoIiuQFDvq8gTvWTAiPd03ecQv7ar+/6T
2Q99GHyG80gj+jOHq23+u+3OuokOgseMWg+MpypgV/MyGluDjOIQIKi/Yz3B99caN8Y9UatI4rwQ
51w12DP0yxENf+CJc0aWjHFfo0y/ZJf36vqelIWuq89XG6v+CGLW3S6HAW5bpNqpH3JjptinsmjR
Katwxyjm0sn4FGHHFQQw4loBPZe+qt/PC849tCYqAxNLldq4MNaDxMsa3P0hXLp70EDNAz9Cs5RP
+S8HgsiqfTL/VXCrMt0xvloYZspE7dY5Ts+RX9cTjnQGSMps3etzeqqQdpwq986W4LbvlB1CXxiy
RJKJPBtuzcs59+VK7PLsTT9duNo1BKM0E3WGptBtjV0WfgtUliwaCYjkFDE9XCq3XMqZsNT0BkYu
dI8QtKo19E3UF7Ti78cRNHqWIVcLgTFfXNiUH08vA20vzzRhrAMl1JwFW/1y8TiXr067lOVEXuCu
IU/pIiBwsxVTYCWcSJQfOIZv66aC2iJ6y8cq3J9z6rWZobxiH7HnOfD/A0UYOhDbcrgog67xe9H/
X9FuohS5qmb78Pk4BriYULPXXb7/EvtErO7VWYLDf3UbEjx30P81Eq5Qe7H/QYYmR/U4WYehIB6f
8r6v9NGpVhWNwRCwgJ6/ppznRSoRF2R7AEwP/iSO9QtMF+SBP/KYlxX0PUkF5h5jkCCsd1UxH4wa
/fbHkRfDctCXnprLbZ5iItQjQoGbB1gAL1f+UvAxR4WAOumbsNtJ5TVqquw9RD2qQWF22PcLPF89
YShCMwsBe72W3rC6oFJbniWex7oxvM62nVfAe0F1FuVwXrXIhxeyy2utvxBkvX3pM3XVoD+z7P5r
jsKiSj7hQZdxv1CkMOZ+yC/CV/v1jq032ZBQzX2MvR6iy3rVy3L4Hqa+x59Z3XNG3PHzfnWU+oFT
dRHCJ3NbZOVWCGz46fKTrLKZLLoMeVTEwcA76XV60VFcQLr1QXKYN6p9Ov35Joa/ujHRkhKwbmoT
JibfxJkB11wwFXzJRlS/P28V43chs7IHkRKOJ9SHkm6vgwJvTLkM2Uj0QIDG0TrPSKnpUwkVFXE0
AbWpZOZG6Y8H3jqMXFNQ+VdyZ6od/XCxmF7PDVBoPdMA8say/Bc/MEObsS2t8UIyIpLnOEELtxBw
gC/jGXDdiIhZLFN++yquOrlgZpobFmIxY/fWFT1/oeJiVUbhHD9TYj6BNbOffNGcTJHY7HlpZJib
NFXPpLAM4MDwdiF4ppdt05hPxzEyRUAT3CXDEsuLMu41AamIme2J9Qqp5HzohHZ5/GSVfHDzHqOS
59Gc9iREuz0scR8t6PhzLdWlnKMKrcbO/dUmw/Yu4qSpElpE5jo/LJYYV//jV74gCS2R9/vp2980
KiI/49Q/6/ZZiZQpuU6sY8EkjvNkvfLmLJyYXFuIZ+VgSvub6YmYFbC7988VJ7+jmYLmKUUIIV7j
sFAw68blNzcDYlZdjRene8n7QlvPET0w6TH2f3gB8YxxBrXmLQCYHwMXnPRyxWBtn1grsvJHFnXe
HYGnvaET4algq4KZ7uvSJVJM2Xunkn9+6LZvbXxCkhVsikxyaL5e1JyzyPe8gjLxhF7XiNAjhqvw
iVLZBY6X8NsQ2rxXLr1SGYbPzCC0C0qR8Ni0gcEZY552IJtK7/CzUvdtw0jJnRy/Hrp9aCjaJIvo
WlwJzTjQbREXcnRdCpDlv15KfjPXqVtMncnwyzyWnpu3On4VJRwbD8Vx9eRwaVH83VF7N1W4qhYq
MjLm34hlRTyj15HwB/vd5zmg/5LkMKSWXSalqYHRUZaoIOk3mzblyOd1ZwIl+foBdfkK36JXzTfk
Vc3kz6cmgAUyJX1xJJqcWPHgmpJWANjm6GHH/lSRlpWCo5cFunuh1H+tDN6MipiykvsyVo6MZiqF
K+/faK4MCaE1ycf7PKrGoo566gJ6IEzI8ohgR6dtFjC7vHBALOkU9kHFga0qA/qmV+fc59oeA8XC
IDS7VtVu8Mxdy5HSEmVM7gN93Na1gqRFFy3OiThhSp5ZKRBHia5i9qhORc+iDZSIP4rGTgGNHOHk
zCFLgRW5s8u/CbbBf7LcRAEcNtfC7X9v9ZYaKtM6EnNa3XUywojsXZWGNVeXvIP1hC7n1hzRVazQ
YON50s92WbTV1zZcJLSimgYtLE5Y1DFu9YmEF416epfKeaazH5PZspaTul32SU6ehV83Cx2V1WeZ
p3vs+ZSh8PoGqXVM+OPQqOgL0YyO/7be+OEcSQrhosJUFN1yf+bUTCraV5xN8HWf2b71FQIOWSGt
uZwWXgNrVyvCJbdf8098xnsw1DU2tPCpeC8JzFf+9txTb0YULkd+CQsUWj/vrKnsd/3g/25r/gT6
ngSCsSqrdqCoxodWtyjJWgd17a2/nr3dae1PztJdpVBhbWR4l0626Q0Bwiav3YfvAduLJpoXd8dU
PIu96CrUgQToKSJtIJnf9caWTsSEi7zyrUoyG7bjPURoCtkAaO7lVA9teMgXATZof9jyPPYv9BZK
mlDIyJQxxUSuOE/3c7bx5dNeb4O3I83fT/gexXg0w8RtlOGta6L5mKu4VNbqzVf5iMLYIsl9zAoc
fFSCvfZLyuhSZH3NhglRlysFnbPMQbyvttw6aK/WN4c/NhwtAgg1WCQ0DrBRNLcRre4ig+5ZZ82t
lU4iArOKFa4+AdJF3dIKSTKNcRzaAwiaEq5pACqPGKcM/vlGqx6PMaVsBycQtylVXHWlFkDlGXpa
/hFIMCtf3hSjISOjYF9QTR67Zr/GNcT+UVObEJxmOrZ2AeTfrLmMcFtFYssyyOdrPv6Yu1j/Q2S2
fT39eSX3Efm+sggUbZg9KnNFF71W25H3UxJjV9uhgtlMS8dQ4fW8DxmG5hPT1J8JXhdn1H4T9fjN
Y3Z5zEoH8PVMA1uL5qYy/a8VJkPfuPq3+TnuXkaDuejr9AoJvxeTiUjnkZoOpfSRJ0GTb/muNP6s
AeNmh0yV+1Qwl0jctwCJeEn1Oq0jM0i/P8OgONNowa4gbv6eBSjLkcVjSlwWYfweBSs18cUNxUko
hXB5++tu4G2GhfOBM3FEPU+dWfZXdMuTfGak1zynGtyBaNF6rSF+TdRbB9LlKkSn9w9QrPgmzJOL
1uGXFlCvW4HCqG2DvCZ3PK9OM/0yVDyCbWImhCQZho9JosOGTukSkyYr5/t63prkz0CQ+eJ/jig3
exjIlTNvaSPVMs9Z8//HRglUt3mTXMHRKjvmaD/D+OOqIL00rUfTr+GbobakzvoVc0MqbhtpCu+i
+nCGoLESHS3G8I4M8q8OaWv574tPWoy8aFK+Mp4dprFRa+o687Tjma7K57z6ZaRNhyTf4786PoeH
G0kLAQD3TcP9dULiZyItNab5t95raY+ITv/6XJ2HjS9MDbf8Dutl0yTG3eCUbcQces6K90ewHtTl
74j3isB5Jfmhmjrs54lr5qBS9PZOnqIfaQujtsxSSPbRF3SiLzM3KciphcntCo4pcswKZCKMqnuZ
ERUUeaQvWamZZOnO9rXSHvD8p1EGfSJ0ryMHkQKMlySisd9gnH/H0ClI6E0CMA/vDSFYLHyBaNqd
XYgaLXUmllcQ9+TuYMDLYzgCqvhPttd1v4TE+O3LfesT+oGcw2AJmipBIfZqG9tf2bXzP0Ru/HJG
F2UbdHHi6qmUjC+tPtrmPXVb9cDva3sJogbzxGBLcRdGDuxuDz5DtmZ0+HCmi4WluiW4+C2ZXIwB
UppsETgwmVQ4t1NsxmLMveZW7Pi+Gq70TB+GBoGOauGXfEXStzeeWJJb0PWi7ZltX76SKLrZPblL
SoXuLzk3cXcfVc0HCnzLX7E3eKN2jjvBLvnyEmoKYyAomiaJrpxi3jnjc+hiJm+f7Yx+bVdJ9cl6
usarnVPipD+3Vh9VpsH6NAz7y1b+J0CKwFHYYYPvVW9XjqYeV764AxmhzZdvyr7MwJuqGfpCvrBz
bi8MUUbzDgjMP5u9+y0W21ul14bmGxzq9q/GCBDaykfg4aQNFJbLI631CAdlDXpCdl2VH957RTdi
I5XaiyshohW0JytDGQ1LoS1XwQ1UyTQh7/VEWKs08b+oxQfaSkzqBha1u7jTGxcnTTHQL6MmN1e2
1Eqf2YeLiLNXLfRkcW5EIN9tsTQekDQdd4qU6CvguZfAuLy2/D4cnYSOFu9K1DvTehtKhe86zm/N
LplmrG6az5zOy61IhLf2fWdNZ/+moyIG+jrmeWsTjp3EojAwq8oCrLeECHsOV3NbUMT9n0vrz8JS
V5LGg7LUT+47uoitidBWXY8sXw19tUNzItSNUk+d8uotdQ1eR5ArkA2zvNxkJQiACh63K6s9pr1E
rcn0SQdfotlK2x4endGXARAorNrSmeq394TIGTvnYND7Cwl0nUEfW/AP/jZH1BVXp/bWiNzHSR8e
Iocm7k5QulTL5uBhzmgMan7YuYjSlIlLx4xXq5oM/+tzhhgz0JYqCzow0Cxml/CJ4aqIzTm2Wred
iu2BuC+0kAuvMYSAtKAfBC+G5D/kCvSG0qZD8gtPcSdneWfTxciSFnXZiLvI7tJfOfzNMcXqhZa0
SXZV8aEjQwiczIy2G9Woq7YxY239239qiaJYNnDHoJDg8pMR9VAnxnej6Z4Cwwxvy8Oerpiwk/YH
x4fQMlUYNus8O2pZ5fl5cqed5zZMecOrsoh1r3qkSVYSYQrcMnVHKyMSPRO8DVkt9I3l1bHc2wOE
cELuAOfhxjHTyahCblJpouqsvXbfndm0o05EiXWdlqRBrX367h1kYXzT1jnR39aKYGpWc1N8NRRS
DgJs4VUSje4bDApFPI5cZyx+hD22YoMnV2zMwj7ypUSnwYqHLFVKZqx981CPGQCzgnRgVL29a489
hVFjLskfjbscUkn//q03BESgs4vUlpJNW0+nRaDlSekQVs+VA/k8qjXcz3K1U3k+vcSHBDmvtS0F
3kUgnnylsQ//PohwJplwoI39ZkqTT/K982263Kt0nmNoic+cwlHPdw2p6wJth+sgQTVo/gbAlSWn
V/yLdVEbyf4miE3qUbYZw5FrSL45WEehFbGz80yqKaZLOo52kHoZw//gqg/0P/VdTLJa1aStyw+n
BJepcfG9a+FJgyO2pBXWXFdmtBNtyGQSYUG96sTJW+uXbtxCqtYFLOK5DRqjIika04KUeL/4lPqm
9+v/5gNmnYQZw5SC+t+4F5NYzqiwJks5wi5uPckEHmkrZhGzJbnYVt/35+FmJuNi+uu9MboT/3lV
bCN0ldNkWyX/D4hPFxyXLN20IWZ8Y+bDHs63a0pY75pROfyEgleF0B2sWWfeWEkTSRq9mXFrdQmD
Oqn0qFZH3JWPcjsK69jqpmdHTY3mapXAQZDlppX8HBshhoIZexHALoMAng7khN+9tbboKQOR7BkH
taejhXnW3ZkC1CEra9BFTrdIvnQ4ixCPpBs/iVHJwF0iyXCn9RXSvRnEyd38CU3GFJ7GzdAjSAoB
9nCstJLT6/4LRTZWdEaF+1BfPfVQHhsApZEMs/zOAo15aZ3aJZAGp/KKyhBLAlitjPKWUaqBm/6j
Sk/TToHPlU0r+i4yGLX7xmZlthfulrbRJ4psKjloUy+GJpDW529CPmVozs5BzvLrkQKSgRRQaUJf
ovyjxLJznEd0nOevlzcGEWiC/zlVMu9qvGovObciOBz80E2qHnpcRWGeu3GVMIS/CIl0V/48wK+d
wpnUHMOz6PbjV8Wo3N24C0CJjTLaXlEs9oqbZZaQSe7RYA6BHM9ZxTwxbYRkERpMfGU6rtGizYS2
tb2Pe2LesiqmDhcfqQq3Tx3x1Iw70+vqAULH0djWuA8yB8cneJpp+h0KX5r9rQrEMK9wXyq81Lom
aHNhQ+QVu4aOCvyc9ppemStUzNtnBof+o/btR/WSrRqZC5hH9Xxq9gPVpyo0685XqN+bPe5MByVk
/IyusVoY6MZyKsSOlEHVH7UV254lINCMa/s+Jb8xsWTcPHZGkSUzo3j1q/uliF7iPA0cc+fSdlWQ
A9RMaX5Rl6DpNwCp06g52PSdZqS2tPBZ7w+g7zQXzYRYuI+9IiarfzkMK6/CUVS3welXT+UNM8iW
bv2MIZocUXaJi9jTv94vE70OthJoeFiYAMH5i8tTJxrLG4Z6PniQ0cyOLCb/IarIbGkmVUkwd0Hv
Avvl/JplcHKj9hyJeUbl0y5Cd+6Nh5OhoL5d+43ErPZlij3lnDvJRP+Ovwi67I+5V5MFGMXU2V+s
pZEUW7qFdIlQBay0K0kmUl0dhxiuuCCFXEslI5SqRqTPFQnJzjSwHny7gUojHW90nf0eGNMKD5Dp
R1xWdrXmW4Ct/iHRT4jZVToGIoSYRJ+ONpY1kQIMvZz0ikifqhKRxWjQHS9SuY9VAEwvGgIDjE8O
hyCOwjm6aUpIqEymWxCNRM8LcaQS2sXNDix2nxaE7zKgnR2vVYvuvaROSxg3ZY4uLHVYETp6ANRk
YJCtRybAjC16Lup89POpTyE/S4WeK+lAeXcU17bj1ygklzPXK+uG+p/2mCNeslWfqygzXfF/PDDx
taRSdcNq6pDv2Exy05pChVj5ZAtVCDTCYY7ciHJNLQ89KIUnwCJvxXuJm0W64bWl7jYqPdhImUsR
CQHy0b0UHR7iOZUPlTksJZqbxhbrJJlnlZ69gWuSj4Q9n+4I0QZ0ItmEyhmIFcEref6gze++RCxt
YxLyaiMkfMpXJgSg+9QJba047GkL1eMnSSFlkNFUb3HYauBOBHqRPkILScEUer41QY5frWf+oI+A
L2ueg5ijiNZkx3UVuRhJ45twWjkyF5NaJWlheDvkL8lQpfc4ildr/7zQ27l70aUAGLj95c98dBla
Dj6VOJyo61MylAXkYKtImpy2Lo7HB735UDEpYK5h0H9VFl04ifLFzjZfhH1oc8+9fYKPpZaH4U4Z
atuyxN3YiKQjgDGAySmsuEuPoqH4B3cvRkys81sXUMJ2t/a4tVcoKcO3ogZoLnqA1VpXnGCn6ryI
SDj6tF0DWNbPtAb05PmUak48iswQ1e2+rca3/OQ9NAUCgOsqp0/hwAu3ZpioxUIIZZbW4WE5kn9o
YBW+cvDfWcP7tRb7tgwSgbw/Icc7imGLkLQOMKf4OMJLbTKXfFcMn+q5c/iN8q3teBlDGTaPdxbs
w8SSidXVNHCL+c7r2o4J2ZFHl/oy6m7ipyieZivf41AQAwp2McwN+DG7C3CXin68zmEn5FNXlcnw
JfkFy5TGCAArkm9nShUoqRFUZGPfsQfr2EmB3SkV/xEmwhaiOfVKCi6dEu9uP5nu5+5U/Mwlj87M
szqcMXPRtxR1Fjy8hZe7fPrRpYcQmb/zXUWvI/hGIBk0QYf1TO7Tc2ysDGU1XNy+SBbQYsHT/aAd
nvGijgv4sxNvNXyrgJN0bTgzGxSxm20esPpJ6LQCnrEuj5lD5JGkAF7taAWEELVH40yLw6LdKLmo
Du/KJLh7jFqzyFM3RBR4GsaMUOn3CKpa4ktvlDmsW0Ln/l/G9gBX7BBi9mS6aX9WH9q16A7dSrex
HZQDumXFumWxY7gkw9g32XG08OAJT99U1xKVQiveW0/Detm1U3g7U77TLpislwetepYgSWOkKhD/
XpLZCiymT5OCz1Incc1AtQ4M8HEdPRhAd2gPU/aRoo4JMJu1GuMKwCAkLJ5/hCOcGwf39rOJP9Bv
fpZUs5XnYJmT+sUNdq0STyj5B0kJIVRX+PB/wbIPWvgeETc0HlcpllHdXZ7Ik0Oe1or/8DzryWTR
ZOXbR7rip5L3wY5bjmw2J8W+IqNOmCGHssG1/EGStcHJaCBQ/+a48Z007Ls/BvjkgLR7n8rowjfa
b3nADd7jfc+M0T4YAlrSDwsUVRjrMSHLQ+E7Gt4z/kcxgC72YAO/UM1ZCJS0P7v6lV7cicHsUZBK
FezuVpdsBsmmufHcOlkuy+icbmvZg94l5mWR4wbaqIo4/U3oFCl0qQAcGG5N1rG+1L0yr83pKAQZ
esIq8Cg0PHtup0woq5INRwI673W/omFF11KJVJRJsxiarnGaNddbl9EjOAh0pK/s05Z8CYAahtHj
ZM9GBKnxX6mgj6+JBrntDKeuKTmB7NihioxivkW5cp3Ao3HhLsufEdZ8KKwbTpVf+RZIYJyEzpDJ
iBIyi85GG+QxV7LkmXOk+noORk6d0g47BLY65MM5t0JfgHvdgIp16NQvLndCClJLNSJMAakEUPQG
nOkJiblQUtA77Wxdx1ziFjUABrRDhb0PeFKqxVW8nS2X99lIPjY8MogVtuGZ7b7Ua+EgCbqsOtcq
NiHeS8aB9cE//RuWGWkb6RUujY3q0t0OXipJjmPgAygsgAwB6dI7B631f4/i4AIMl3Jsl0MsuC4m
V2HvCj/QsxKTUxNhsC3cR0pOVX6epUsIHLH7j5eMvC423fqVuEKzADxCcEtiNQ1YIAcZdNkkVH7b
TUq1TJ3pOOSQR68pwSaf5oB2qs/wEqI+OqxLuDsbPcn72GQC5wucJoxFYnagklw/zCW/kq2jJRGo
0pOKtVLC2nCTMM9jUy9rYOFbJXuXr8omfzWCAfVvPZxOlEjLOb6svN8ym9pIJcqEaj8qtxim5arL
b86YRw4AYSD4DFFMchQdUwU5fQVv+e7uNUPvPt41R7ENpUdQTQyRVUtdJ4sIuOBEzfhOuOt8IgTp
VmKD+/oner0dx8QfJzOubr596OqPhXYr5KzgarLzeQ8wRfU2wT5u+SsFAcb5dLy1vGXBNrgwWTSD
bXqeVbRrvhdk3kLQtJj7XQddjz4ThcBwJQUFWj29gAOCuO/EfISOOkY0+hzKXI1KX+FZt9vu1P1r
noqq8gA6Czool3lja9ivsJSZ3KxLFApPgDFS5ETCkySHrOFAcYUCpNg6I3yWk0BvG+uHI2RsfizF
ViYppgkRZcI36OiNJzpYR9YZ9Y8Uucr5JlKoR/jdhGMRoVhyxsegvoHgG+xHeQp64ABps1SjMsiX
jip1e43cyCZWoFcbJ4HhbcoAqhG6OmlhrzWRe4ZTBOeEWsx43vGEPDDoeVY/nvWcOTbmTlWE/iVj
BnoKDhUx2U3K/IACdTc/gvCEnUl0FIDeT3HiB1tjiWWPK+ttewZG4cgKtGDy1uRv8CA2q0SrdvIO
mv118qxUFgCDyvgD1Aif1BkzkH8uO0Vy34bo2MR11SIpUgul4EpmuiE6xrqFqNPPcEwL+NTqWmiw
uRv6lU/XrEh5reLiRKKseHyAHJ9snGE2Zu4rli+7G9lw87TAA2naHERC6YGM9LxdItkiJkQM43H9
jkjY23jiTF3GR1nsbaxQS6WHO1CwSRxnA2qMrF8xdp08D77L9LEef96BgmOXkfOe5kCKn4KF3OCB
yGFIm4Zt4U2iZWAA3TS0kqmbIvejtXb+9wEGQ+Tn+ua/aquxKQltyy0n26Ph/juXgNornPFWAabf
vRvB0Ngfv6nrw+RiUT0vk/ISvgEQX6RzlfEOr4wnIHoTjREhkrPiOnSKf0jlHuNdgIgRIKUtCTJX
S3cR8avcTacKhnNqdqIL+KCPIdMyroAea7WTK9aX3FrT9TVklkADxWdr0esyInNlUMKihp3YB8t9
WJA/0rpkoYP6NeYo7+GGSO6c3a54+mKJSG2VHvAtdISWQp620kqxa9lZm7aWdLfyqKOFiXJpuOGB
aGqA1SrP0WZ4DKwdTr9TT1nuPuFQaVA+8PE5iz7UrawuJUwXq579Dn73qIaqeeadSuh1jIzteKTn
QxAf4Lr0RA6SN8fxTnFP7v1mhX3HHH9UAVD7/cI5m6JhxF7BY/8qp16cPCU8PN3nBV8FiZXrC2sM
i7R/NSwNLZ1ugeLjlksuEj2fv9zNdf02u3lJnjzTKc3aDgVmHwi27ddzXbV+QD0syIm4gM9alhnm
xxiBD/D/AFgD1IdsrovXawrYst4fF36Nk+tDhBRovaYwNb+DdtY3h6P7iT7DB0B6d7uqencnSPcF
fqaWNbgZAwnUF9epJpezkC139/REAsUmL6YTgZVVN5NZ5PKZM8wPfJCnrKJi/vZgpsZxzVsst2Jr
6ccJgUj7XaRo8w0NFFXwXDAQ7INenaXKz8pd2Yo9+0WPMyBWXxqbyILso65jeijju4CTKGl/QtNe
xaqRcJBKkzL+i5CL+8VPDLRnroPZ2VYD8xIAufRZkaghn+lyjhHa4sL28m+qvQYNcTN6y7eqWKih
DP4g5cNAibG7xzd4WRQaLY7IEDkBmlCH0SBhnc+u8GqnxQZCbbMkMdZmnUJDxqHx/GDOH4023lyz
TqYUyoQfKhI7yLAhxfWt6maAcGynkgmMrakvhls5cwPXT+k0iMCvHI9B1NJaoCZSw5PzssEJiYIi
IPLFJ2mvhisJcjePfQc8/GCJw7O6jZMid4Mgg+7yfrLb++D1y3Ytn5TFyodoTuo6cWiQ/2b3KcCc
dFLIge5LByQBs8qwGW09aFZBKKbMj4rsSQ0F1/ZGP0nNl39eKQAsvZKt/m9B2vWmiS6h3LV6OsIj
5jH5CHP6KKdPuu6C7DiyUuk7t4o6bmlabjXBmi/44DJNXttUR72FbEoRX/awDczA7lB6pJoxD5ka
DQ9llYArtpRO4mBujq8n6+6zwGr56LZuMyWV4Ox9FbJph0rBI/Zuqm7/mRsjHqenzx/4dZ4xyHM/
lNYwbJRzZVgo+bSR9SmYjfMINS7Dzr7EGUiEHw491f8qf0a0ScOlxDaHanJOUX/8LIlrklf5Mizg
ggnDbE9PfSL56A6luQAnw/qc85+wKY/pNchsKjiHbUoi3hsRLD3WKK1fGyvKZYhJ9t66S+RuhEs+
U+4yoHls7DAy28+BA4rFXaKz0cFybs3HmsFHdQhWJTeFn+ICac3KSfyHlpfkyn0SruNJR5LnJ0j7
zYdFILBH9nEe7n6m6To3hmSN6hqHwMJ8fNOqg3PHPHJfpvbjkteGqhplcWAAzn7kxmOpwbpbhmlf
IBmwXNMkgLe8Qgz6+y8TODGYqE0rJf+d3XyAGm3P84gKUpa2LewYcJPOQHGQgNgJuJvBE7BbxMP8
HWUx57H8tIJNY34hZawR5IF5uNxy8aQNw0pQl8kvMQdf/mgnEh0q9xDjn+b8iHEjql1QUB81Tw8/
MUD4EN80O1GFSL15AOcLIZF2lrEkzGL2iZqy8C1uxrx0OH/DfT6wTlkRdvRJXSaDBuOY10PRCuMz
wB4rVVLUeAhGvV02kIFJUSI4JVsLb0FYRoziwnRzYPMLdW/1wAoMDAlGgnrSML6H0QXjsY3Bo2iu
9li86XVB4pewtSZN9ueb2uNKzFuSk+a+uFFA90fKECPRDRal39wz1QIQpDqzB2ZZTidc8X1TboSJ
jDLxI1JFyC0SCEd46PDFBAVmdVQ7zyO+U2APtZAPv+Aljey3f7Mbsu1wdCjh28g0P5mfPP45qQ5v
Iz8Y/QDpCuCMD10nCllhvvFptNqiuG9u9FCLwmXGNfcgdVXCqYZuBP+OrAqgYGtjGg9u1/lgTavJ
phxJ45CAQT73tgyQj8iCxjCcEAVb9XUU6kjzfKQ5pwYypgQGSuA4d1Y+95AQ+/C+F4HWUqOk6Wt7
zyN0uMZnt01bB6EjEUrKQZz/J40MNRUyuIZG5Cr4TVM0RHwcXl0HXn3xPw6qJOC+fULGlTid70XS
QbqxZVHdXcDm6DQ+VCejXmsFkc88Q2jURkyQ3F6G/WGoeNGubdZOLaB9NpHUlr+H+5AvRDkqaWif
57Q8xPcAhTD4Pw26UQIYFhWuGnoV+DLqA0NK6hAwsM4OO3PKa8fghXS4Xg0dcoA8vcaeYHOZlALn
80PQRBdDo0jkj36guSjxYGDs+k/m3IfpZlrr7NhoPVcS+j7JAlDRXcdd71z+UOCAsnICzpRPGKkf
nAUeH/v52h3ZrlJW10AN7bsjeYb6DtfAFNkRn+lmDck7vGDFUCOAOdp0ozGr7zsq1ScBUJnWEciT
jJj1DMByT9pt1rzAoc5fDIG5xMkY5hOyJH2agsIUjkEM4lXPE/V1LugCVHvuHtqN12rTgulT4KVN
0KMjMynikcMYhRVNlHakRC1Vic/CcZdYn5Yt/aS7tiEbLc/lk7waIfaUnAY4yDWsDRfmufloTlvX
02npNL2LpLZEPmbKzj3Z6p2g0pQjIM50JgAApOrL2w3W/L9WAYcWSowqn1pWijuHel6ya0e4o9rO
Kf3ykqTIyWszmVXfRxMSgt66iOZu9curRUVP6NHkf93OcAzniG3gsfhy2JkSx1KWNrbFlpmDXuLh
nLj5dt86O/QLrwOo73by+ROi4t2ZJFxK03AX8yVJY8/aHYGX8zZyyk/MAoEH7293yqJgJS2p0XIm
MHvzHij4e37UDlp97/8b5vLmAn9/RYdKefKCueio4h93Rn8E704VF0YGdf2WDwY2AHldfUHyn5md
pWUsHu+9bWz1zoU5Y0TxVM+6fnkzo4WHOP6Mac9KyUGhFD2ZDOJ9vVxbtO+sfJSyOQ75aCs2obuo
7qMB58CjFRvqPNQQ829Wn9pJhuFG3ygRY9w1rpbfPz1Gt7ltNYQWPDWtfSlUv1BdsI2FrOgAA9JG
MFFI+rEBrhZfIyKT5mpOU5t0yxnmxBvSBxeVNQlUco/0b2MiZBOEiV54VRlmvVessNLJvNVpwLgJ
njyfZazfp0kQmY5c9pPKkwvhA8C9Ey5YXVTzhdNDZUQgUYmSoGHUCClmKMXORjvL7FDbbe1zI0jG
hLcxPuuNXPCwtAaP4pR6xOiOUQPJNAHDjG4c1c03bZvDhcE74Yc9RRt2j4hhisDwAln0AJpAYMGj
c5cxisRgOvCI18YOb9RolUtebxWy/KdecxhneXnYdxQIrBZ7ZjXHgC72vHwXCNS/4PFc8GLQuJcx
cDPBJYqCawRgDUD2h2sQzcVsYr40BGcmiJJFvigaC55PsuQvlrfKGXEorBYRICdkSkFP0URFMaKy
EQ2ZL7Z38nBs6JJSejfNnwPTqNDpAmGTriTv8vXgIVidei7nAmcogV5/v9jPKrkizCSvFXican3i
QWxHDUicVaHIhuO2NC4VmgwfLg5XK3cp2tq8y2oAf7b/JJ6uu4NY20SxHVntnW6w3LsXKhCRDtc8
BMwY0eMJTXCEf1FKBbkaCENLxW4zsQePMRkqxuruKQiuhUYpXTJnogNdLODoPkWCnsM64Kka6s+/
GR4D/dlyWWxOf2vyrF6sxu1cM67mp8sDhI0AXPYGqK+As0qfKtJ+YtE/xO8BtGQ5bqANWOmt2EGQ
PJnPqr03njZH+Uoy8Kff+N2AiiQWhSTKKNT71P4caxP7KOMki+GmxTPMqrnxUhHY2AcDipXECwsy
aSKCcyT4VdOU/zIoz2ii6OPU7c+6zqzN2WjafpsdRKhJtuuTC3H0tFBLvEYFvRxMouFRs69R62x+
GEMhySg9OJy6Ts4twZPAmOcaUpDcJKI+xU0hIZNKB1dW+UMtYlvA05aJWl04VCeAHz0ctEGNtaix
QkEh+lVR1njtlxudtjijTYY0NJG6tPRm8u4IqYGdHW0ek2JMADe4oKglveusGGTn9SBpypTELwZH
rcIki3z58/ufq8359m2+YPQTvWcGmPvSRA7mnHvJGDoAmJWtV/YDW09GDDG2AedesdiWTYBz47zO
tIiVfxhrvaPKRrcYmXhQrNruhAGmvJRTxFVCimWoJ98rYWTyN41aXhKoAE8tCwETkzGRuXYvO0/L
BTMTiOdTYsAm0tVCYffeVxwKkM2enwFRnUndW3KrHkyvqi8CNbEEonboYhI9TGzuM4AIKTtFyDoG
Z8HWj0zXAkisGuFh4csT5BnN4ejkLLoqZ42zXH+dqFavp/iqbqDv3D1sJSCbDnptWTbHydgR5rqG
mQFgcBY69DU9G6V0eE/YP0LCqYlpnVsnQj+zMsBIrLgsm1ZrJUkdHXGn1+w2MNZF/WBEol0FGzIY
o8j01GWwVSO21HvqdQv3sces6Zqsaz+ln1TCevPm0EPcIe92noRfkEJ4i+PYcT0ZXaF3S8Q0uBOI
fkmNqnTYvmfL4VrEF4KlY+T5AXCknR8PpqmQBXUiaNVhGt9g+0eUTFM5cjKpMRKarlmTYrW6rd9z
9N24UMGRNT/LiO3ng3/g42hzqbqNvB4XoxM1yxoaUXiBjTbXgpIIqMPYsmIQyJhstkqWekD+SlKr
j3X5m4CyR6UXAWYacO2x+6oK3fVe9F6AswrdyA0I/18DpJm6WEJcCWIR6DcmarpaZYPPsNzJi7xZ
QTIOXkHFLFZar6s6SAePvPTgrPb2iBOD1MpzD5uNojx/dZPVLQgOu1XOPmuPnvbW6zCl/eajoBg+
T6aeJwt8MSv63+3HqlMFDNtlgM7/qy9LDCKOr4SSb7TcTLS2tVEt9bRJfxqPvns8MPkxsq2UFKag
1zibpjtU6wWsVUPXy32eimOGzbVK6SyhLvvu9VjKymDKz0qwVdOdB+BTSS6lrFIxaXYC4lboGbFX
KRTbhSJYnZgmPVT2vSqIsv6md8cpn5T8NlZVFMba6ZuqY83o2nfAdvD572BPqEw196oK0rc85bDg
hxIegE/56ia2ic8OpkDXwgLImgUumELS7lpNreOnVCc/nflSIMm7vC5oeFanrA5LqRDEKwL1U1et
W8IlxKWVpNI8t4C29NRBssMldFLOhZC/hiGUSgHuldfoEt1S4GR1f0F1tWKHDu8eJ67QzkWm8fuj
brY7QxsG/cb2125KqVGXBbWhCT4K3uogZtfDZI4zaasVRsZxsnay6rqgxvrCITpaYjkMgdqIHczJ
/1OtKnKP6Qv5OTmvJq+0gk0XYtpd8oH//cRr/5Vt/lKpMCzhgtDg05qQVUJfoWy9rE9WEfs+ZgSt
b4Betf/Ru0+XZ40NDi2eKzs93VdOHqk/3Cg+EMVtk3Jo6xgop9rcSzQPn4Qs9WO/xysrLmbJ/hS9
y3DfxJgH5ql7Vkp5BEO1rQNVeMiw4x/JeMdEFUuaA8UX1OPs7+nysEIuMxJZuptCmJBIdmHDmssO
OMSS7CvbhJ+aVcG5TEaE5vJCTE7sh7hp7csAyQ+jgnvl5NCrIjqYlFVmnB0oAtqrEc9HWoTcFLsy
nwdO4ZIBkS1eWEvTmA7D+dlwp4szIieBKNyDgnpnlbL02QrB/yCZudZNeEUdoCQdeG8RkifhcT5B
GJRc72BFxynllgzKt9z+pZ49PW89v7NREQMxSGB+c5uepx0SLKcevoWYCnsmY/N+d9Qd0L4R7iBV
dpkTVsMzdijKxyakxC3i0oNbZz+9SSlIIHCwxwP8rOTZM+TJF8qD0HjWTsOEq4VSPnbk0acTFOHL
2+220MD3cbleLlBBEuaGajTSted2292RO1yVaBUMMhAyGP6azHfjREREK7FIKHOPGcpH8SheB5U8
NIKx8WhEvKSFJY8tMBwZYCFeG6k8AijmZO9aFK6E/5HWtEDIGK+WOlx2+VetvckkuA9vVCfse0CS
XVUFUpO9OOJzNo6OgGwrCD5L6z23GLFCcj6c4HYpwt9j7T6hBIcbGcky9Gf9p4VnywAN6VCR6ShT
Cv6bMErj5LhcF5kr+CFRkPizW/9ZX+Kf2okWm8BVi/mutrty4djZoVqi/+ZiJJFPn7HV9ZYQS/RH
Et1dw7CRNW9vHlYPkLN5DkUPKdgAxy7pMhhc9F1b3DAhI97+zir13zj/vl7K7zgXIQXP6pDmsMIC
vOIBvqORxiy++nCOtkj3DbOxUGzmmmL9YI6LQCVrRw6y7AzYpK+tIkwu4nOuDqAvr+1wPQCwJDqI
FPhaQfPsxEA5ECj3DJNCdYBiXTopZ+0ng/7kymXhf1pRVMa/fFDqpIkR52IjnaOWJZQTlLIGREB8
7ieuJ5+do5250x0Mo/hBQO9gWeOHpK0cm63tY/co3g/2hm5U+YEpXTW4mdRxIhaCQQcPQui/yYaK
Vf2MGTjoy6Ecvki2uSFZuLj3y0aGPYwi7Y/5mkw4Ti5pH+SI6qhU1ALj4NwNf+x2UNY5S8lRd6b2
E2zykgqDgYkXSNCxudAIUD/MMyu2xht4VnKRCpTzH244AJnR+ypPXBivyws0iVkk2WBD+OZKDOd3
I2sSrDuMyybgYIsN1Kx0E2c7pd3Qj4NkxDRTHPfcsnE9HJnIeZqwt3sya03zwximU0+AZvcPKUgt
Dyjjgae3WSt//i9ZLN5ti2tVK25R2UQECjQ/XSXH3m8rkigcc22oWYA0kKOsh3nuEf0muHT/rWJS
vZtg8mKxW+r5SLtQKlwhpKSKKkFSm1vqDxBl6iuM/1joMpPiSjMIZIP/KvCmEWAa171ezl37T4M+
XIloV3PWl1qkjjQUwjxS+cF02DFjwpgAqWUaztCEzPIbpJbsqJ2B6o/dY6HAig3h5IU0JecySv5P
2H+na6u326zC5+RMvl0cB4TBQbKmzZ8DorlYs3pY4ozrERq6qThaQ7lNjw1/pwkOEvqk0IjhbtZQ
9ATspfJhT1NXdnblvOexC2XazldCxQNu7i3hYllbQIaJtAwHDmqT4X43mYCgzf7BkX4EZVqVvaHG
Qm3UYHP1khY10MSEGUFF65JvqvSNcPkKoyoMBfsSRGwKCcGdD6jETnj4224svGrZngvT/0zcN5ac
LXwsw1etYvcDaAZgC5kBKIvVvYBNpVAJY89lPxH12AP3Yn5Tvg0tRybWIOYMRYxLF5EscYSZFCon
iiOc50LrFQUUmg/VKYZP0+JdxLbyTASDNRA6G62smqcipaUsAYmemd9utDVfmPsjSvs8PAWtJTPv
tulaeQBf631Rphf7MM8m0IO0hc3JgWlQLUX3adPcYlsMxjzZtD97T5ra7LkQmcT+I/ayO6YcbVuP
eGfRqpa0zRMouMXjvhuKRr1BX9mlCXtWcLMiALGEw6QyPvghB2/P47HlusPtnj/lsg4jZpvro63G
11wPjFKo/78qhRrONgCV5kXjfdBvvE/nX9mL0CPf9q830/3uSJvwORIuLN8QzGad8XPsqmLZk9vR
6MbG9pm23fhpa5spHSDj/Rk51aHCVy4d82NbTIgnbaLFTS5AqxZOFtOC6AG9LZ+M30CS4Cv5fZ13
hPSR67Ssv9/t33CaiMp2dNy+5/eaidKgx9jsdmLXrqoCAeTDcsbXRGtcbJaupT23bIsVJSqxZ14u
tFSn7lgn+du5T0BAf1RHS0/zYV5CXjRBCG6RVmETeCLhKyJPhSzVLHx5IK3oWsM1MYH9bo6SbqL3
p6R4Q6oMhJoGzGKQxkmnjAXOhAOXbbPS8h1Nse+2kjcoGpnkoa6yn7bFXGk3E2QVxpV49AYdF9fC
Wp10AsHFkuzROPIze1PxVX9foeVikuS6QQzWsnejyHUMmG6gc2XcemnxySHkvuF3BOPW0Qk0uJc+
ofmCjPkxmhPWcaJt3iosA/F2sulAOk9UcGIuwcOFi3qX2cJxhL5p3nAwnuV0zP2EB7xOg9iiYfYx
oQSbSezEQJ7YGvNTbrSJt6e+bJk5xa5Cqkx6UnhE0tZE7BzbIVgHXqq1/MfI2edjxw6hLfLSLb/o
A9rxetWpAQxj9bnfMlmszfdbqIRniibI0bacg58WBXZYspeA081sXU9K67YXw0TJuUyyegaFOYth
4+JGbHQOuS4o/+H5TZoXBVYpW+QhUXydcS8cbUNmozUEDxhnznDIW2RWQF4bvTWx90qynbdMHiSV
evWVIYP/BHRY5JdA4IcKYKrTKQRpsi4ehtmdFuRQWmgwt9/1jGMQG30rjQCFOBiAgYuSkbOQvqd7
vmYOEWxjT1JvVMWu5cpbEZLMjyALr0O111fR0mxn19mO9b1TYYj7Xcu1na2ZEOW9pwuYCnZhQ9Lm
65+208UpKolbbs4A9KI+t9LbAuiWkHzmLwGbbpR9krXHLuPwsN9im/10IsRCyOvkpXjZP0N4MIov
XOc7eGUx/zrckH0vkuXz7VgS4V1BPskXRkNq47mTZ/qF8vIGQd4keU7NdRTf3YhoOElYG7HjFnkE
XRTdxTa6CFIqu8VLyWos7MtOgu2ozxVGJPFhDX3TE3sZgEJx7cLiE+rQRUl5QFLKheRgpOcK4JPG
kfIKOFFdBnAk4+/UjySrRRtA3dfYqCvHz0N0isjqqfdQCzjWvvkQKOlbm3XKRVlj+k9HOUuRQjpV
0+sO2vbwWbu8Cj6DsL4avneirb0jmQ9aCA+YAvip8AyS0acmHr+cWEC/ZmNmVEtHNke6qNLFmHUw
kr520unFmr0LhK2cofjoXMXp2hK8Y6PCmFc7KN6HOr58zITBME28tySHIuJUXTkuqifLzQwHzXzs
DVifWUx0cesNXIlP8n4JzRhC+PEAEM+2VYNxChSDZsxs0XUThIiNDPonNKSOjeceJ9CnOC5SD394
LtuttaYI8rjfx09vjln+5mC4hdzMP8p2eIOEKhGInPS2Q8QH+zy0t96KL3QWDIjMz3EcErb9VLNs
Lm0rL9IAO77Mook8r4VeAHyDh0bGJM0CIt6Nlbmp5aK1YCiPKs3gRaieoXG4tSrEKz0YXSLFN4wz
BDdLi4R/bJsdDopqfZS9mbL9o9eN66cro+SMxQXCcg3QQE+ByiB+2aG7dfkQKPPcUfhwOLxCXiJa
VTlTwLDZd/2ObF7BD/HzEqprFhI+C/QlAzRw62G57Ky1d4r9JZNyqMj+helzpBL1RriCdy3u2q4p
PhT4WRS82i7unqzMP/lp/A8QFZKLcF899NewoO3qF1qL38fDwnvTsS5ZPF1e3lbPn/LppDXy4eoj
MCrrh1n7MxVbvp2XVhwUslpOJ6LJxKIL4tdxY6/5TUN5R4MfWBMjGvEiBqHc7GaFIgOmLF1LyeUd
BEk18pt5NhCRY2ScIaUCLJBr+R1OgtGD1pdCKwvMnHHcBYWyZNeqF2tJGKl7JC+8PsDYHgnZkkNy
sPPRPVE6ijHKqd0xc05FqpJpAl4v5ZpeXvtcNhsGtf8dGzTUb2ib/koPfHE+d1rYrLWvKuklOsF1
7SRmKLz0MRyG42JemQAFeSsCnAh4x2nDSyqSiDQyljaLhqfCOaKBOl6mokd/wfi0rA1DxDuANmuJ
jRdmf5gJUNhOT01YeZWSZT3PlCogT2BgJO/fXTmprqa3gx8i6DuKUgStgkwqYn/o7fhTIzq5pVWQ
xEOckf6uUIqZWvKXhL79slvWbdqUMNJKSS6Rm2tY5H0mPWPLUT5vnIyE/1obyf/g7VlcC2YO+IKw
6/5pr+22Riia+Ll/RAFBhQJXTPI9xbHP74/d9oMgMIRT1as/8qaAuiXnI5YR2ExUbdiMRQgBwrkl
gFKEFD/Tw9ySIrlVcjg5KIuAOhMNM6tlP4btID1cnLvT81VWAZ0VHS4bdkaw4/iLddoKySvkOHVX
IHbUcC3RTnlArNiTdc7kwCHb8VWa6eh1LDHY/nbxlIjm10sjIpzb03oOIisAytIvK4xOqL2EYHBF
LVCip9ZzLZ2Yo5irDBhcXXMuKYTDJC9mO47L5l15ZiSGEeQz8qP3zEw3ZOfcf43TS5eZO8JAFABR
tjJ8guTvV6IhS0hc4B7gVKTzeua3dMY+AY8hJs6lTuYw6ZbIOPneEi3jbsUwtMLQd/+rAHfzitdU
Fj088ox4QoMD/Je5M37WK4hP2gC+gcP9FGCdGRbIWrHlS/tv7dDzuSKPMrVv0aF6/sS0ruBzIow8
Znaa6dQOPTVlwSbwnX0KBlQw5XDRGEZflgUTe7NEltBHhS/LUprza3EOHBxW0DA6ZRB3g+M3Jqic
3BaCQ1BjD286kL89Z1JxI25JMl/ANzuCYBwxDKKYv18nAuIaFR/TRWkjWeUr8hTr2DLt62onq8CR
nek+7E+JIRDE7UNOd2LM9NaTYP0W1jE/xqiUBipH1qEE9GVN4uOAD48awgUDz6y0l6jde5laTJI2
npI6ai33bA/kjwP72jsbz5T4KUJ2vjAuE84c5UAyU0FI4SutUJ0ebqjIfnmug1MokboDInoHCKhs
Su3sXNUyJtgdvU4abju1I/FZ+toLPbTOB/vxtKWo1RKKAVWYjLxi4oVWQOEmDPPZz+M2PPN8vW7d
TMGRVf4EkRYKDAivEkkhJe+7tZn2sSIa93usopoLSWLAj84/0fPyW/NIa4OB+QWF2YZ9TVwbxCRt
JvzuDVLaoBBMVbk8JOcpGuVQNj4vB7HxpW8aJ0bRuUu4d+TqiYWmATazZv1nHGMe/7nL/eMrW2EK
YtvUa4Ctu60xqHSBuTPHymWKPWAi+46aUlUQTAxF1aHmE2BNnpy2ao1qFUX6W7ESqJ/qye9Npsxc
Zt1uedOyaOkEALp6RJD9LGozQtY9KLRMOQy01vdxmZ0O6G6GBo56Y26NdGCrZ5PU4tLzkwb99ozJ
YEnyPMtoGYLqtuJS3VnEWc7BH8j1Tmqk7sJFUb/pub898ErhTUTyJ/S6pONad8A4XrFyZTNKbrOl
Vx1YM5QvVBnOYGkwGqIdQkbr0cv/7DgNI8abTzuAVJPRZcwwigKKIOA579N8JrxLwvpOttsy3VqI
LDr/wpU4jOKfBGP74ubYywn3R6BC3dc4XoqEIMTa34CVXi1/xG0PcQGq7QoBBhHe6t1vI63SpBts
BqKx5XKKVQL6J3Zhb0TRpzhLbpcnWRipbpJnNsqLhzMwECLRVsJ4Q/FAvoYgQzF8KSqzAOZy7rcE
BRDB+SzCZ4TCtfDuKbdEeJso5Q/mSMXNL7cXxsma6ntIFXAxcJ/Jk6Vvib295mXLAIp9p7bpHUPN
ejzfjYHRBQNtevntGbTq9TBNBLQ04qPfFikuROYJec11ZDugGu3TvnXQaUJrREVKXBwt8CXyIHvQ
2iu3sNqGSwzeIEB0uumzmsG+Yk1H0cWT5aTGiTC8VQsWkjLbQs1y5iQRXWLQ/HySGgBodb7HmrjU
TNiPS4WIXIzlj36CMamF9QrHd1TmPWdPgKq5PyN1St3puJJ95voCDcj4l2T2CyFRqDmsp3M3/JPx
B4Cb4oanYt/FrLaQhIB0aAHu7be+cec2lJR0bkKDT1U40lm7S6TAVJ058Ouh5AKHEQlBE77mLKCM
1wX1xHjfdQxAwofCOyQDEQRxhKPviqQ30ViFPECdgCknvljvZ4WQa/EYBDj9C5IiUJgKg053Dho5
DCtvq/1IQpB4GUmvLyiGkk7MhIokL8dOXGKNXILoBPZ18gPwYLzrDWp68s0pu6yjFniRYxIpedYe
NpgzAMCK9lIGiiGT/jt14O6NtlxGEWQ1SpS57rNbqmwV9f0oYmnSyV9Pb/LwDSpiB5Ve5V/xLA0B
R1gaBx5aXMiW7SAcsU5sCpqmUmwyYbqIknt0PMQQ1560bfMvhGz0m/zMkkP5UIxZQZicqfHLKEX7
PL25+uaznjY924JSn1pw9ZS7vdaGXi9CPVLVIWztyd+qxE89MhEx4oEaJsWRB0hOdBTlRJj8ySTE
jCWIwgriysdzgyx0gwetIMLL+y0dIR4fIE3LACdHBOg/2dVi6x39MlJozar9NCCswb+xI6MJviPd
8sCDDau06tndqrvHJ01SE37/jkkP5zNfK6iV7a5ZAhBbp23UrKjgTnTOCtjep4rJ5VhCKaULmv+h
R6DHTYb3slivPzU6jFOsaX567EDT6JtfXVeS7weT7SfFLm00ZCxRKsKRf22BMMD7gCNzhjRqEXH0
O1WrChYWhHUnP7abY0o2KpNIaphWlU0JCEtBDwsx4ifMvgqWQovwu554tjuMdopeUb3+Sn9NIato
aZDnPKB3y4JLtpfaSYZZa0F2Fs/6lMeZ5S0qnsC250EfPPESzOVhrb0cuMW7CwHe0+4F0Yz5mmg3
paquxjA6XH+JgCorEcJNB3E/xFTYTB9tb6EYfIWmYmpxMNWmYvNxakwN/cfQIn/XfKtSouSFxObO
OLR5VTd9+TVm7mCRUoB7e9o6iSqcy1M+rBj/9RUgggMS+UQHeUjSqC8ktWsWr/iEESgkRBe8wOzJ
CqZ/Bk1Mv8gnh/AAEFWG6OGxMH+fXNpNBuNEZQLpm1FP1WX3uWwlTUPmYSHBUhQf60qbCSxNWJco
uoFWQnOkLlYW10iELg10a7nXi6EoQnMdX6Z4VjYiI4eknV1lUG903ASY28e185uMEJ9eEPV/3tGA
Owtbl9sy0+Zij4y0imGuRWHnjfwdti4GEQ5d+3wblQ5vqisjL7EzPr9xCpNGrmFMcHW30AabOFUA
H/V4CB7Ef/VxuOURMtYXEskpZR3tYtUiFBEFPsmYDMZEFwfqV91wfkIHDKE1BGNWEgzZtQojPMDR
P4ldvxBQ3piUiK++BKQVD3dkgGTh/AkTMsJ0B/LbvOk49r771SLMdlohFUcox2VAAgSf4p3RnZcX
6qZz6CrYdOX0Tw+/NcbKXCPPkHPj+J9SCTAYDzpGInPXh0xkj1ADVdIsP2l4wY+7VK6WGbaAiikZ
/LrsZoSn4Iclggatr+/XBS2u+cQEBOxFR/30WrCMHob9krc516i/kNURPCX9ADc3DaHd8rNaSfPf
bUixVbBvcg7GFiKZGJ15WEqI2IkxZGqximpw988P2+W60t6Mk7dC5BrBRnD4l+k7HXnvBV9Uo9QH
T4jdwA+9X9j0gc35RHPwNUJe3Uet8UgosUdawFmvyXpg1IHvlXUZtv9SBvjp8bEQa08RXKmhPSja
XwSUpBZfL/XgZpczH9OuE+pjCe8oZu9CDsuvBEqg8H19B1XUjIChYH6QZKeLRH3CUEH/aPjkhrhP
RyaOJREQMg0RqyRQBu2WcZ48XUVeQaSp0OwY5vaHqPK6RgOzWtJ9PxBl2BI5Tq0ySaordQTQIrZ9
/3UbpPOQZ/u2X2ZIYmdTztYLxr0tytUH8g3oHj4oMQMARGQai+K1AW9XTsBm2WBcq/UfRxEg/koU
xkuyWb8ogWElOudtKln9T+LKytXopKrtrHC9YaxwuelX3DWrsD7l3eMEAipAbKisfOSJ7XUgjpr1
9qXil6GLi4FLDdYC8ExezYNj2DBAmzS7ZLGy1Jqw3xfiSdHHQyzYMbX6nkCufHUE6Ke6jdyVK8eo
5+mOl9GYtU0E7awJd5eVrNz4BeBCmu2gWSxcXWWZBG5jkVjX7NbSMD7VpOW9qkwuZXnRMJvQ+J3H
aRxsl3//zGYGxoiEvS6cIF9wXe3s8LXlIct/3Eq6pGz3MG9ZllNKo8VeDEkiJCFAHtw2UyYMjjps
s/dIVoqqWJlKUAWJtcKil6/JnR4OtVFZoRNt43rJ99XGeUtb172NCDidNcORY60OmasYubVGA5uR
AqfqVA2H0aYOZeeKxzTb0vdTGwRMhmyBO8Bo4wRk/ZraLZncu51FNYytRjWV1LX4hm0DPPpxOyLy
89CisT3+Xagn3sh1JQP3ahX8dcXntszYDcVdk2vvNIij9BjoyJabPTYRkl7oTpQfinSGciMih1u4
NISwYECnx2Z6I205A05Kglys6A8ODwzeldPNe9rJNTnTCnBX/B/ZVY1lLOrO16y1dwOrrHAAOSf4
nruhBR/fDGGFj0jRE3JeWjpTvxP6sXnZXCxb84GLwzFiQsZWDhaKklDmBr++h6oJLxya9+6bk8qk
KIyoFfqAi6Osd9yxdw16AcEe8dzyjENy16lqB6tSkKJ+Bp74YXELGMjm1Acwbcf0dndS4onXM5gb
kU6pJtRF9z++wo/TZalo64i9/nLOZtPWkMDlBbc6BYVABvO+XT4b8E3Lpoks1yMt2G2k1ie9J89W
Mch8yWABNMZStm2dLvpmGzISiVf9GQaIa+KPojQ3XphAjST7x+X4Renz5trmyXApj+SBYA8CK4Vs
ZK8C/N4h5GK37RYkm3zzgpD+lzSanTRQfJ2zmSDsj51dteZQzLYjNBKlrakIJfRYCwBCGAbBYIP7
T9tHLs9z+rUEfnX5+mykBZtyfaK+PNjn6w4wnURvl1HrikD0Wmehv3FRBwzTEiUHOxLjN+bcpvYN
7/XIDBuPrqx4CmDXcUlGX24S50gelLC7gp4UOklLWbUoSJTprrLIR1hl2VMI6+Teui7Kr8RCXlME
u7nH/tNpht4G8UaJp6ZsFnPL/dVqrEcRXi0trD1JQ6BYY8atzqOIgtA/hYSvxft9tPUASMSNrVFy
yMIMHD0uwQ8xKNyjeO4IZh1wWDh/RxyyOaCs12S1YD+1jyDo2WyvYljDPmRJ9Mz45hZOrWBbmSFN
dJ1+84rtUaiPh3CxyQ+NLxTxiFEo9bKHY2nCFFLAkdD26L65umpfmCnsI2PRd6z2ecJzs5U3K9ui
yGXrAzQDb94EmPtYpsN3f/8Z7KXz3dWHYh2HEpukcjYBCFi03PxxEWZn0f04Ok2nBD9rYfG6YXId
hKZORZE8cFBoaosi1o1ZFE8kP6Wlz2tIMjgbGJReGeJ+vOpG0fd8fJDf1auIof+0bbWK8qPTSBOM
5uJouh7MekUkiQK4TSg4nSNY5CHpoibAJo3O60+f0yWsL5ic+2DJDFp8E9/tF0/fJxX5wO8QsjWk
DXJF1aSor98VkjwheV38QYWaxoiTXVvzOcyYWPLwllv2gVC2+L72AJI5bVsiacGh7r5EI7m6sIXS
x9b8SVIANVoIB8Trrj/oPajjm+bbrsGKPbvxBLhRCnh7LAbczVEV9DAHrdnVB6JwnBw+V1bp3O/f
u2RWLfS0Wum3TWOCW+Z5yiPOPu1EY2fOsokZdC8VeVEU8qBE6kUqezaDvVcQlM231no96uaupg3P
JDM484B61Ad3hgHnvUUW9Z2jQI1Jq4ySjRVHTVAvTiPx1PEgvncwTbbV3eM6cvcL3Fxf9nunn0rL
crHGzUv3zLOvAqqgXKO6MlXFiqKOO35nDye8hmFc4TX3e3UfU7Nh5tBum1f1yStFoCP0keP2kIQk
MJzdBHxOb9M/9Ul27a+Fzwhm8ymoXtC6760eHFrQRGer/Bx4uIcMFcUR7NGgQUGrnErupoXdJpOl
nNQUsaCtIQDS4sAf9CtUOscRXrQQPZc7cE9nGOuGzMGgbbQ9X97ikZ5+i3QbF3ZuyimkF0sbPI30
SIgGfMI584e1Aq/IVbPiUhzSQJ3nlQYBAeYkKR+HI5elCl1qUA20x+YgZIRQDpEmAm5gxsoc8gin
YGM5g6LvgYTLwor+Yw8orX8/rJGWjUqAy6epqdcmq7rLovykskDbcPdb30hgZDLqNt8kAj9ndQoG
BB3vpcDNmuoTnouR8EFAWmzDEzHGxvJZ47UBD6FwIcz5S/Ey79FL8ixBH+PzLeKErp+Mabo/EaLg
k6bEe41vvkzjB8vvozHUZnu6jWBBEsRfpvMWOt/dJS7h2aC6bKlztYuUxn25kzbS31jquz6g8PpE
/XgJenGajBDma+oLh6QVJyudjaam6FIOO2h8HM24T/+ehT/rQr3Zlu5oHgRFl5gbFflX2OjSEO7s
LxHfWECKvmQdUsBKsyYtkdHmV7CDHcVDBVUrVdzOaZufeMBG8jdM1wPM14OYJMaXiZ5OINnL576H
nuZsviVPWNEOF9Wd9PWOFCM6d5Erq1K4bNbptgeCt6RkMPRzNd1i1zFGFYqi5S8UnNF/955/LsAE
7PrZXcfGaTbTF8Q4zmR4sELzQMUNZ9HX3ImOwIHjzrrXFwkZnX7PtsvGTh5SqMq6VA5Geeyq/Aof
upqUhwIS8sGHjW3tym0cJKvqjPKeIwk/STsWsh+igww+xI5H2RE15PdMXc1e9ebDzK7Pdy0whPwz
tRk5V/iyRQLpbSgRsCfbbI9AOfb7Mheguqkj6o6dRfYFRewjYW+fYq5UCNS+jHGb/HB9VAuB0k5k
zXhWaHEhy6pGNyzk6k27aqVpJqyUwDT5FeaWpDWIiPaDapy7W3hSSYAkoB0mE1EK3+dEgttKtN1S
neVPjikelGDey8hMFRom1jnOcCnf1nW7tK48ZHXn7SHn+uOGfho8JW5IG8Ll4Q0+W6bgfTfOjgPS
hpsMpYchae0XITReZxzKF1PCsV9Kr+gCnEzRWCUOFpGcqiT+tZV3nBl414Q9BI2oAkkIrJIEar62
tPKshj9Dh7tgIvg4rTsVSOksXl6UOWj05H7BHLqGMokbso3+wLnEX5xdg52L7KFcYqxXzeWmEjDC
HCAkBxcYF+h44DVSzxKGCXguzxTuZTIHCxcTkFx6gPGM8XdDvs9SXcJPoeavURLNcBKSd/7yGAP/
EdezUr5i+4EqEwGOdC0I9uEkYl0dgH3sjJ/m3WmPfKwM/plmeSK0DE+jp8ZyQHn36fJKrAGBINrs
eAv+EBgQzjwwhBHRpTQXdEKW6dKdP/FgdIjimNk4/WggtwdH03eXc3YshdyIpWY4gPCwET9SiB7S
FnWNzuZTEZXAKnVdUx0pDC5DPDcEmCsICNnKPqN1fInm9F68lMMD/YQishk4dHMhHLWzsJtAe0P4
6DJbo/Ed3XY20Iz6nixZUOk6TU1IHD9rXgHl5/ei47JFYkDQzZE+Xnx7xV+k2cZgfaHWYDd43dQn
mvYrFhdh5Vi7RqhYCTJVgUNbvWMjhGOtHJX/TNSiyxLZ6vWZbOQy1BPAuabMMMwWezNEHtB/P+2H
c3YEmsqFShXsmuh0fPqRpwM4LdTuR9WjCDkN/h2bgznJHJ6vO2Dt8DKML1qdck5VX1C3LxBkXnRU
HXQv0h7YnWcAJVHrBUP6STa5R/QZHaAgbPOe05Zp8CrN1sDY9Jsve09deBrtN6mMqCRl8NG153xe
cjkcSjiC88YubWqe0WDi+M5TMix/H/OTCKruMqRhOTcFQS0UyikiRccbySPXHKfa0Loqk4Wa0HgO
jcp3xwv0fPvGVPjTXPjwCGSfosPLXhjgj21SbLix6sdMMWW5BU9K504hnVB310DpUiLm9vsKwqmO
as4oBKgsYasD//kcVuv4Dpv6QRF49ETD5J7gVWCQ/cjerjh5tnyERnhXXAOb1icIbYlxx479QaQp
tU773NqLHLHULbyBd4g6iIOT6JAPo20eAVO8aeh4scqp2/RGojwKhowmYM+nen/8S3mPEt9W6Qer
RYlyoRzWvN0F45i6aaIaw+8MS8lwPSvJgQBuDDEjOKeaHx4qFBxnLf0h4jYN9NFTEb4HWpm/pK2P
KHgcQwJIX6FpcrdVQgcbUNlXlB3asnin5S7TvZpKmdtjFDlc4YEppnAzlwphC0mRco8uSw27KNfc
UHc9TqSQStrRQgiaZNYCNdj9kwrHK/YC2Ck6fvOQp1aVm54ib0EzE32Bn+Y3dClj4S9zuwQxOEHg
YUfepeTZDxu5PRupmZcGH10jGy3R2qjMPiDBuFXQHPbiYSRxGAI3F7A/Rv1Cv7lgkL4T36vbqHNl
OzEurFIvjOztq6y9vzH5s9VEArH1NnVlIhFm5KsuMaL+7HSt759bzfEAdhH3Gh3Ki2cYy51kCTQJ
y78HZynBKdiD0PRQt6UnxmvwI3sfBQkeTpdGFpPDZssDUHB1ByZD1BcsyML4AXfGqxsvBQ10Q29a
3xWw8oYG5njzQmewD5+yWjypbewstDclIdbRw59AGhjVOMHpr00T7CAZGklvQdfu9/lSjnzwvTUN
8AUOGntlpROhVVRE6GWvKxAuW0l4YSOLMf2lCZJMTGGl0Pn3Pmm1UMUI8Tx8bMYtsOy+MuF9wko/
QLxnPJQEBJ4tmf3ZSQbl+Nc+hqozOYLPSu98tgIlxGMOeo7JpnEVE5u7XqU+vTt7jfnmOJ+49HOa
UqqV8Ru6k8cnaIJIGooU99694jgSlbkHmr20Cx9e6acfQqglEaNo4SKpi9zyzw4QNNcC/OoZxIuR
KzXU0zhA+V5mjE/Ure+YmqnP4m+mAAQlzXI0FYTjkBxDux5Ndz9whdsjgc+wlarRzx/sG8RihIyJ
9SnLS6rYyIWIp61DeynlLShh0i0U3+BXieYdje/WAMfVK51P8pRgGwshmGgrI+4CKEKIhBn38Dpp
JM7iZc9Qban12EuRsiWLTmRQar+oRUgiw54Ojo5o+V1bvzE1zRuiCOXVa7OsNVmvMcdWSxMdGtM4
dx4Cb/U71Y+8UvNJvouRxZAKPmTgZlDEPOwkidwx3TcwDGa14bDx/bAT2TDz1DOPSGhVUeI7vL+o
X+nyz5XgkJIzbc1sQ7uK6DK+yrFzYlJlG/NPe7tHq77aBWrNvZwA4MvJE0LDyvrzPtqgBOJU0+lA
/nvjA66qqixUM4XiEKHFzMN9FN5TrEhPfYQ98ASk2CcXHWqlUoWzf2mNAXBzF9/B9Ldswdnokp+b
W0P4Gcshc9H5Yln2ylM2u2dEaLjaIPoeUitHljO1EcJQ0WqwASuS7Diny4k+/jiZeh9NLOcyjNLo
43JUZ63IzMhICyGeM8xP6FjfdmIxIWqkSnnA9zY8AIzbfVQmFKADxNYU6mkjhRsYqw9948DjGyk0
CAEdc2CvD7iLhmwWW8xXhZtz1r7Ulk97gAdfO5i0pSyDWbkh4bvpQHYvlLbgwtWEHsV9TgQDlJbG
lkOC7pd/GeY4/LcIo5B/PBMcVf1uTRqfzs9jrwpQOk2hciwjLdExcpCBDCK36cWRzR2b+PwwS4ON
4p+N5+yr5shMLTm7y4J4YlJB6Am9Z2NpT8i2WmjL7uEjUB3o0d0obW5kJywPH0IrSRzn3IS6gxaB
QupE/krXpmBSs1xjN8urOqspZiAuDV3Ml/FoK4zMWbvTS9JoR1GLSr/+36txVjonFS2ezxmHvr45
b4V4apaOFvkdvk+Ng38orRNY6K9a2wo4gT00H2KrB0o3+2RoHE4uGDNAIrE7wTIOTYPp+/zqLDgM
unacrqztz3+aadbalH4x6Hv125hhXw04DkenGW8a2YzQS16O5+sWuic6sxBBaB6MRd8gBUPnVFi6
Nez9zB+rxAEA6q6RRI4lCKVxLjMHxe12TW09Y0tljS0yw3A+xOABKNoj8vix6yUWeAgJcj9MJd6O
MDii8TaajCncH3OEgyPJKkChDAAvHxR02eQ5/QDcFjMzybDuK9fzFoi9Gpnc4YeRoRR6HlJ507Cq
l91CPkW4QUL5gQs8l/lasmO0ibmaLtf/jjinYtdlfx9WM+bEJEKZ9zmw1NE9cbXjfK0T/aIC1bpz
PyXBZ+x7TnQAhdQgkbJeELCVuS6EjDhtgt9BjaG2wqu5SJQS/GR91sSmxAEZ/DrZeYltTMUdbJV3
klsUlmfuE7TIl+DTziFvdQBI4HbZEIPo6oZg1RMuUGDvGAaUID2yh2SmA5MBTOUl2c2FFli+Issu
2/VBnihTo68JO6Jc1wflI+Pny3jDWJC+wzyXzY67N9UrgTybAG7wbOM71DK0Y1qxi/cTzsuKX4Bu
coMbO7bQI1ScLYiN4XzjvQwftgaLS4RipkIpCMRQxaTzQgtrOKOUKBHorOHtNhRKbWCKWBue5IEy
+eWpq6VWUTY2hrV5uOv7RmYjfZ7tLmcOjXo0p9d+wD5fYdN6XedD32QN6vgoE/CRBSNZR+Geh+CP
T2GhV9NHodVvWNzcg24kuVwAR341xXq9DOVIrQTeqZEZdwDK67Znh8F/LsROuobP5ObQW6/hkBZg
8vHnN/mxj20UZxFvV+Lce1l6aHo2HZX4qJ7PFL/fGGQzgZTy6ym1YkfjkOqBVDVihOxBOILB4gkX
EV1F1yVtZOnrv0LKwho1dLdf1SEPYSDLh45YrR9d0qgRD558CA7mZpXo54GhRm+T8x+LpMLQR3wl
y/ndEFi4meMkfXUiup5ipPUSamig3wugjqognFV0MUV23WdPpih0Z759OOseVGD5RkrG+PBill2d
jfofbJZeTmJ6wCf9lP1TY3TLb+Fw96lgN6WuD6vGPyh4Jn5ZzP7/kkbt6+p3oiEVMNcnrukgUnn5
6Tlnat5Vm9Jx3haVzdlrJvZmxR3wOzxl+VHZhXwtncv3xE9S+DZgrcfunadsthOUgGfc8vwBPaIz
klrYiEZYDuH9PnkEAH9aNhpDRpI8SBJqYWeqQgWgHMgUD+5CFszFuzE2KIEMyFbct8Z4ZzPGRk3o
oFK4gRyHCv2kmDkWar6LrQxiP9I29cijtp5CNlrheAUUTxPCs5iU92Hfe9Lu+Q4ZvVsnkWARgpgI
OWrA5vbhtEGJk8jsgHU3oLLH/FOny1upAmg/LRcLHMth5FvaAvEE51GjomAq/EKkYOv6M1bEq4v7
HlfbhgNlndy7C6xVg4e3fQIgDsvyN2CGKCRBUgBb+/L1lQiGq8DcXVphbAJzK0ePJRtNZYyGR3uz
+ZT2nPl9cC3g/lA8C6ZlcO/4yePU9ivhswS6mHHgrH31w38N/7qIlhvF7o8GlTACoRQQ2vCwN570
WVZc4somHhXlVzhGkMAetNRaik/U9i5N4oMXplrNbcROFT4E45fJYEu0bFX6SQpulNmzzNE+W5Zt
qx+F/dmZWWt7KWzjdh5jL/Ccnf+3AlruF2BdFzkGNSKR6TgSIsrXSczsj6e7UWcPGjzPKvyHoQMo
VBaUtaQ3nnKB6adG1Di28t+f8peL7wgL8fr/WDqr4fK8+sea2KGSAc/5Dl2D9B4RAhGyzKn6WEl/
X2+eZYYUPLk5Z1zSDXarM8Co4hqAYIS8Xg2wrm9iuU01KVqRzKL0gjk/wyw7aUJKeOG2kpj5Uas1
/fd5STg4Eq/3AYkHg2/uiVcew/Xb92BY/ilFytwfOmfA2Y1uUqP+DvRGcMwEPZZzYXpylRTDQdU0
Hmck8dVv0YkHeItF/H/q9cAM40QmCXrFCeWvo7gOgBdYEhwrpnCRisubhfDI7pyMJbQZGpS9+QYr
5JEabVky7RNuYNMoY77+YXKP2sCMPyaAqLhD0agIr7w9VS0fxxeWrX3ulxtQ9FP1JS/f07LMpHCD
+Gtn1t7hpX8AUomQ+NoxKlyKfWwyaUbPO42OEydCj5Gc50bvBZEy28b1fFqfbCwV9swuBi2BkR24
xA7rq/oorAR+XpHGbUVKWaV2gRoNEqmPm8QDyrHczbfXmv5fa8qTsPB1aFX4wTtKOkihtD7LYKdW
Tz3PF4mTbM8etycMM6IR0Vpjr0AInvNPXYqtlEYYav2OWWZcsg3jm905lmotptDDh1VwAwfwrMA1
n20Muy8MEXylIboU2mvfrBSO6+ohAPiW7aFpVmj8lWr8inKZwiGqRrDJJjgM/NW71c0TOalOBGQp
tMEeZ2nU8+f9+jDgSU+UwuXjEeVjw3UXMlr4yBGWXYqbagvp64AahkhqZgysxzkse66VhByh6wLV
r63rIjMiZJbvXL6WySB7wYz//rGM7isz59gwlPdQDa9XgrvJMv+ngZTvCLXXeUksvbwNm6nl/Oql
viBsQyGWdHOXxHagyPfBQfEgSIPGraZjU9ofpznxSGiuCbE+NEBrNdClFNuSvR7uaLVDIa2xMJm+
h14ZHrXXxIQQIFQoiJNKTSEKQzZ0F1eq4oV4k6dlC/sQXpvNlKAX0lKTHvXOYxcgD3xmJKl1ZOld
8ws/20fz1bWKebbTr24JF6mf0+TMg74ZObE0bH33rxgIFaxyH5bSuj8ZCDn82qADzLgxzI4bT1NA
LIKFfCVbuymBcjXOodX7xLZ+uI0oQQ2Qlm5oBfOoQ/Re2Hsk19evRBGB0wv4jMoCRxmBPPLq1dZT
yfeaqjap4nibbF59qHydfB3W/akARU5ihBw11e0J1C1dWQBp2U4hr+3W5JyTi5vnMlu1sscVKhuW
kBs2F6O1xGxw+4KPhsEK9vmuQTO+QusLY4Ly3Lh8FjgEYAzAdCUu+Zay5qJHrw2eK+/xan5dFKxD
B3EhLmVZUcI7MGwNohgJxwYnj3MsTbowXkIc1M+a0j0CsPYZj4y4BxEZ5K9qackLfQRTJB7Ggg6P
JdaAXgoB7MGXIMf/9ngAgIHG0SI39PxigIN0ubCJGIeVfa1cNpJgF1t8caNk3Y45xIF52Ca7pmCz
qGPDf1y497tX2NQ4UYEHiqA8/kbLf2asAnZiDitHLRnl4xqiUg/t6jsxV0aNqmvbJ9Qmd9wmGu5P
7CUqTr7j1Hbnu0x9f3Z6ot53JQfjjVRg+Z0CB27Ymj7sLmoSSjQieD7gWUXeQqvFl+FZl7cx1tKq
xHfy3Cf/UKj0CSGdenBrRldbdeQMdTpFGRPMIuR9TWLpoHSo21apNekKSdYDHdKbM2ntiC9Bd/Mo
CRg77x9JkRQife0vH3wBEkkDcK0Q3gWcguCvh6s8vaa7gysMRelWWUzwMONHSJ5zy1qwH0lF9opN
YJzufPPTCq7VZGaTlI5Fo6GCJ2EWQn9L2JITJ3j2FJAkVqerLBLV1H7fW458I8hpwSgjWfqls9Mm
RjE9biGAeZ12kcUjUX/VUajbQCRE6KfwRlvHZrgRJQs7pTS5WcRPAe30TNQwCmtQH/NbriQFK5hB
ZUI+186+tJbD1qSWyjKhGhmvy0LUXHSuVuT5TccrTjhcijRpj5AOELDEfdnFYsDk0ufUwFnk6Wj5
oGfWGmanCKCl5+mdvotYn5nI9mokzvbpDzaL9UNEXH6tgqzHEb+JIkaL7RZRYrAkyS9QG45ZDzSQ
eqS2MtzHnPUEk3yhRoglPYZFR2XCBqcTQ/kqVnmEJUTiF5o1EB+5FsHc4C/KOVBqbPZsXaJ1lwmf
F6M/BptfwrqCbKRd1QBFLtppjtdFkDEqOniAZmd8ZzBA5c71eRXiqLKxd44H4M3nI9UbQYABO6nG
36en6u0+MW2pCR6F6T3B1ZQMj78kLAhnhwglKNigy3QRHAO64a9XnT2QmQQtj96BNAFWAzGImx19
2veFAzrG4ikuPTDTI+GjkY/22lBY9AGUYSDtV+ng1LsuXKtmq8fRtbXEJ+X6hGsD7b4Z0Yplam7K
LamsvsEQ876+NHqym1EEwwAEUHL9hNGTp3PFRh0xgJBD66yXbQ1UDZCww3L5NwM/sC6VWz365aoh
XSMGCNhr6imVmgofVfB3fP4Lc3rmkGkQYy1mdTFi1IGlJKlYvSK6aRoZEUsukwemGj9oxpW6sI45
lNu/ooYWhOUBLaWVtgS5VgzhtPRhRSJuvvGma2pAB3bMjfZ+JnhzrMSecfeEytVKknPlX5K4mB3n
iC362z2I1uesa8ixRuUgdhyShmn9c+MMzPOfCUVL0OhrUA7bkTC/mg6UYtIRv8z8c3XLD2SHo5GD
MtVh2YKivYHQ9l3ZRawGCzY1w4x6YZJ2ropT8xkWhup80FE7gVqt9SZiXYMrI92nPo1T67obyFGa
N/p1ePfNf2AZBpqOeNpQDObvHNf5fPSJw9ZNBfgTCo3l3fOMtflXzbZ0CG/0S/+BuraJfn0drw17
K+otIrhiS59f0Aiul6pOpKmJXsHxRpJaSbRHRVIU1HdvFIydgC4TpU910SL/5sD4m3nQp/JHz1Wk
HDaMJUZqNOsoLkctI25u2fM1F4QCuABEyRS8+oKAEnDAHjXoA5JiZyRhXMdtFPjhaex6kVIGYqop
zDoQsxnaTKUDLG3q4hyn7eHx2jq4p7njuZqTaSXCW3+QP8IXoO8+uTwjJCP/hete0FJ1RYHnP2Fw
UwK6eoBzFVyVbNoW6/Vy4O6cWbg2XGMDpMgUjbDrrk5+4l+EZKIQc1J2ii00ISm4VjPKfIfrNYbR
mM/24Cw8YZrC7WVhNEmsnuam2Go4gq+ryHeyZK5v+mcrk2KPQlSSlm8fnUqcyB4GEQmYFRHR8uRT
r1jXaQGgh0shgSHDx9pIFYpI1CV+KhPKXGSsZLnzz2coGehf2wkiK0TGDW36OtaEsOLVGYgr2KPC
bTNuZ2YojRjemkw5ciobNII7wQpGmxsUsxT/bctPfHi28haBLTKzNi9EAKJiyRIzoKxDQaFki8tU
nI45y2bezk7Q9yacubcBh8bRdYgCncwvOj2vr6tWfNrQMb1TDHFbKjX11h4jQI6S/1TZHYYS67u9
R1ZSCsVjr3kVCREmtH1okmK1M+S8IOC2KVLoMBZCd47u2PpvKdED2TrzdTZlLQztrxl3xb3XEBw8
vo2zOBmgKpxXLQXadz59nN3XLoe3DYprVR44bZGgFUZi/oAAYmFdmIoj4fpKYxY2n65z4Rsk6UAq
OZltwTI5nNug2SU9RMechI2Scx9fNh7Y7dXQviDLWQIS6EyCC9apzA7UCc3Ee195JuHgN10HFzld
sjEUVU5qyTsE9KlNvICBC1aBdghY4Zx8If76JQfwkAvvcI0+SBnVkvRayNw76yH/cFzWJ6/ncEbk
YQRTegvSZN2UZhW+CmdlCL3n4DjcwyGdVU4Oocv42NuS/3gEkrhcW8MDmBcJOkLSwqKnPuL0wlKa
eQViD4g/UUWRRlHwagjdRPImKm4reTx7Qf/aC6aTm9GBs8gi2VGHyaZBQB9de3RRzxWI3ZWwlnNX
242I+RJGXnTgmdaDwsbp1EZ2oqrainF3UKnC9d+88cXrgI7gon3QKLGudp3i1mcDqkqTB6aFd0ak
F0tO1Osdz1OY81z4hs/Gf2wljVlDkgXRUfqCHDFdiFKKO+Gd09P+o5C7qHhNdYBYeQOK1Oxtu/aZ
hC79tInaahEkO5OE0BlnO07wWaBfo1M0BNvG7Oyq/BHUbTKOdK+h2qzr8Aq29J451zDAHtac9vyC
ICpTdJmAfUJyZ1d+cAjtEtkEPGvOQc7XUNrKv5l1CVkhgFvLYQZNjv7gsd0L0vERFgzcas8TDTHX
2kDuv95XY/Uact47UM1Sojs6jGaVst8YAxx8ENYlHUwGjMMCLjN5qvG4B80jqwrkdzHXS8RZIHUr
goEWBg6YnX1ukqa8M58Xxee9MZx3rgn4PRmyOFrlPRkZA+uCPbnPe/vPzw6TGBvJxvEKEWVKe+I+
3BLxRWJZ2XPQm/k9uPA76C7rWHMD3QuYSSi7L8sNWsDBhP16RGw32+NZDjmM+ff7xO4vZdzCXeQG
58l2PdaaiYrEQvNEc45KvqM/K7R3TVus95NSue7IRMu0zfJNs3LmP+NRjUJy+Z7RoOmwiqh7X8F2
eJnNI+r2fCgW6IqtxtNmuCabV6aBSbd4fLqWV3vp+IizgDi4U0o3xjpfDdHeyobNq0lorwlSYqXE
RZe/82Hew9LuNQZHuKqlQrAUY37Rw6ft9VKGY/3gVI2cQtD5K07e0L5BHRQknmm2uhYRz6BLpaZS
CRXdffyuT+euSJHerim/sc7Agb3iu310SmE1bj3GbE8o49Iyl/8u8KUP5aCXmXwNhN+8wYpPjO84
gRSOtqBz93uJ0Lxg7RP0nRKUG57w+Fq4YM+Wm/h5PWRHcoY4uyC2otVADwAn0Mf33W5IxCXTfAvW
HTMbNs6Hj6srSIe3CdnThvnmOC9hWqGcNX4G1gaEs3mBOgg1xl2214sO3CczFx/Wn0hawiHBsXrS
udPPv+NqK/miH0F4VFeAGTC1W9IaRoIKunQ2AgjLTYDa+Sq3T8Ds/pETL4cwIq+AtFJQOK7gSoIX
mShNpS/4lnXfHh9Z64gPZEXrlWTAKaneMlQWPQLXk/5ei4j5YjZ3A2E1vSjoOG0Ew7+9/fVCtkXU
P5TuBSQftsOzz1thLHNgGDR+0ejrlJipgAdv6mgDejhuDQtgjvcr3LfwYhG3LXVgcj3aLFmKZlUu
JsEAcJxmEQT6ODy7mymzjcV0PFlH1VWAGFqOo9+q5Fobvptz564rTyLkS8+0673gnxuYVDDN5MQ/
Dk6zDafBI69I446n3yvsgJTgmH6T5LYEnc8Ezpi7ru1q8qqizK51sNfs5t6eGTIr6ZGFMbZoWsuE
W3oLkSitMMXDif2C5wfkpJjF8ja5FtynzmcpBYdehvlDPYh4y05veYqvB6B/SkqANhE8edsSZiOY
M/SU5QRslfy8k66zFPvilk78NRJAeoXrwWc43pz+NklGXKUnaqs2wV33C428Fxb9Sf4i5hE6j6lQ
qYsTwuqeSMYna45L8w3zWuW9XIT4rFVMCKzqZvC7lDLTd62zifG/5GeMZnwL9srf54PhTc8wvyQv
BYdZZJRv2J6BMZQWG3qT41NxwbeM3ErWDTbe9YNfh6y/xNRPMboyH4EYfkHedrgka75GqIlOs3/w
7TuIIKKPCz7+KcMOxR5EzyRrMZz8DyoPsupUtCVxRr4gGUAV9c2WViKU7AZ4reQdJBk49VNPdVnv
LbyfkdElCJFUn9D0GPkZ/tiZ6evSQraNnFtID4ifSDQf9cLMFfBenXv9iHROKSZHF95XW5eSuQ/6
7H2Q3TuxgCpTzN0ybksiHsHlSyOh0iDOmQ7ZGQb32tQkrV4RIqt403xg2WAEQu4nuT6mBVZNY6dk
z/ridLGyLXf6r4rFOjUXk5coh6/BOxrM1xS6ijKXr5WX9A+YtbWD+uxlrVAv72SzFvdSog9JX/ln
ORVOgBfz1E6yuC8pt+GHsr1NoQo1ysPphc/TR0udSwvMtdvC2IiU2For82CFPC905KhSC8ruh7Bu
WpzRaamGr3LPkGK9WRzTtFOuTqKLBqOw5nGH2I1x1cRGifhBnFt1pBx1jtk1x7ie/CYIklj2YApb
i3mQVi4u6slKu4ztOPh+gO0CO4wLWS0qmYrCG9Wa1yRaLX4DvpGzRAjE8kQRNJlrMGDIwoLvl9uP
9LlIxlNSAaITXQkFNkCa7wquHNhSQFTVpyVg6ZCTGYwgTMZ3FriegS8qloSRnPaXv1YGWxzp37f1
Te2/q0iBUAtWWX1zRyHBpdJbKg0dWmdpDgLJ2TxOXPjdL+XXv4S7A+g1njuNFj4nDn99K6EsC10m
21ncF/v481NEl2/ijPqbRoOAoknuuXZHiZxL6ydz5kzTipqFSAP4WJVauHpCMNPMnEBqtBcT2mcC
b3bGLeKWRPcoAioFEdnCfzKAYtUXMavmQmQg9IyACJK28Xy5JH4DrR6q2PlWob1nFrU/rc0f2brc
eWLCYLAmYEhqK5WelsuKZN8kYMHqaY9swXaH41QdW6B+JDIpT8Sj//cQZVnx0Lt0hclQGEV6pcWy
A+UjADBFU+CbK5dHhecwQN8SUCL+dnfIz7lvpeNMEL/2ebqcck+xno8JLDR1CoSEVKWfJfx5lis/
P94Zg9QdqfVTp9GRfKZMJhQ1pXuGhRryxozjulj1TCz2976vLOc+3qUnffmsMtk2SEeUnV9Jw3Ww
M36EaSCgM/wuZuUeixxnYDawyH93K33R+JnYa2kxhqckwskoTZNA1DgNsw3nSTHRkx/W7u0qb6mv
izEjKi2yVy2MessaONTqVa0A38e8DMaNRMKGlUX1+L1HYks6rB4QIuHc5bUCZl5Gu+CfyxPAboGF
PGUIubdhk+Vii2Iy/AEcXnF/jJW8/56g+YCFdElDEXQrhTRfky4vxKr09YlTgZe/Fg40/v7yNOnc
oY3RtOiMxONAsTOVIql2o/duy5MbgQ1wMvUGlklLR3FfKODUMU6pudP/kn6w5e7jQlkDAgowSUGx
ZrhaNcpdD8IuWWstE/BEXp7Jc/izo7gagkMaJssJXx1puryKVUS6B8o4Z3wKgarw6ICnHpbGpz2d
wwGwwnqU4JXDZMcElbMaJZlYhxAxc3e3pJrdOHO8xm2Rvy3cZrsljykINTPukfpdXK8d7w6bnM3G
1pULmS2TW6esCp9g4iqLlhYBqIGZ4wq7oML5Kc6rh3wYedvPGGjcIQdkJjsmwWoKPAGAEYigxzwn
FZRN9j9a/ijdskvI0I1tXq8AuglFb6RT7yFV8yt8rYAkX6hGBUB97ZWTNUdcH0a/Pq2+zhRqW2o3
z9v/gIy6mRDAdT4JEFTjsvRzq+cVc/fKFafsO/DIE+jGkNwz6hBK/q7fg1cKv8nIZLdokJkHYtCw
+vLxsXfdVsedoWmZhokL6DUiLz1WNIPtKQ6bNbzYxoslJh+65PaX8tvHQG4JbggtxRyvXw+vJgOA
2Hd7k1v3dN5ugpHz59dh2qtkT3C+pVTcK9m+PQ+EO2YgsPnwRaj/o7lizTmQsN8Hsc5qHv3qqmtS
yJOWqg5K8/uE/xsFQAgT1b63LQ81znoCVMevpzQjOqqO/Ctfd3hJBC2u6eq9rEevt/C1giXZLimD
aDYBPIidKDsupoWSbiCyMo41j6i8rZBFbua0dwH31/DzeirsQGZIYWj2K3jKdJUdhGEw0GZqfisZ
yGYP5gnLuYWcCFUvtQA1yUytpEAA7h1q9o3yCa48s/d8+50WNZLf5UMWtSnigpMungqq4rDVHyw2
7v6kD9mHCfDhtaOg1iBsWgeZJ7B+RzX4Y77VpmJ0V8ugLblS+mn+VP7LTpN30034pSsXcOR+1lhe
FvLF3qwCNnJkX2ayxuNnpikDqvGg+cX+RzmBbzqgR10+TQ79ZQDFSOyHXI6mA0EK9LaCbcFZu9+t
MgGtV4G6yIwd4mIgUyhnauVT+jzGilfxnJCq64v+3hMbn1RXR2bUBRTmBAVcMJdjT0+9oW1Lkq0n
nHuhJUEE0f3euO2rAOq1FhvrrY2xwJkkCudzTepcY8kEqNzwy9jQ1QbRNfa2FXwTR/ldA6rI0BJg
f2FJd7ZnccI7vyu+bkOb4aLu5vt9rVty52F5eRi+mPOQ1sNH3EDmh5zJSpGQ3ppOvXF0NulW/6lq
xWnLz5FRv84l0lf+xVPBgLoUNBVwgnPQd7OrOBT6v/LyMltM+9qjygZBOGUq/Ez3khGwUO2OUaIP
2kQF0SVGAOMXGyDtV0DAi59JQ+TDxcEplQc9olyl1Vn/Alo/wsOUqgQYCor4AyHGwgllzuNJDTHb
z36aL4LaSfISzohpng6pBnecY8UjtHDpmuvJBZL3wJPr/XkYMT4PFdWdUFlHDoyHRn6vOSGM5oe7
QzHyPLo7IxGK19RYRf3DsWXeYoC0sctvaKWMHf8PN3mPyNnMaatmGdPAWsaxmGTals144ywxKD0r
mhvE8ptvdMTPpPhCb/MyOup1d8G96vgG+RjeyyEM+XqYO9cbJat3oGtQmeNW0Ytw8/08B6+ir0an
Yy8unQ7Oh7aUJpmue9X0a5Zq/30/JZJGSkF/WOmuQD9+tbZAtLoFZSNRAGaAVFB3oYQw3YQwP71y
7o0jAaETjE3odZKntvIX0aSUsBW8D8QikYHcLpyb5aAy7G48DUheFG90BtGANsp5N5QoEjtaC042
EZvTcH/WgSQ+4mHPBtqQFxjqq6tEp7asUsC/Ey6glsyoACdbOmJbgswUO4nxjOYy4JeYKPHwgHLr
bnalK6dMWSJsXLKPJ5l/PESlNVBn2jMU3zAWFQ45sD+5F5UWgEIxxayjgUXZKBC+XMOkZNw0OItA
+Yi9a2r4nG730BCuK5L2pJ1CuTm72LBjHnrwMLI14YTAQuzOtVkardhzuLF8UIKtLmQqi3dG24Qt
oQjS0XSaDn18bYM6AJ+FLgv3w4XnMn9oBafzlzYKKj4hMUws6xlGXD+OEke7pIMjsm60ZJpKO9wE
/0wKQnUQ/VtkFalS0S09FX5IOiv5q70ZKChMkcjHcljFM4BtUiw6JFZEyo1/N68/9E2iHnTMkcuB
C08+K7cFuer06d4wJND7XuofZEyM2DBI0plg+yTLOzTk66gdt+U18JP3rrkJBNbjj8oeKQfCt8Xe
DGQufGbqqxtMB4zEPJpRSMuMKBOEOYnrbjPI6n94/lkJ6kBqOlRtGz+qsq+p1snsrfTj3795QD9O
t+WiZfMIYDK9eYOzb35LXVJN5yfcZ4oF9VnymW8ZcZloCPVhtgW9AxlZsbHVD1U9lkcygpQO35vH
5je1qqalAB7UQ3lZymjUjstb1vCRf1KOTTdjUO6E5Vr4nk5RrLwLAw9GjGnxdRQCwUD8YxOnpao+
X0awDldr6xbX9bcNnVNDt2Ovlh/QsLKrJWXKjfAY8fjEff62uFRuuXWP+E8EjBUYNqStIkE6/Eli
4AP+uZ+wSOMMHrgM4oU4ImnEpK3Rvf0B9ZJFj7Fm1sMtcba5MHxpdNU08xKDqnHOwz5JP4Tfmxqm
rRSdzQitkqPyd7GZ2Qa1cE0G2nDFs/qJ6fHEbqSEkhckVQZweXDbn57N10dxpHzGUCIiJ7+6Nyzr
DiODEKxQxhfl06BI+GTBXWtmTge5/FRy0pKlLFWTMkNI9dxsyC3zWUJjMOrKYJFD3UZp+ekZ1l/K
Q8oh5Ub/r8YIUmWmTm9A5wVOxb730Mg/eqw6QV5lodkCwaWTR1l9d183anZ/p6AwtSo9zCp9MoM6
kmRom0jRaLIdKOfndsSyDeFe/IZf+CGQ5PunDoxYJGsK6NWYZJOZYuVlTAuJyPGXc67IMzt8iwny
Eva+GDj6sRXjEGXbPUhgi8JjWpkWqvMAUNA1mrSUqAoLAXqIfHq/D19GgF0bcafsZlgNbMArhHRM
H8w/dmicSHf1iUodal/Efty/RHd9avkoWoZf2C85MLBoI8VQOWXrVb7X1oi5odKtkV5E1kkd2yPn
FBwdAtWgzjbIBXl4Ghro/N55SBg6p06+u6zk9t13Tar2k4b0Bp5+E0r6tB7sezNmDN5SmYUWXE/5
kzJWvZPtYkZtk9CboyiI445A5B6ZovORUtd9jX5I6VW6GXQBp/fvJifinmEA99gHXiy187KQqICx
C3D9FoYRXWF1PTmBpzNOvf0HQBSK0Ena3UF1RsPX8BTFbB+txfkkhy23jF5QZpg+y8njINYRWLbQ
ADVm1tKRZpcdQuf7HaD2g8Dte/E8cJ/Pk6EmehvA2EQdu6/euFZEqzQhKPc1uyeFGnqrzBj3/2zM
cd6kv6cLGRApUEoEVsqTpcqiHt2ARIXRS+kR1vj7avuQv/pV7ie7JgQ9Xhf36hErpwT4lcym9qZ+
JnFHq9kQaYKpv6rU3FVZgebZ9jFBx7/eQNK/4dHA+IibrkWJjXcBv3n7Gt6Ka9ImYDClaKdAIJT7
3Cdi6Dyh3WK1SbDiU/WYlKmsEOxk40LI5d5NRNfcSJOzfgin64fFlle764Bw2vH8UevVLbEHMUNj
ncCP+2bKbGiLHj8OIaqS2enW4pTphObuTMwLdyZvMDWogbt0aNshhtGDw2rTq4ALF5snuX8xMUuL
gl3vUHiCTxMkYgV/VSyzVckdqewLkHqA9IxwGpzR8m/FE6tG20P5r9f5TQlQvQdxMRk3ihiLvZoB
wnT4/XH4k1i361BanKLha+OtjpOk8WtFUxZYzkwdBSWBrQ6LIt09DzA0TfWsFf7nzi7kO+8mOgDc
zj2dTZtqqOQic/ZOEynbl2t6SJJAVsPqMVLDu/M+2JXQ2XlslLy4DxDNMdNBK2AWftc6ezypMaaf
SYA+P7eqJoBaegwMJ54ufL9YXsBe17lK9VHOXnix2OE2Pr+Op4yFEQuoaxnjppXf5fuHs0w/wDVR
jCltDBAGAiQT9yw1ql0TtA6raZst+x5BYTK0Kg+jxmTV/tw9vG1FSMIIGvdrQ8uxJh2sNtNbdKZ8
CXxeeb+92LxooRKAj6WkIDceoFsPHlqBmavzzdxPsANv6BV/GT+4gHYZe+5ll+DUGzkfpHJk5iJs
zxq000f7+9gbYU7Dtj/h7ytfV+Iw49bcA6RPublCeUNLfNlD1nplqEG3EN+zkQQcbYZl14bEQjYv
QnxKrZuH4u25/ngPE9Lm8wgZjG0zvcJRq8b9cYr0fVMTo6DQkSf3ruM7nqN/NldBgsxT1GAvdCkv
2szbXIty4hjW7nFUnlK/hg3Y7AuUtWRBoZpQ00eecH0bQ/IBCBt/cYWsHc/VPQ44Bk+ZJv0ketgE
OET4BSWAGsiJyOOPJgbFKnbUnSq4r9goV6nE4xiCT17gxok54keB5xv/z7QnVb/xKWakCEuUvdoj
TQ5LDUB8nem7ZUJJmvBvj8xrnvyW/y4ffKCi/Gf2p05mgojghxb8Dd8XGD0d8UA0jGTIM6jiYeai
6RrcZTi4Y2wJmUKmWUOqcOnCcxa+DfeLAJHe3bH7oZE5fKxYcYkzqDvJxK4/gQYlpbo/T45xvwE8
UwU+2KmsteJsGHIr/RbGXBqUcJFCwF6uA3QN65oV3GsKgNs9Wo8tA701iNEXGgt6eOuKCDLCBCv7
kv2lErKyimqCS6IuvYFEtz6FMlgpmUFy8wkS3lTwmR/hnzRo8iSckCUjNh2KYsvHmyh1PgbkdO7e
xXaSRp7bVbuFE4wYgrIpsakje/AHWek7su+XwMAK++WNfClpzgc5Ln1/8kHnWW3XQUqGQrxOhndU
62lfu0bn+QiJzul5vW7wR/ysXATxntECA2+Lxn6uQdoMSdFaqcUZ8M/h3OAtG7FfLNrfh/Wgxle+
VmEkfJK8+9Dte4TmX4zyD8g3ZafptKooMFS7Zow130lvs3seaAICdHqn0LMdOLloJTl/lR2rdz/n
hCntEbmuzYQEGbzANIjM1nID3uDQG3k+TW5RxT/hz1VShWZnavzO5sBJzdy8EKHg7HNIyhh/0LzE
muyer2duvF/RbsaCfst3Iu5eCyqdE7O9K6zHoHNlYKlBUpIaB7Z87NBIUfbCPVktgFefC+yNeIRC
pL564YyY4tmSDAsoMLyiO3LId3nbO5f04I1wAZmKkyBa/NFLQwbDnYcAsfSyXB/Lqr1gVWOl7nIW
Y1BqLDjESi+SeqeK6eD5hQPhvH5MA5Lx1bAiB49AR5KeFZPnWIO1Xv5yO7zOa9Vo6NfpzbIxyFBI
rLtEZ2W8/rQB6crb0EOEYGpBdrq6KGhjrZUHlVQgwEl3YwFauhvuxUJBi7Pysb0IXahhf7gj+5j7
O07RjBZ7IbCqtLJ4dKirzwfmF7KPkct2zOd5ijXdujufn4A00O1kHZihs5d5WhMSb9ILQZWb/saR
yxbg5JsYmBRfCHRoAOWXmHGfv/KlNk+T6nQM9BA8x5A6/sBjjRAyNQ9jisCfUl4HbLiYUTjtIhOz
yutfENSvpOGCPu+iYoDDeVWd0dvY9LSgkCLjjCPIppaXTBGSo5L99CPHgQt2xgQboSQnvMGQj6KD
BoPGsx+mhPd/QAHwHzBKhXfSdObSXLb7PW9pW/vxBL2jve2o3H2oXdyk9LZE5IRrW+kXatcePs2h
XFeBc8JwHI11ffp7F/RsPcHXR5jxVH/IE6+3OEHz0U4p5McHcT3tE2Rr4U7RqlpweI3XDKtyXQPv
xAeko+gyvIFc6gc/2xzRValCD58NRHM8vGC6hF5zkc5bf1Q6+PqFsVw6NnXjdzkIbhfbwMSzwNlf
mpniqrVdZarekZ7JBim+Bwlxp0XcyX2r2+Vnumwa7X9Ggt2KFaXQirGI6sI/b6QmTYzwVFBc1oJl
jwpIYikEtMT0VX2tyUul7Q9F+bvHTAMyRqqPTC6YYxifpCu83vVJI3WrsaNlHIHUvq4XRv125ByN
YfLQAjCblKWcYIEZ/8KIYSNUHwriRcC8M/4uv/rfPNYHtZQC7mIi8jPoPNw+d60EgIQ6BM+f/RZb
dxnkgIk9t9HsEldFJq4wkc0EBMbeqXi1F/qzItj7qrOE5Stn/m3hh1FzOm+xI2pnz+9VV2EzMCL4
6750tbfZDqXhrIGyYMTlmmqPZWCgn/inIPZqCIF/J0MsTAwURSpzBhOz34nb7VfATjiXgd559CnL
DtGSAu5tnCQzVRQdTh3Fy3gudU+G9Zb/XP04AZ6eD5tw/9YTewy0KFZxUD1Yek/JRc0ZrV/C+QMn
XSTRiUPQBdEyLL8Dn76YZbD6SFCtLZblz4/24OTyEBBAdpzpB2TxugG6InF8aL4amMErRfKctZyZ
BOmNMt942T6HlOeJVk0l+nGVCzlYDMwcdHMBYxCiOj7KlVl9Tqk8+ioAYJH6C1cw/tKo1i5fV48v
dwCtPowwAm/KmKwn8CFe+xF2S1nGOqg5om929lZRvbETbTdtEi8FudWkVZ7FuZGJnZklEbwrV3na
ZLph/wdyruOrJgFcHKk0OizAhcF2NIglsO0JevlDZomoT+J2KLIfI4wzxliWVeqFt1UOCugR7cYV
J6T18UroTpnemjJTzoOENfce955o20Rfvli8ypQUODEdxnLUaOCP7h63IaH0otKP7PJo6R57HKZD
kHFYFe7H3MFSAhoGU7gXvIykBcdRSbr7NJxx9m7xCPmlFtIQiPL77fAIckNh5XCjEKsld6v3ZlxF
oAbifAJeeZjyJDOFFgb15Uxh3rQ1EITuk53f7J/NOirsvQ4+RLdHTeMrCafpC24VnHYpm/tPRReI
QKrztHZc3zjk3tJHGCXsrjkxMJNETvkxgcx4nDZfL4OrLpCKDIkE7Ct6vcxW5QaJcm9+wEEdcBb+
IpoUHjNaT/tAE8CUybCZP8Ja4ZjcvCOeBpVSB6z5TY1ySCBkZptMiof6Vt+5sUtzzrqnjG+G0JYT
28ilKGO0ENcCPlwZyNzxqe/hnAP47maWFdkY/Ni8AUmPF+5fF0x1kpenPVpr+sanWPwttAt2rpO2
LOHllEa8P9jtuM+OJdsuwQQQ9C8vA52kWLhqlRlxb8IMe5HLCSNVHjDxgslWn7VoNxBXEyrq4Bqz
r0jz8YmGCCToaCci3gZ5H4VVsXkr9chZkJo64f0BISz7f0KIcH7msiy0FI5sH9DZOOo13nzO21sy
DYmydZ2YAKbG4H225NrtecSIsiFydEQzlmNZAezFFF6mgyAmJAzK1lSsJ0qBbX9IGuGgLUycFYAa
+pkohGHnR+5BfdSjCP9jDGEJ9MjIuoWuWDKr6IQZGAxCdU+AatP9GvADsF0kR/+Fa/1nXTrgqpah
MqOJwA3RAwO++QOueAGeK8OE27TZkDHmX3TDGWm05LfdZM9hlwHIdwRGG71M7gdBgZ7wkp5qIw5o
E2m1OotocbMBMA0cTW6lNTFBKNl5Da32S7/HiLsjtPskhjiotYk+ByyyUcMSkWQAf+K6VfqEOcyr
Go0tkDqe1rOCJOM4Xt2rc3N3W+Yzqoc4Kp/67esSiN9jDWMEh8sqXZ+LRQy5OhWAOyzQ6uxnk9qN
upYGoT0SL16oYC1i9PoLOrSsoDkQLAB61cqYM63M36I2RdUqC0gl0cFzf+Dxe2GKlKNuZY3kxX6g
JrNBTDHNGTpmuO4NKJSFW4oCJC6zzJZ5fCsG1NZksCS4leQe9Tf7ykFNnjkn/GZDttL64YOglGDs
Fg6/UHPD7NcNzGftFcv4NfIsSUqT1rVJU0CaMRZzKPDX9RlYV+AYxq/OODN/XAD6aHRXzyisn5eA
5z7S3+8U++54citJu4f+0W/rWDiPLi+Wa/uSn2v/8lrh6NqqnzxsCZxinv3KQU/YYyOk1kBuS3Wb
/1TygSQbSYzNmoJ7UOJI+aqGDZxKI3anR6QgvtXrTx0dY9SrkptWnXfPi0TY6aXL6ZRfPdxaQyOU
JNYvvV5fqomVSZ4psgyjoxpoV0EoNT/fHKNSPqRGne1k2Lij6DtSOixzSRehPIsatJ/r2DYKW6Ld
ZzkyZmxbbjZtAemm3nFPMgn2xbDvkDIlk5x45b6gi/LmqsUGvTxPZYJ6HkR6KDpMb/5PJvIt7OsU
Fx+HDx71MlWnIG2PUt45rXXZ+eovUFKexpOuKMxH2kVDwGc0DWU/Lp1r4OII+J03GLEjUU68HJrc
SM7ir99bbf2k1k7qqCCDbPDHWcgGKIV8kt6rLDPKMHj9USyS5XbddSMmmpdqabdqMU8aKmDuv8Uq
+1NWC9VCYEmwQ1QdJ2zXH3Lihc2Gz3r25+1Ve7SmtX5ow4R24dePk3EN3wMjaVq/1MSXda9Edpqx
nJmKt6tkV6+GAOs4XvMnFzsZ2K7LfApn4y8AKZYNOQPMrbOnUXgHUoGMTMrnxTQuIqPR/Ml1ES5N
U9OFQclOYjFTkvmGxR6wEKWK0jKwzr3WI0QSRdUL3rD0d0QdPVCDfFZ8Pn1zLnF3SFuXhuBncxq5
KCQdl+z7UJEVJZ7hoFw9yNmvF9SMEbvex3kVM5AzUV+kwcd9yW9dCWTw6Gs4/HfedlNgE6qlcoQa
N4Fl/PtsgP01jUjE2pmCQAC5WzZPvypT1mfje6bNovuYkuHo8kHmdT8SPtokmbOdn6M2hHnvY0Qy
Ce18Hixw4R7EnuILwP2K2Q7PfrClc39cxRScYIb7l1OvXltb/SaKOkANUZnxJMUbpUeivFbenNzj
X2ygoC2lWxx0TjT41srnzYCfLSANVnadTH8EL9aTzxRsJF0Ljdt3oDAqm9WzvB9zsJEMdjhXPXnk
sumviE7uiPOr+zyjFv0cpVohtgWdB3AxV6rCnFSevXqXrihP34nMT5P6ja1TL1IU9WddSMMcQ9ng
oDWQg0P8YjDVnV9KBu5chL07INWzvcLnPpAdErEnGAsDxAZDSIrXo6NDO2hR1WBFGQkSncaI4C2M
5yI6YabHolj9+Acr+B21wFs129WDdtDPOQYSncYbFnuVgvpnlVLF14KOx5z7k5g1j5uB4lmbSjxr
Jyo6lJflqqPuRbgk4kGys6JZ1IAtjfsRO6v/AuiEeu6CXMiX51kJYyg93dni254GDIZM/YsV1I1o
LobpU8gfySDivVVJRh1LE+QTkpxjoQYjWjAkBWpovn6mYFcVaQyxVbdW5eg8yEmDIlZIM8RY14N9
JNMWWOsmE925UNLXUj0CmRP5p/L7tFLUFcGrd9T+mcMjNSBQXEB1r+DOywZ0I12i1RfLe1bZy0wF
DQA9J97sAVm74B+C14Hs01yNhSvr/9i0q1tVBCan8ed03lW5ftMcRzCQg69AbCzqqqUPcV5UJkvJ
SWeo/oTKGw1+CzpTBYxnch+vMXZ5CTItySjJRjHL2EbMcSSXAFEHMJZALjMZ05PTahSMIljb0JiO
NxlvbWQERvwSQZV6hZpuVB0rzuCwYmQNQfxSP+SbXlUvBU2Lo1SmGeAPLb2Iqcvx1WWbypa36rtx
dcM2qcdR3ok4W/PI5A2P8GjPC0WRrZbhzcVeBjJSp2ocWD+MkJWz5myZzVzfZH42sZsf4vECFPlG
ca33SlzVQ7en2Z1ypJzWyGui3CKWvwj2pv6CO8frbals4IKZDacAqv72M2sxLOh+GdufoKKgBuBx
yyLkXsklu/99pt1/8FCLjRKsAQhmp4aGHvlC54gdVX7lA6U+jf29eMvOAwIpZIwYWwXvReZtjBs6
j6guGNhssJ7KE7FT4DnGz8TqWPFBMM/00Tdw/gfa/FpYv2FD8eJZf8VZxMe1DViDq21dDXCjkaMS
wSuQdvuf4QMKA1BgqvLP/+oFyp+46qnrTJoFLwWoct6jztLcHeoso95PCaCHewViKOufLE3Swx+X
M2rqJp8rGdf3c60KU5ZY9UKrSavDb7A643t22jl4bh6xr9VjuR4V/r+GqdBK10rtmxUdordGaj45
kQuNJEGamlF5gwONXZItxaV3tdnT4YKEgWsIaV+/5OG9a0ro9TdApzvBAjDyQHsdyrhA12oagD8W
BZ66RIWjjcRCzR9XKHCEPK5OLOdNzOoj3DuNpAQyPNUzJTiUR/zvDrdy43IKn9Pfk7/VyqahObPG
aR2UzE6s+4hE3as8J047IEPxEvrky5iR9L02AIvxuRJ9CJwXPekXP2Tw5Vt7+9EAKdshfz6ne38n
kjkNee9/YnOXrfuJDAEzo2yCdrXQddmoZjdqZ3h7qM0Mg5dGOcHjhhCTg1ele9iiF2KuB2X3OyzF
v6USpzorz1QdIC0DpFBX5QzvZtnWlSE0xi0RpH3oSA5UYu4G11HkJZ0q9OQ8xXlV4asrpeWPxGlt
FrG2rjDtrdO0asTTMgSjs/uP3dydhY3VK1FwbZ07EVaDs4nTIZajno7/ivetKKn+TXbDNWLJoh0z
DqW6iGexSqxX/QH7aedVhvLNTjsyZReZ0Sw7KiXQpegv0BV7dAZ7hrUQRA+TIc33Ec0JUXiFBX1V
Z3FCHRPhNVWVSEgY/Q9QH1jlxb1XnBwACvT85oV0mc5kadxFFfDHvmgg+bQSccjHWMLW22xVgkJH
0Q9YuV82KwfXVmmrL2SnCgBNWOQARXm6jjurbxDX3Dd8ko/g0mEgsOFOZJWjLQdzTWUkuYFZh2El
g+V0+bR2kgivSp215BMw9EV0gdan5Nn9GgfEwaL1gSTsrJCmUqkNeePbnt0iaqEfgl9gKikn2pJg
uCzgOnMWDnQEMZyhJUi2ELA8cFZBZIuWo4nwnMt2tiaAEk978AW27mlZJ9kFlGROBU4+5lqHdhft
HVERcb5+MCss3ke7m3CmTTGnPUEhX3qjrFwOCpXvqf/JNHB9uuj2rMNyPmRESNXan8Dr26CcukYM
hSRtnc44iIks71D45wxduozsRYWN097MZ+F+PjM1mKVz89T9ZVP7ME1Kjli6nphVnk+aeSnoqzcC
FzHPJcNjI55onSM/moFBJ/BXZBjMkXzZSLdzSKheGk0Jv1zjK5hEK2RLkBVGeVyDJEdhEgilG9Hg
dWc67KhO31/H6pBwpQRrkdFXTcgKh2IaDFkzt7XsXL1Mx8dRcQ2MnlUWyjoQWZCCXInptpDTdOu5
X5anmx6dmOJqg7uuIh4gYya07bx49fdp1wOfmOQXcJ/gYZvN0pYs7iLGeYcJcjuDRGph0aDAFd2l
CN5aB/H/zri6qtzGlRCQpPpwR9Ta0/0OwlT8p3B5aP+VUCH2TqDwUFaWxeiA/j1RvcvEchOV0Cr8
AytkYN4FVpYVfs7N9IRY+EZZZlW+7nGKe5D7oUirSae0muhhQB139Vq1/Bo4RctpZIPDvBBowpEN
XAvv3jv+V1DV2Ks4nM0RGIotHu7BuV4PszwOe46DHMqrqqPQ+ZqYF5/NDKpag4Q399nHjcAybX2a
T2oAe8s9hvUU1P4KI3a0FwUbzptmfInhPI46MHOMZ+rKdB1UtTukqKq9e/q/ByjyM7haIRJPIabS
rY2/wNHi4C0Zv8a6jLT4mkvwtMXOFP14OwFElfAdP6hPQYcmmi/lLclFDE/Bx5Wtkty8P1Ks2hRG
W0g/8vi9b8XUgtiyj/UXIoYV1fj6Aq2IFumzHoq4xvYKgYNX5iDyRj/LoSKP0f6BrsEwQaXusB1g
a5PpEAtN2rQpTG6jeUQoo5qzmnQpuVscj10Boxftnppd1fBplRed7xbF1tRJEOVy/emKPLZO3r8C
0+QbwQSAXfOhKYWfiwo1eOm4ncBFIEx+Y+eUks+8jLj9P9s5Ft0+o0k528ikxBODcAyNUSjJye+j
7ejYqEygnj6aesxFNs+Am0CXJ3aO1TF8RQTubF47GbRImu0eFDK5NedD7PQFDsApmkLVsOMW7h5k
bD7qKYRO9n7ehtHVDR9fxBBOhGIvKqzU2fEhnHy4uS7anrV0kMbvtD25/+EXokQu7Y254Nt2frb1
tpTl+MJx6+1iNNO56LsdgPFwb85eo0OSOwQILfgGV6kM8hMHb6jbX5SLAk8lSWQDbLbc7Ghttjj4
o+kTY8TGmYscql404NJwHyD7BujesZC8T+eYN5rtlZBo/5SWLdpPXT4uuJATPGzU28zOeV7Br9xU
ztDlC4k6xEN9ef+LUs4xKWpWBo3SfJSfTOpv2v2/nCzM4bRLicPujkR3oQ09TNlgt2AuL3TXFTKa
363xoonmuVojEhZDHjBgmvz8weOx7jOsKSZpSDBQJ60wbEth9JTQzaaUuYSqQA2HRaDjMIAcOOdP
H8lcv2Fk8j/Ggvoq2vD39qI81acOyWwcYEz/W26P6tggbiTD3KjQpkDhTdalvg1S89J+VveAPCM/
nI23VCMOE3oQr2osM8/+ftlOt/DshkD0olTLcvzq/U/BCXSwwLj9aSUtfts5PvWAqYbKrW6ZVmb0
6ycd+N8L6EXD28AVMY47sFam+FOoE2Spj5nob4+I9FFlK3RbcDGe849BlVFuiVaCF2aO52nhLVdp
4aqCVtizW4Ynv+manRbnAu6cQL/wr3TERz3qkfB2WxOG6F0P9MBYME7baVdJfyqvHT5q0fHQ4fNT
nLmdeZJgQXvHRH9q/ppThmklnlrbukDeBgQoUgVf8LLK8N7lgcd9RI4xqvmoBsrLwKVnxskX/jFF
ZkV9lPK6gOzmcp2WDT9+YEM2P20XJrs80cSPskRdNqhKLOPrssf7VKWrO/iTCT/KEsk0NNycFHQC
TYsaa/0JdVy+AF4xSWyS3Jqrbtw7a3DJpFzqp5FS3SbMEO2AzE0o9xGblat9CA0jh63mv3E4KN/i
ZoUSZ87ulf6JFs0O7mbnxVJOg6hfDM1J6FgGX4eNvC8Wi/kCRWze3eIofiZ8EyorOcnYYuSWeuYD
H40FNsIHKvueAOlciF6Wwv1TUxNrgHXsGoigKUVXSy6ReYVoqGPz9fylWqDgdYdUwSYZy8ybBPab
4fuF6qICV7M8p1ge2gP/pE3JdJysF3kleRPSHlAOVD/hw68quEZqeCighMQjSa1zu/Po/FVToJZO
e1DudgYHRwFm3qL1f1Rlnb7ttDn2ZW/uggAZqfI18gJVn/EDUP+x78Zqq5blvfaF/GtfEbGlxRac
141P0KDc+DAxcMHy+R5gajDGu5p/kcAtfEQX7ulTRktfK+HtrqZlyGMUxJEal/UNBc2TT7U77V2i
a79sqy0AiBLLKW3B6eOsTREZZsolf7eSvLQR0yhm/ohgOXL4AXz+R8F0g+tifPRDbLFt0mWKWVvF
P4qoQUfqAzHuQdNDcDA5C2cF8koHOmYHHxANpoTuyEIQNLizV/6wC99v0oWgSzp2sLEuOa95/Hh4
v71tc+LdvUmOautDmYlQtq+8ZysunZ+e/BboBO8rKKEHYRGlN2XEuEw6ELPwQpEEzKLIm9eR9MWs
axhi7hPg/od8aDXhwV/3w1Z0D4b1Bupcw+YrGHo+rLv9hHenxNErk6Nls5f9mWSL/Rbj3V+rgBc8
OKdTHSxmfsHn3Iq55mwSNUHlws8dcPRHnANEPBtU27RXU5ZnaDapmJrvhGNWygRBovPZBZGVtvpa
i3Hxp48paeXNGjmH54yRpffH0/qMaPpVtWyP6AyjjqiNIbCoVWb8DhiRmSZ/+IoWcUh7MVWiAUuK
QRCccqh8N5OG6jIXdeeBxI3/3o+0FkJxL60ZxBmJM+8BfCsAAwOOAkAxcM6s3NSz0ScEnmky9Vkn
epyNnJDX4kiR3Nt7n1mh7cZOhUDhjGps6W7NSPcaVChGo7pPO312+jmgEZMxcf2a5ASy+2HMaQvS
2IrJK1elXb3HGqSw4rvL8fzXPMp/6SZfmQLwRIxR9OjTJsnErRdCwh9b3PPiWkFCyuZnGHKGcd6u
T/XdVhs1/zBeVKj/MpRoad9TaEiER9JzLQERxwyL00U8X4gCYIupwzSpvrPcmMrXd8gKmnIyBfN2
tmiRk5H9zDXmwwxGUdI5jbyOHpvflj9o2gQbHhBsf/EFSp0SvQ5fAbe5DWF17/L5WbM+72HH33gM
fprYrVuYYIlmRjPeafWuLe56OVj32D+gyVFApCVlvDhz3ZNar8+N9V6U/y21H4tK3goKc0r3qju6
sEKtnQ+PTLnA/0L4reFMnGeWcUCL45o5jVPGT1s0P4Wjxl8aOn7dtjCZy7zgtRzORH2o9uckHTWN
1Wa9oi5p60As/egxU8+D4okBIDxzAc9evWlqbLSQ7f6kbYlZN2oahaJMV1hz6WNwUv8AYadFaw3j
COvXXLjpaI3otRDWIlmmq/vA+z+Mxi3+ofiZ8cY129jT0pTKvkgtM4fL+t+V2tWwKSSCeOWuVGRr
QzzmIIT84NDHFlbsYvoXQ0jzcxf3C6LhuIaFdPQF+jcnvGZNAtrJvkmBlE4BLVasPsqjSIxCjdFY
SdkMW7A4nj0TcEhJkP4YTx9Q3gz81dVJrrZQPV8t37h/TEqxg9UI7MmaWflmoj5NKFA+K++SJt1p
kJWVQBIJrkC6UHVyF9ubonQmF2TXwo9AItptMfIjHNBVo42zM16nWFsGowPFCC7KhZ/eyk6lGOTw
zM4SPWLyEXdlO66f3hlokC8NyXNJ8Oa4n++abtnhGr2ipVcmeLlmm2bNiuUMIt3IHJJOp2csyfrV
uqtobVKqlPcP2G4jLGG6VV5sOSRIEX6qGZ7wNmxmxviwSfgigs4O8GVbN/jF/4X+xmN6lpvD7yBv
GCHHem8cMactslKh1RjilL+YeQLK3szQTDNrBnUJx/axUHNsSFdahmmWxyvYLcVKoOpabAM0Ip6i
6hLeQRqboHil4RcXiM1fHtjZUUh63+VQprMJCdpPkzOqgg5vzlui1vNvUd2FUyH1NknCQ/AwuH4Q
ZZgjAGOsDHgh8kDSG0eLglHaK3K1cLzSO+x+AlMJu3TL4lWiXJaeWGSKkI/VgtL6ffDpk0ufHP+S
DXKUAILUAtNCqh5p/Ml8euFyEDwXjRsqLMbQnfQjHCKgp7nAfabfvA2ANPXYcWfm4/BuQR47wGI2
bLQnQc47oWgfa1EpXn8NLI1Cu1Q3fkc4ErWyTdulxHnngn1TPIyb0sEMGmiHx2llRpNNFw+I2emn
wtDS8isgp147hIEaKMG9WyENXti3F+ieyg/jH6rUHq5gjebauU6mRBcIbbMq9h8yMLL51PTC2npb
+E5/+5rYf1bItefKnB7eiOVL6EV9ARPvxHz2QsF3j49PX0/D33rs/WfOIrLSxcvtOxM8q/XnCUol
kuW3GAVTpfobuQftyCVaJ6T/GQHaSSXsGWr4SICMZ1ULXfdQcq3AwYwgNeiRu2t3YFN3wYg5CBXB
RyqZhvIGjstGysP8DFPbacq0Qzd9Ce9F/jSP8ffEs304SAcmk2k39+4WCe9eE4SWPdWAaXMiUro4
1SZcnTFdvnyvS83519M7FSJXzmM+NVuRfUEsoQ+r8iaa93CaAF31mvPE4yVL0QXVZaU9ahz9GpN2
lpW6yS75Lv1TQfEfjLm+vbRnGhc2y3laOFEkiNs7VjtUkgRye0D6fYEj8pn+4eSRN0wdElbr8f4o
1ddhVq/oW0ODXThlDGucxB6IiKq/c6svEtHJqeTObh+YqTVGdfdWksMJaayG1HxJ6y4zh3i3qmCB
V26AQS3GcfpO+/TRr9O3qHtIMOTKJuF7ruKG79WCAt0v7XlSWURogJoFTN0DoyPsizhag9BaaXRQ
0nPeHt4CVM8Cm+dB93+fwJ2wfX9P6M0bpWyBmeU8aIxQyPG/gF2Z8mS/DH4KO2pxylVXKDIgo6Gv
qD3VBpAvBuMQOtAVtxqsS0xOgc2wKMkMn0JkKL8ANclqhPO63OA9D4QHOfsdBiZHMrwVJeyADdEC
2YTRoCPnIGZDedCmzJF/CHQepy0PTiuebhshgUrZzXspeG4VI+1fQciJiyPcOkW97D/DfOwjIFf7
ER8BbpaIDPuwuPKt8WZBgM7qoYJqoPHYrmmw43hAsNzNQwqokXJqG628ezxNpMiYKg5kkzMnkwou
+4bYLb0oJE/pwicJP0UdOEs+tw6piuqw6+S1QY4X87Pmx8WWx2/ByTDKojHO3QnISHG7L5bmTvbO
BAOQrN0bnhnY+3HjJcAAqRCMxblctXZww9g1Ys7IofPKxsuycsFioN9h8BH2VeDNv2k1T0oTmljR
L4Mow+Vlu0dKwVnN5K8Qljqy6iybykdSwXh0mSyEQUt+adOHm+0ycZOcYYLMgewCjze6u8eoGJ/j
2MhdTBfIKpPbOjixsWJJKvmxfm0HPKfFsU8dJ1KZwbtIwpVF6VEXUB4HrSMI0U0TY/GMlcdFwcZ7
xAu+M/9OVWziEfeCweP5JC6Dvv66H/6MDMLxem83S+A6caVxs44Q34hDPAFkKPGtO1N6pOb2L6In
uuRWycXKXLKoDf6NfbcqSq/GCw/lsuN/+3xYxxvzeQBOWTDcQ2dXzopYPr+AWw3IbfTiiQMeqXHB
q2eNi9RFfWMMTpfdcqgY8vZXrQeEFrCN8LwPTfilfZ7fQRwb22eFBHeRu5nTBgpH/Z9VaChGWcIb
qpBO+NVNFZFqst26gevQhnRBvNGMifCzWYL9agDMyPu2cndaeviXm5Rm301C9Ae3mAiZWURSMZFW
3OWAjFhB6MO4knhtBSlE3E4kkODSzmOz0Ffi3KHAEhJb9+ys+bhzxLbuWse0tWPSVjYcBoaAT3on
EpmxzpkrFeMgdJ0Ls7TIS+kdy775Sft/DzvRtYFKlc0Mf2KUezeSRshBZz/EXniB09HQOPdSnmDC
mukdEM/9HLe9tqMe4Xjdl5wTiix7LD5el63mXFBZSSi9gsy6PmFUqpcOpx3z5Fto3U0BLjl+i2Cb
ezMeqqeC5WPy86Zy7TySEIf4djjoAnAh8rIDN+rrkY8oGxxGPC60Q63HEB9qVe7Gjkzmw49ySWit
5bBS5pCOPNGKaQeX+KlFSo2/hore34ejgs3jfSOZAXHCCAWQC2m3Oqu6mYaF9mncCpedGQ7pe7eD
43wNXDcArGCFOp/llHMoh5bnv1wx0Gjt+PK2wtxdJu852W8MBDOq0CR3o5kkecCGIGGBLOxUVXm0
A2qzqAzBSQsNtGv+AyGAPHTBbiF+aikI5N9YMr2xVLcj5tdtbY3dcpQc/2kE1iWpfjMz5rMwM046
/33mOyNiJYQ2SLx/9dwLPklFq14SQfcljj0w1E5LbjtI5DdJ/8Z8At3Tax+5q2S+QGrVD7WuCy7U
jULi4xZ0h1wWbckVTUgY/CAZGo8htVaFQc//KdWmqdxA9saKLHZaePH87LoPkXRrfHo1vLM7iy7A
Wnbcij0gyi0nbLRvYxeMN5RuMM5qFcqQK74GlChweudmoOnXhI6k7BlQsRopDC9/r0CkSVUkIkmv
525DP3UFmjAVa42D88HXSsOAgoLXK17YhZde/1Zz/5UDvtrQ1MhebVk2k467V0w85XK2gH5wyoRx
iIHOj0bL8V8ynviQqkzbGFHmMfbmCLzgRckvEtMiGn5L1HkFFQiqoL4cF9Op0WqbYK3nOX7y1xZS
WXUvsnG6AwiOl3FJ1T1KXXCBdu0z+3kp0GseHqLIXEyV2w5hazsYhjv+X9t8CAm+GP1dkU4wGMna
gjAxxAwPZJp9z8AM0cUz4FkQZ2iPRYCPfa47Whaa7VCX1YvALuJ6XCRaVUKU5qtp7b1LOlRCTeVw
6sDgv/lPTZ7WfoQziqgvtKPGXzmiAqZ9uPR/lx5LmeyxPbdAUOH8R7B3ITPKHdPFHwrTQEDajbQa
6vzxdR3t7DWC12mvCD8kHdOQnMEbWN7HtEAJ03ooG1VaSYs3PkYOnec30d+ADgD47dOkn8GCElXF
XGT8wjc7T1C1YXbfFvenXWjRhwKMihHNPzrURPzG6XDCAws0auKTR7+ckl/Xf3tCpaZAco8akVR5
mpMvwdwsDvkVKnvkRoet37MtabWFfIfsWTyu9qqT3KmyGL+BAxe6f2H8Sv7R7dkN6GEJNkTQHMUi
khvQmQO9Upuap2KfztiMruKe5MgvgnNbuSiS1LxgeOqI/uYavxVJBq4NFlzob/+hj0g/rAL5uedB
pt1TeeZmuRf6BbEOABeASLMuNMLGaeQj8KBXoWuSZOO3NL+o/REYGFn+d5pT/eYww18CAUwckWh6
QfVI7iIPZNjsAyGYE2CitaWPZwjsDLzPt88HqjH+i+rNyuOUDp6fM3Yd9MDwhB2ban9iBA82h7eo
M1VIf705m9DrnqTKHkX30MArPzMFUNByzCgI9N0ufPppOz4D9GITuBhftGf3hRBcSH85tJw79UHT
xQGL8X55vxe5rEJClYizMAEHiON/UuceqXA/sQpI2hPUyDiU4LzfQRm65b+G549/ira3zdiLR6cj
vtwxvQFztY0zTA6IiiglrXQvMKKnNizPjsgtaW4D8dkkqr+Hzgd+F3kLc0bcuz3dcjbdH3U7Garw
CReWuwFnYUDlsDLLV+VzoUJqujWkPGYt+BiCXmmWkeAn5yzwCAZseYkYVnkVH5hxLB+AoWNh3Ww0
GnZ9saLm5KG1UoblXdSek1IszxPRorQu9SBGieQb4qv3yfT76vd6q0Tk+IGaxzNXD7fe9gtJXYn7
WenfFQliG/uCZri+QT5g4IhP3kRe8u3VvgUl/2um+WD0nSwEz2CafOZO4w0TkNHwGQKn/Bo5YBqS
yjGYVCtcgJ7I86KKQd/JfhkD6APStXB1M2jVY/MWO+ABpQAEIBu6X8gvBvPlqBoRKBJK/bXxVVUU
MC4HqBewZh7DVdsRL2peH9G51Iyy31ZON9n7+S+c9vphWHYEhNaSxRhxtdvqiSkLqnpwyWMb3SbK
FuxbuLIAZKFG/lnjwX5ehp7UOuIECzOIQV1b2UQ5MtkgLPcBQr2edg5WQIzL6mpBpR9kWzNYi4+V
ENr5qxYqJbHXCctPWKebGteGUm3BlYVh6OJ+v3sFM0baWwzKuu7Hij7AXE05snFNpG0e3lc1Eflu
3UfMbaI4jgBZ5q5Dj8idvYyH4IwQvsuR/5ajTOd4tu9W25maHzU5e70D7sXlSMxjrKOwn2KtUqf2
Agha2+3+Gfcs7CH1DvwSRU6HurlXyv6h9LvFGmavoduuIZKpaE03qgxZgn94/6z8dgR1rPweRXwf
SEz/qYO9Rgdi2LsH7161RtLN0IxOxD03gnC9xLKeLkWKHgq4Unbdn5Cpo8XO6AtT3jvPozuca9ht
urJO3JG+WMtGDlFzDHAg7qRtPU8LsxVrIe2mJvpGcF0jQVk8+aJM57azGvCdDIe4psIDMt/12mf5
IaP2EgNAQEOdl/ffp6AI8nnDRQRLILKwDb72Lman2ysYwP2Fs19pIsRI2QH24cYwiut3CKhX1irE
5ZQeqWa+3LkrGXy93XEjA4gT9/P1h/43h9r0NGZkYdZxqJbnal+qab7w+TtfyOkafpWPMyOJrVnx
IafKP4g6G+XTzn17VUFmw0bPug6Yx9Gm9cX5WVWbJLy90ORPg2ZhN4oK62sK/P90AecyrdnCgiIX
nZUDPQQVkrOjKo4VNf/2LDWwbr4CIGkeovdPPk07cC+jzHAnfi/kkGqSII4qa3eqMPJEtP/zgiEf
gmy4feq6jOGG98STjIKKhKPqvT2u5MRonRyONoiEi3KUoIGpDLdn0PyWjTXvG6kSo52jsJX4cKv0
FCLqWUFnO4joWJUtfPdHTZnhsA2zSotYExfISmmcCWAMdJvCtbTGG3UY6ZZcLGoxxxBuLPI7O4nf
GyV29R5o4ZDLyf67Kp+s046S0wPF7F50Im+tyZXyyuhJjZ35WpC10u3QVnj6LfueUHae0HLHPsmf
XGOWKAoOAxPqaJgZXGRBdMq2/6aswmjBi28TkPUflEn2BlLZ7KLTj2Cq0MbJKKYzlB+gomMCDryx
lDm3uGdJw904z9Vj+8ivC8eaGjxLn+TmHr2g1hlcMbBg401cY/aobvCAplXsdjhUJfCEegHrA3rc
2VhF5tcjVcKOfgkc0GXA6XJNV9Y1AgpblgbqzHrIeHU7qLETQxP3EhnOMg0sKE65MIEXzEtEAefc
ZBu4iA0vkMCn1pPf7FU0BcnRTOhiPXqxQLmTt45mW8Y/K7l7IF9hr7ABOuJ6xglGRehV3MfPVv+O
GcaE5VhXx42UaBW0qRclJzqw5CWQKPl8+BsG1teRjU+RG0DOrWyrjy5ZCK7qMFhxci0/e/hZocVj
w5Z7RUnYA7lh9cemT210G7BZiHKQu0+LNqL5nqRKMLIUp0o+B5MHE8dbjzlRNMpPUJBv1skU1pET
dRlaDtrhAD7aLbXOzA0R97g2yKFSN0Zu+WlGu/8+abnUwzfKSSHM0TBaDN1ZDVvxU3zD+50teW/1
SRm5X6wrUB49y+7p9C0byidkra72clGvovryZ0dohAltoAlfKmLvAXqUDJUMAIrAvi6k1IEGeRG4
DMz/6SnK74VkLlmw3cJah3VFj3o1DeK0eFJYBEEMJVXAh1ZZT2Fcr5AiLAasvVEnUS75J9RocHys
2JV3M107abEqR2KKnomu4g1HnY6kxJ71Dx9lozn66UGRUsc9nUNxiOUSchiUWc+CQhFlKzzmch82
Mes1wlo2ZwILRej//Svx+xnZ65FvLqbjq6PdtYXuqQ3SWLOKGR6wbERrmST9K/kRKrgBL8JZBmfA
qxdJ6DLJwIWd24L7mueRZIyRN9js4mY/cfLW+RsUiKR5yz3Sexnaxg59K2vJfDKC5Y2x/3Wda72d
jO7mqaHuiWFAOOVzLZmkpPZY5Y+mBQGmJhQ2tgnIDao3bde6slrsuTyTqjKIoxbMqY22AXhEn0te
cyc+slEK6VwK08N44JnNuV8/riE3vnb0G7G+4je2k1pX72SEgiZoS3TYegqPoxKypG1FtDFy1RNh
L2FDacCxC4u/VhWmls9TDTrB9pywNj0VxZJEU57yUdaasw2H2XzpLYfds2xcYDmr4+DOaXIElG+q
yYvW6a7/PUh/G38/eL4Rb55EmzS/8itYOyN0sEf7JODY6gXUqduXX+2KnLx4vpddLnL5tn2kSnfM
hzYIvGRivDqhxYR9Jzaq6YrN4iGhx0NfFpGGdXcsWxbYqAWfl6CCQKWgRQBkfbL1m16Kp7gkAL5F
ddSnP2lOavdaCK2I1cEyn1+JO0SDLo+gwJxOkYraWLfTF801CpLrBX2bAvCPiuTN98W6+nSBmoH+
WEprmBtlYaVBtuKrC6gMG2XXaJGHYk4MUIAqvJHyTDeygdGEJyQPgBNefOFXsFcpATFWrk6Y/cIy
GnyKwqctdvSyz6cZDMm93uW/4JAlW3xbbLPFGn7aO16Yib46btS7g3RH0WnWrBUacTjX176H+jow
ovo9vnKXqtZmBrheNx4kdtL42RmGTU0UgK8GPjnqy9kBBbLs9FHKZvjTuQYm1JPQZYY5yWb+vnbn
5uKU3gT5GnzOzeGlQWtmAwM0CNKR/vptinMgL/X/28SEIJ92fZyjL7hU4ryskFvmZpjScDRQ3VQc
DSPraRYGel21i7o4KyUldG72fMBDnM7+FCTXbd02cXvMNgp5ZZ+86QK1xdLiPSGGDJo1ERPiC8S3
xrs3wuJ9+58bjiFBlC5gSWBVIEBrek30PSbP0NEQ/rtE4lsqi1+nXQ76A/Uf3C2s7zgg23rpt2F8
aRJcravB2O5isYnrJsJriwMqQGmYI7rmdrWKrDTVXT8vaHDDT0/3Li+mM2Ek13fIxBT3a+kPTN6o
c2CfzxJz8uWFDa3UpWjyQDpBuVHRDMg6TajBTDF+PGNK8R7/uJW3/K2/9/4a+g/+xr8kwwnf6RmX
op117TVdwvUc3y13k7q3aNkbpXGxduVXx66Q9tQEYC9H1ZSd1VZuXZcKKOxqttbLAjqterfzlXZf
T5ftmwJzzz+uKzl4ab5Wh8JwHGUnOn3PexPeIJRx4vLmvheH58org5VzTRKDPCKmO35CgTL/FxDb
c+JF+NRs1HjbHjYif8rK9IzIgbB8YHn7ldrDS+KYeK3a/0GtCTVSRagZ7yR33J1HhmtsQLTCqMi2
mRR+d7CIQ/PAFo27adjE9eqmyGyyPuAoYnmop199+2u6d4+EdqRTPehukmmsihbQewTE1A8yEcfM
bJpWjd7Dc9LH7FzzywMHKXiBDBKgYVdOBEcysIVJRivcjv8COVPEeRSOMV278qp+znm6PdAjewbg
u3XVQu3BKho4gz004FDaVLgDTYp8J4ZG7Kx59qYC7wnwIfs6k5taPXCQaUjD6uj8ZprupB5iyfN6
3naL/CTMc0T/qZcokZT1gB4qx/Qayr4gPcQc5T8y89w61l6WvOgogLS0Gw5fYOnUzpGeM0W50xqU
a1K7y+jdC5BHMDB/xgJaqlNB55jfRsnZEiSBy3miDx7xH2q4KBm1vD2x/4xinUJchehnRvzpGovK
HrpXfm4Hz0qIPHIpewmHtx3B3h9YzWmvKZ+8l2hqFhsy8XjlhPWYfo9b+2GzinicbpsLppS0Qybw
wV7sUzSxygLoQ8JhDlGN9MhqH8nKKeIaVi7AVI4+31VKf3+bc01QbjnxeVEp7giNf9l7c2Vl/81r
fm4FD5DPRHaZE9qmbrLXoC2ROltygP1wQCb4K4/z+kV75TyISHWg5yCe0zX+ItO3FSA6YNA3O5Z9
UZ0lLunto65XSsBO6QRwnET3tb2ppGhgzRw1CLxNy1dOZ1StjKmmTMrx5OUEtvpIR+9KlHPoE8p7
nc6uDWgWHeQNS9v4U8hh7BB4qGDRSWggyqkGO+bKF/O47dwHkV6xfEkKlzhR4dBPZmLs8wpsKL4V
VYPA29tq5NLVPGxPtc/XL/3ga2OSFCD0yZpFubAmsJRBoXnn2wHdRqTHzP4auRMx7MmCpjcMk+lm
F7JirUKq+/nEHIELjo+S4uVSnq8T1LY0ALvckHyd8XzuYN78VV5aQufn1BkJksdHFbYul3b0ofjk
KYI8pLsVWUGf3Q4P2qCAyj3aeuBPsXnROPtiYwHtAS15EzompF6Y+iZCmemTsR6ni9ezjEKfs7OV
YsZgUZhU6FOKmEDF0aYbLQvELg8SSIzKX+8KgUZxNwiqwcRPpD5vCC5xZ+yygQ8JA4Wz/FidkiZN
x8OC8PlVPPxbiioJ7c/0xEsUiO+4YbR6JXmxK3sL9FEdYxIMcQjTMXI6kjDihiXPQzp+l/vUE5GO
Eh48oB6KwR5D2bL/Nc6I3eJ/ghRQGv5D37c19/UIO3ECo4OIAXLjJmhGejJebXLxwwvnUFIcXmcR
gQxTx78pqzsPKpfFIpYBeXsHUfzvwJL/mSiQlf/voPnAJN8uZgcxB7R0vo3TKMN4sQwkK84uGGRv
fgJ+7OvunU2rHn/r5Zn2KNOmEdn+pJAI6jzcDzFplqrGUMp77FsOMA5lSk5D/g9dBN8/cA3idWb2
EqjqswVwk/lOpVevo+5HODt0Tb1Bha3t2VZjcJkPLapbr/Fs1sTI+JrG9g8/Ovb1OSijLt76wC/w
2m57a0Fthcb9lBcTjZN/3zTdgQ7sfqKWuIhTUadUepOw6l4ACkU16u78RE9GdE2D9w3YVLfE2A+C
zJb+XrEChqFTpQo4eGoVp2sCKZ3YaolJvcG9zaedsA5+MyR/MP40fp0ksZVOU4otUleZduU4S566
n9r/haEgvdyDCZN9QdEnBAAB6xIo52CxA5LHOAJ+hawVmTILDWBZoGX8tMY1m5X5KdAXvW6vklla
bxJyVDsvtIJn7FZAyuDOrIeQMYPURce94C/RwdJGn/EmJOC6K6NurgG3JfOU7xg9LzNW31lWUoqp
N5OPaVQ/eN0nip2ecdbpnLVISf4OHFpIz70rT+K0Eo1QW4OB77/IYpgktUQAFPLh6OLZlawaDZ21
qYwRivS6Ydn0jzdN1jqgeW/oJd4A+Ce26tsgp8YlKhy9MylaMT7pkLGTA30O8/wpTS18PdZ533eN
75rLK7fB1oQ1Zg79GOYKDZ2G6zyeORgbJuNpadmM7ObqY/dqf4L9E69u8zlchbvJinlk+u31HaaO
pY7CdQtG5aU4PXjYwb1m4VfhCVw5meP4HXgOM23XmQg+cMuGAYmyMsk9Yeihf4jaMljwHaWyhQIw
jkfu4mdF9GNpdXylsAe1wZ/Fbj09zx6OyixzOMW4HS/APSupcaqGUSya5TvIePm9zjpYJdoSUydH
WTGzjk6GL2iRG4aTJMSxXkJktdUugxHl8jr00gQKVkEGdGltUAh1tjEzWVfbpVgJofhgrcM+pMWW
5bBfzoyYDVv7SUEhH+ns2fyDhziqSKH6CqRoYenX2AM3udx57L86GhLZcpGJWQtzJc//SAuaW1MU
v/A3/3G1rgMWXP4gv4GCIs8XoP7b1Fj5jJqMfBb57QnCpDFp19t7jLQPMkR/wKxqCzuWjOOr2AOP
8qMycdR2KxkKi70TsqVi6FRKRKvYldPef1P/UjBuGbw9QPTTjhLX4PfrQCiupLDQGXTFJvFwkiC/
mGPuuSlotKP1SznDbar/LN87MhuK7ya0VT5/TW1c+XXejM6M94ZtxbFOA6G4VfC2s109dRBlpaR7
v7rqdsSIzEPa8hqZ+5lNddM8jCW5XQfb4X8ZybdpT1EdnhNTHzehMrQ1/4A0v6JvuO2Hsdz52wyl
xF3DXqjtMBurqlVZ+Ah6vf6x7gsdfvJtH8ouueAshNuMAyWIWt4qE93BD5VtuZmCxbbxQ9iTM3B4
I0jdPK+bBn6RKz1tmXShv8eRjCIvVtFXV4Wx6oia0V9LuHhkqeR2IqFh+SMC1lNz/GGEtWhMyCNF
WK4826niG/UtoXWhkF9arhJTCr7HYK/zckAB4I4rUDh8Ylr/ht4heENR7Ejm/P0TamX+134ONwIR
AnJ/8RhWHl0Kfs3x4EEZf3IA9w4NQ2wH/KqFBj1NkWvgvRa4zd/IS9Bx3Prgq4cY6A7G2LKJzDKH
Ztg46UqR5EwQwd52iRwD8RlpZdEgiBI6sHBrrFvf2EMITNHRvi10gX5VaFUFnDOJZza1AjRtMGY1
DBrIA5VXGxpjTWHM2F893lK2+ooNkxB90fruw3nzGxPXfkojPzJI4Cx/yXu5EpM3/SJMcpOrxP9P
wdyTZo32wQRXVLWrgKN9B8e78pvnFFt1l+72joDi81Z/tDlu3H/1nAPGDKfVAOH7XtUfkeoE/VCw
qgAtV+sW/zm0vTjlnW1gwpMHQ5u9Ej2LZ6YEV4B0grf/JgSC43qZz1MyemjePZOmzbj/ytTsTVDx
Ov68UASgRLWPKsdj+phpCVP8ILyFuxIeEfjCQ8M/5cbXQ2pFClTVY5ORmDnsJWp68g7HRVtfpOgt
5hvr2wuLlX+fkdSjrYwh3H0iKYtvnNdmMwDDrPjhYcBF9JJuK/d/Gn1bKVRdgtqH4qbCheQXJI4C
vVKMiYkyxPJFIomyNQa+eKPkSN9s1P6gxdDrL9VlXAHhRlY1ikl4z+ZizbPRnTSI2KYEYZyEPaYi
HQMY/qA8Y7zAJg+4kg/Zhb+FDeLfAuFWdeMnfsq+q9/Q68SEebXAk50LiABWz/CjaRAaF+dJD/Wc
A5syRpahJdGejqDC3TyzLmcl0FS+kPRbQRfTv2q0mCnUQ6sz4Spi8PNmP7vsIlJjZPzi37gpJEBh
nTOXydXq7ztWpE72J7JjCMR8Ic4PITwhC4tzhyOu3Ik/dDs6MFzmH+LcLgaPiJT+mz1cABSDh3zS
TgID5IwYqbxGh6Bm3ipys+eC7cnya677JLJU4Qf+5jRIomkyClJKbRmVMj6knOze9hxasjXIKX8W
UfXATSYeFaf2P/n0kTn1jCgs93P28plV2YDBqqoGvcaT9O7UJGaFds8eaBiz3ZZ6Vi8HLVawOTNv
okyAx34IL6yeG89YuVDaFmmAjdvkLV6py8KNTddaJoeKdlFTt3QKPKUhbS49B5B6M1HgP9OQ81Ms
2Jfd3TsHrsVZe6tR2fkVbqkprSmsYJVYU2pD2kW+2eTK7uYm2rt6bbfA4JvhBssONbM1zkg0be87
Th1+SWGkeG+l/TVDDW9bdMKwbdETtf5bOGV896ySk9Blbbr9uByd4OwKvXN0fCzpEiYRuy0SWztP
reuydNdWeVy7W/7bL3OTSLpk2DzztdmwLFMC4WapJW/qcOz2nSs6cuajchFHBGumMVz5p/rf5e7N
0KLxTdUMbnHEIqmElOMtw+J9B+DBzbDJkxKpYPUTDlO7/XKHAe23SU9uIJM4clpLQhcp/obn/tc8
T9gi+H0MAjqPIYPBJcAy1qpVeHMq+IMAhKuQT1Ywzo2l+o2BMTLHGeqGrDRYPCRG9YOv6qOqHYtX
d2c5PR524PXkaCYAIK2wOruY6MtKuwKxWFtOZ4UtADsMhxI9WlNEkwcTz7OIyygA9at2x5A+Llok
cST6dXzJy6wvxit7TKYtSu8zGDiuLg9ePBwyhRLjKNMWVc3Evl1Rq39lf8fzkuR8HT+iMqSpcCqn
wumdQ31JKXIiF6J4k9k/pp9gWQZuVJ2VFobSPbWKXfhO9TEsu6BKm4+G4QjS+v4pH7glSLx4rFL0
1SZynI0R965KN9rBsVQr1hyUuJ0agL5ppO0rNHAN4hCxyHoFVXv8bsuYx9nAd4rWSRTK0Bz+zLhC
32FuU2P4G2VN9gk7L4G8QMWQ8VxjlZRUrbuTDZsbMmlkwrSgpMVu6C2FzxlIf8yQikpaNyeLueL1
5BxDen7SQutOlXSEpm0/ZwoYz79uZ6XAGqE1MLmAacmbfsPLVgZX8hu6Ey7CdAkD6BGih8r0ONLf
9CUW6geE310Ng0AaeARR8xTmFWtXDBh8WBe0uuQsekbept9DilJOUfLB9l3cbY6yJoSP40DjH/7y
xNoVqo/SdFXgwPq4fbygbYx4DP8hihQDG6n8pNYfhAAnCy0GDJYt51JgFs9A8pKp/yki0TBZUsUv
8VYuLmRXucudqxW9smp0qhCFQHufbWZyNJfkcOsNfE2NnpFGRnEVqSFOzI/RyPlJxS9t4e86hC8u
YJ19/FBsjT9GLDQoxmOHN7SjfqYwW02ehoQCHie8hxbZYq5sEuQ7Z7MH2w1m22H2HnzREo/qvuUz
BWJ8BRctseGOMHzm8ObY2HdnWfu1/pR4flMO+kZLPOMEO+NJepilcrKFTux1LIAd3s//l/XvYTSu
8in9Hw+/ZonRyYuNNxP6EZL+YQjoRRHDKLXaFXWOEgO/srdG1Cihdp/RD7d851Mu5YiT5V6YVCYY
aMgNPYV2GGG310eCukZhjKWVIkDTVeQ4Yy7JCixv8p5WPFHE0xuITSJPHM+c+HQCes1cU5Mmx3aq
bjZfyl01FD7jYY97gUIQLh7B1lp6Qhk97VKQDSBmtgYvgRpKYLYi5M9ZmFzm2OsRXkyY790LNTqU
4xxjj3gR+mxd0+yItOMhG1TGX4tf4Yn+qNjsgaI9Mhz9UCDX4PHoe8mqrr7i4B0hfKUvidSHz8jw
VZceOZ69+1M2rWCOW6gvG5Tzi6VKuCcMbURf/KJ2oIXjli7fPJPHnpwZOvilw6e3LCSUO3kmFiVL
QnvZb1DSsaZkCGindmecLa6vgJDcjX9wWQMQHt821LPt/vd7Tfno5fdW+cBkO2K7mUC7ykMlC/wn
KGgDyBDHwYY1WqD3Ymh0UJ2vvOXLkjll18joqulXkDMsk0orovFCTBirMVj3YcsNMOYQ0x48GX3K
4zTG99klRci47gkhafxuABnikDeg79Ky5vmtvVMItzMxF1v7zQo/vLO6DlSdqb01q6XdXPQ69cj+
5EhpajNDNY1eozImyJ6+YxXEfgOBRdc6Tcc5mCR2iFKkHVqh+9htNzF+/b/XcK6yLwjCVygsGtul
KKeRDx7REVUxd9RGQOLzSWjtjd7OycEgp6UOU+eSFBuoKC+e475nOE1Xbf19guTD9DdbMp8sdNfm
5TvsCCg+I1IT2A47BwLFsqCcuRDa7hKQuZPT4BYoBV+KDftGnjE2DwhTOMhnApaUmAv8i1+J6CSm
z0hfzn7AysJUqofP+kNrnOe2HlwSVL5GC25aqkjoT/OtLR24az3KUDR+QUkg80+WenIMPgW1Vyes
A66GdsrxsClb5qL/qMOi73opF0JetM7IaTBBhaWSmwG5R1yScxXBjrxdnIOKssEhGG9bsm3bLYoF
xpA9JLcjfL7/u+GdjjVDj8JNG1/a0RicMMePIEq7Z67oHVvVG7H85Ct+1prXbeZXDBtTJcrqg6wh
Ac3xqPO1Jr4pc5OC+5Ae8agv/IbdbvIP/f1Kc2z5TVB39/vr7WStW6Jwop5W8hZ0it/hLrR6YzD1
5u6KLJUwad1hM9zefloQGyL8PZdAi0+t2JzzJ5KDHebLJpZIlIBBpLHQalCDtRr9S1tf1PGBc+CA
64nBQRKPm8IIztKGQTvNaHMRJmpi0necGf2gHFJDbbww9YivIUFUdeOcmpa8tTaQUx9i2lV7ESjJ
P6d4agJa4p+pel7xcuYmEEg4SoR0HSlpcn1NR48k6nkc2QcXfXZXleAbbCnhZj3VAxy2C2N3LMkc
FbNUTVraAhPDDubUV6xEs1IKPF5gyu0TlFIoytHQnmumqXaK45fQPkv3LkJnZJdq58cG4XIOHSuA
1RwUIe2z7ssN1BmWdxSTC1uYw54/8AUhtoZ8mPaU5Y9yITiTyF/vkKuFSVolkGy8LVYCZppdNq+f
AMNmbnytPJuw2cP5b2nzWydqCBFr9Tcv8QGhfsmGmJmC6lgcxrYKqntJw3YZuhfCpwT9vyCiPaVi
/WogRYO4lbQQjgk4aWqzB3DFlJHjkMcwLf4GLZ26g3zvaEFqKBD0ok8dAlf1f4aM+A/IEftTXnl1
gqfzi5bKsLVVlvfZ/tXDlVwOQ6vb+OUKk96EN5oQ7+ZvU0QbHMW5kZJ+R1bkkI0nLNG1FzVFis5L
9QRcEGGRdCQK8Qs0Iai5m1+MDP1jmMlmKJy0rix7+MqLX+E2nHAH7uocy8YFsybKha7gSBOQoeGp
KucScqoeZeXktBmxc+OFj8B//niUlGyBGUasU2UQmRBfdpPiXiGKCVj4j6VCYQWyXLKAQ/ZdPmpd
zXkC+8DyS0LYk2ONVbjaQYl8guWmYGGnPc3dUha1hVM5/EZ8p/9dOU61LeWLAsQCgIWdEo0c61JF
5qfUSPI2OY/su/CYtBqVxK873TIW4y7uikSyByqDXwif3MCrzZfDCo5sWOYDyIqut0VicDTMybSL
J/LVRcubACplHWAnSqEbjG4fH7BmQRM+sEpAfb1KrIgCNRr0A+EbbL3CEirnV/ZFRYQEds7/h8/c
fjudXcPhFBezFgu4Ms4LJg6Bf13HGqdRIDZNv1nDJEPQs85eky67CFYNQRTCxKI/uYEFAlNqjKBw
T16RG7nbztl+T6VMKZSgXr38WYg3MOFx+R333pkgUT6wFFECzZrkNncel6n45zWVnOBj5aCMEATe
JVrJ7fqQ/0/d1o2TIziVLnLCX93anmB1b0Zk3QxqrpCIpHboNH0pbmbMwigatOIYM+DAr5XEdVsw
KhVPHQ3M0zne3dCh0hyjrjz9tcuRua9epKJSoWixrA77jfin9sJHAofg3tnSViPCNslZh0QP4tjC
tYqmqeTiIK7iskQaFDrQwv06PrrUmNvpCvdhh5ixuexrm3AqDNSGFj5yzQScu42b7GuYHICBswHA
m4FVQ2c0XOC3OCN+fIzZbManUSk+mKpfLKon4z36QSSvFuK3e02nPss8wO2+l9om8hMXRNzSPpIE
JHsbDXaMPUe9LzO2cwX3A7+HCZpVzsD1ttCrHmyWmNvcY6RvGPZzsHBmBHxPTX/jd8oB5IogBksB
M0y8uoc84dgVk5s0+UibuOqHI7Dho242ev2kezgJ2LufsdXC/k6amZTBb8NG8PeIb8mLysXnsSfF
cZiCjP7yVdMMs5jfEAlhocCfn+vKBZJUQ3BgN1H4rL95ToES0ohsb7lzT5vxs1+u1dB1nVeeaL+w
by9twrJdfeGpFhNljf5VSP9coINsm6iKACV8Z6w1ATd9w1Y9kASUxkOn4KpIzAE3wGaQOqHRdQlr
9xMwZ3DWe9A2eMzvMqHdckVLCZ7Rva+KDNzt988o+ZuWlKPpxHg4IO/McT/nhRGiJjjK/YQLMjKO
WR0ujTVAubl+azPQ8h5F7YzzUimVj10G0LuQxA31B0/hKchwkD6FqYmKlXunPogHfazP3xUsy6+l
EfPYzZHLIKA3lvpyjl4PFkX06oLo0bHN7iJyEAKD8eI/usANXxP6TQVchAmzyD2vC7Sg5uyJJ4Wt
TwrTRpvgqm4vWOnYWHyJbCwyQPPZ20rBzVGE+aOo5xq4+ANuXwgtb6oj7Zy7i+1D4menCgfu0TR5
7rydPcww7Ky0aEEip+n30tFuI0iqQ9zk2QG4pxHKrF4WP+ShfOO19K1Q9cIX/AszNZZumoTE4myV
3NYVnKOp6Ba9C9NC/nKE1DQqbKlzivarAJWwwb5RqqNr2F9APv4x3sLeXE4MuCo95a2G5nEv1d4k
1WwVE2iVRWi9h5kUUvN8IAfxCdRNxaWLnpZBd6d3+tomD9yEPcpCD3cu1BP0QPipBgjEBBCLqgCH
YItP6xio/NOtrYUToKvQyFDqGRyr46+6e9YgCgXZxJnKfCMC0o6yLlXPhAwKLgCgHSLZpaWBMHqE
0DCiRKj1HfvIafirwaiv28My3B3ttIP62VMRxM0jPkllPDPysdhPKxk72eJJDlOIaYV5BPu98tY7
y9TA/cfu3YoTLpqlvqS2LW3iiatWwIvUsXg8V+b4ITPvswV0wsPdPpPwMLuN8Pzo03FTpSV0DYRT
kyRqtbBCMMPN48NaBc/3zw19e2lHHjCwFIOiA+wPuQugqEfbAecbu8GXglTRHxMLRZBSxzTTuEYT
0dHeZaCtwXiolKzJjyiDomnOlKTxSQWIhsCem3O7h2SKod4whlFCZ6kuxiJglFJxHx44LEeXOevF
PtFUCJcgTLjQaTmbWSxiwSIPmlb5ZkU3wdfmaSOwziZSiD69RvkverYUAMtSWM9MsBrlf2IlPZqG
aSTOx4dHarb7Y1H/XJo9glObcYiBMfxyX0x+VNiJr32/Waus5W7+vhGm9zL67SI7NTtcHtiyr/pE
vP86GfKAoeMtxhYkv+hV7SF4EMCTNu0/E+rgEPgaPDJndQXJ4MZgnAfver9+gHgS7yheDm3nCE1v
nfX4Fsj/16bU0IkjcGjEKli6BTnxZdHWuCsAAJ5fe31F8cLHD62hxR9VCMTpNPPbTFO0xM8h36mL
vVuTLUVJ6fTgLYSzcuWlJCplSU7Z5WQ7xs7NSLL3MPAa4/o6uhNg8f6a9T7N4bpWd2VC1S4HtmMQ
6xs0G51x3hfSsFNLRDH5PD712vYAJGxUql1mvXgGo5Nf0pAqJlp8L386fBy3c0gWrRVIWmbVo6kr
LoV5hFhtUB1e9GZLYqDdxu7d7rMJgVFjnty3Xc9E0CTKBGgPF+g6sP2OLrGZErEjEdUHTaikJ1vZ
E1CVn0N5B8dCb3rJbzCIbUzzpAaJQft20IR6zwVOWInTjYvjotY9N5GAPkMIrJ6XsJyV8qgJ9n7V
7lfcdoC75Y6q8r9ErOCrl/Ajrai9mZLXbQZH5HSu2FhaXWOTSHfm97ki7tdcIg0iyRbutji3fJ/3
ZS6B3hDwV0CLJBg+2XkxxoyKKMlCKt+dK1rz1nQMY87Ss9OOLd45AW+0KbR38ECGAF0Cde2WZ0ou
4kh1jOqsY9SKuVuQNtUFZ+QzVkzptkQwIfERl4PEE7nwXTYCZYbfaa3EEaH+LuZck9XfXbehWb5Z
65WPZiblRdXaNw80Yy13LGd7maFrMHO5D0n6gjZQ/nr2QchNusJ6SEyCDlwvZiqne1xzBjTJqgvN
XJLy0uALMTI44gLiANVrgW2bKAHZVHqIwoaKNEZ9//kzQ2LByRs/Efk2ZStx6JmLX7yPKzNg1j5i
7NVRiqtriplX1jkesjLuK8VaUFLbChhpuM2N3E2LZQV5mlMg/jbx8bvn62bLzNk7gGdyOkSLdEN+
5gA9bMy9/71tHrNP1My9vgDviTYMtVxs0Cbyij8lURPhM7Ehh8upnpiK2LKWY2kntimuR1/Km+3Y
ttCB/7gbwb0aUO9Tlwsem5LxmsrxRbQF0aohHZIKYYMWajYTk/S3aNgGKteTXrZBozQsvkkZIH7u
zEQSZPQnEeB1ocjID8D9rkV/sX4Ooi6cxk9pcJmFGaTgt9qMd7l/q8Lu+slLhStPlJSjb77ZZ9DJ
uxCmvqeMLsFn7Kj/umO03Z7vlBqhZAtCzKxjKbB83huOq85zRowIr25WzJgmdayqPeqZrjKmCkAB
xqdEDvhZitFUO70RkTci2Xz4riXMrWsZgNq7OUZ6cfsJ2GaUC7vhoXW9pCpf3kbqGWRrdXhd6FgA
jm6a+LFo4BzIk6xac3DyGk7Yd+fvyu9j/xwMkGbp4trrPDjQ1/PY5v6Xv1/TZ1pmmh1KU7wVp9qi
U3XwzO/oajpTisbvPYYOx7bw1tJDUiHA7LKVsgDzYZR6QYiOsr1W4nwW+YfxbT1HnCVZa280htlt
a4DSk6tynsiSpeyDp0se55Dt7PVJXIT3u5VqNHhNiF5bD8rR4gxMRaqGoaXg3xRQuqCh0ZbMgjVI
l8qkV7VEmboZd0NEbTSSj7cHWKmZOhixkrol3ly/k2UKAtxUH8WMqDmj9bR8PJfMD+gCFxfsed6j
I0MNxrwyGUo08TvJKvejFYG6MFBSVyYgR/Gd+Tp+SD/norHkUi5gmoZ1ghO68Bar+2dt4SGKsuV5
GjW1obXQJuDRRs1DOkr26UtySXHrvs9oVzB0f7mkeYkbqG2wWTae9sH13i+ewtUlwOm2uNcOiuUq
B7mERyrUzh80i71SEicjoZlQ+oxU11uiiOhil9+uwUyK/u+4KMGaO51kywpvg0q9rHAFIqFmTvQO
1xjzBEZ4YqbRNZZOr2yKnz05K/fjgARwICT1BiJEAgFp6l+naZq89KXeZJTB4ra1xVGzAkjZ1KM4
2ZWpuVxHljdVaUeLAoZQyCJ1NL0kBv+Vfsi6wT6f1rHiI0YQALfmPq64MIzJr9sBOHDlzvr646Ey
JvPBHsWUn0g1UJfvCpprk87Cl4Tt37CD119IEG0acnCdcNUZqEVSeYE69yXKzUL58mvBfo8pSl07
n/VGC3dzYlJoPZDObpvhYEh/IbXLAZP3j8fTWTc/cO+OaS3Kcex/qMxDrPHV8M5SZgvfQsOW3ar2
Uuk0TGIUNqyA7sNQwqXlUcJ7zc1BbApS2JZjSyjZeR8PgMFYkeFm+qzpnr8IegThjiDY+pXdvX9B
CC7SRO0ZLxSvXfKCTjBXUojpwt6/5X9YLOFI3HNThiFBel4e8ovo+bz1FhsdBWRydp25c0KI44T7
fCSsH4JGE0jct7gTIFw8eGYRBM0tWOHi7Ay3wFFYXG8u7JKoYO9hAp+U1UubOVcHG4IP1/h/KnZ7
fLUX0tR8RxXkLnzWwzXD6prz5dGvsgZbtORqQha2vE5CrgKnbg6mXElim2DErRjWA0aFn97vKyn4
vEscf7Vj+jxEAM4NbQAQEjajTe2rk/N49kgCkPtvp/2Z5/5JsiLXL3mUcNYyHVmkB3eOespbyhkw
8j3JLxzxgTzsNF2TfwYZv9F84hhCR+JSNUp9HiVp2l5YGTTSHUtW8MglV+RjkD+BzQeFv1oxZDEM
jG8xQZ04rEWz2+tm1eftEiYvNF+9ZVGNQDsUbVCknCN+sD3+tkKEdlEQKS+fmjPItDLpkj9au7FN
XfPXf5Fv0iMQOT6hRQxKAjNw+MaIALao923sf+STaQKVuI8i8nXDs7TvZxE+1jgPwvC/AgOv3voy
l4uaS+/ZeG3Y1JtL1PhSfK9ndXGoZ1bCGzFDxS72MbHU1Kp3NQ8dKJ4v0+AJG0vpgh41/jfTw+AU
Yh5oS+3YO+KIVuIIQzENEDC70/OEUR+XYR2luhv1zt1hgZuwRveJORUjLz74LSK9Mxfgh8TFmYdE
X4clSEE6rcBk6mHd+PBN3z+sSq4st4VPBJxx/j/wf3Ey9ZMIeJ+SLSHhS7vsvB347NuZUMxv5M1V
Q24LcNemOup4uF6DxTfByAzQb31pvmrc2m0FyX3RasjWP3ouPmUZi1XBhzu6BEqz+JhS5PeOMjhW
D3XPEhftg3I+9vnch/zKNxYMZV9Y/j8Hj2TxF0edmEvYtfGx5FpbFtq1ULptDPUc/PpIY4m+SOgH
VZGHeaGBpQwhiSaRqHBPQWywFsoWWCHQcYEojNSOwmaU4EhZBSsYDWQYbZOhkEPcMNCC2a6DrafC
0qwvW9Y3g01Q2gfL4EmWRqr/0MwnIYpWz0RwnhG39PSYxYnrDHul2eAZ3Nv60cpzdTuP9dXRO7yU
7GTKpevD2fhShvZWv1tGYJp5XYF/prA3K2b76NJtRVAmPILv3lyw3+WhXQJWdl9awWLZMvqAwif4
NseM0wUouV0PLQec87IZMz+zqf0b2OZ3F3H2gf95nCI3NqUGXXU+Ty2KqesqBT6BVfm83EZRbmeM
grQEEqfV8avSNxD3lV1Un63YtM5EmcdbHLyH+NLxPPuk1gXuJlMUEhzDHSMsrAi+AjGTQnxrch6L
v5WYStLHCOsx5eFiir9o5IwC1ixdTNbhljhoVfbE5MzKrfXu4YvHLnclF97b5p3QD+LI7Q+tBT4+
co+pt+pVBILYCd1qXvfkkeVhLM6inrIDPp5yg1O0wya2h1OjRaIv2Ld5A5jd4lOzDlEdQXTsPfIH
DzSpzAbuvyLu9IDdQcb7JpqyzzCS2QbMxYPUN2Jbpp/XPoq+Z/4UdoCMAHXaDeTfOiW2yuJtlYnu
M2cgxs1VXycImfUQL+DQTOLo6AcvWdv9lmgzekr8AMXGzwiuf98cNsEKYX8R7xPE1vBlPByAcP/4
h7vIb8pojmfNSzJI61elnCsn8NLo6219Ff055KNLj8leN3CIy6tWExtRXJqQh1MjqIln4tj47qYA
saUgQkloU/6P8cwQ/8pvyzupq8kl06q5Uma70u3rkMam0ISXADGwHaua13/seEg/rJaOCcEXEq6m
0sTfuYOJRhS9Ez4FCQAGJBPjxSX9aaNgFXymp97SfFCnlYqDhpbdeWpDC54mG9gw4PXu9fboS99Y
f9Vhwneto7IuZh++A2rwlh672DVDYAaON8WIzJmGKpkOhMGsBAx+Wk8w4hEuEDsAmckkf0KQ3zUs
fbj5ebs5CwaBn/ETGDzOkag4oNpUjB1nOBJpALI52p6OlDG1wgM+g9m8GffXwh3P2CmnkgdYejdE
N3yjngkVBYMG+Dl56Gx2Us8UeKLXBV4EIYY94CpJTcegcjDaANgtMmAozXdkNedjBhAoiyUb+lTT
1DJ9q1S5HirU32lhltrndkLvLiPeqApMd9vyzZmjA0yB+/QdvlpqMw477Tk0zAEFj0BZ3JC9e8EL
7uc13giqb5dgHETqGDIy2fQS3AN81UbPzzuon08R/AlTFLQbXql+hkzdv0c+bWpmsIeLeQxTUFnH
rNNMxpBwjwDhkrSPl5mTkIi/Oy/kdPxUuHWCG4aFV99ITSVXKqzAK78JblDKh43HjWaG3Bb7LyxP
olZACj5UbCluhHe6U708IDL9q6dI0gaq2gLykcbsiyTQDFeyUf/wqFhL88qe5t0G1qUT8s/3FEwF
F+DVMkVszsfpQ2BIb4K/h+P+QzSStWceV9dnx1FuUwQ7wCg3XbaPPH+RTDb7izhpocpvW2Ibip7k
BOHqhnUmv4dfqL/tgTSLeT0WYFWMewc5ps0V40QpAThKBzknSF7pikNPpwUn0NOHZ2b2dtftI237
z7ADfuMUV34XG0bJXwsG5R4UGzkAzTWGbsh2QCWwrGT4BYF+TvmNhSTgQyun1iJWWe5iRZlbQ0a0
oQqv3kbKwdAyqtVAPC/VkyCvM3h/jIZBWpGmayvwVltNUK6MVP61meW+dLgrqzo8hONHqAQM9CAx
0nEJQ7sguPvSaF+YpD0XjVhGZZMnuI4l+BmyLz7j95lW63mgQRPuzI8iiEKIqL1iBihDSCr2yABl
n2UTNf4U8AOKb+VfJL39wLa/BTq8xBawuSQjHXJ9/LkKFur1QrZsOPq83vE5VucRHp63BfLr9vgX
cOzWgNc7hA9IQhpswnsY3lt563x8X4IdzCJPyikluIC7Q864Defg9qJvEGBed9W8khwxkqc9fRZJ
IJ0tx1ThkRKaVrCoBdz8GVwwyFMPe+hXPcm62mxC/irh/a2FRqNR+kUHcrmK9YjjaHtSp2QMwksz
H64HLIjbWdCjDVyNfC8GBCdU4w2UMvVKSJAgr+nqvklPEgmsthsl1Tdz3WuM77UC0rXSMviLMR/e
/E9E4/6Bt25imu5Og4Szyt2S35iwwPfTIA96Mz8mkpSUlDu1WB/L2GxwdgDBrspaRCOGGSMl/e65
eCDNuzroU66T16Zy79Puki9P1UM4ONj9M++7/l5z3q2LyPGX6dd+lovxlaZ+OpnEXNovJt5Xy8w7
kDDgwtnkCoAOs1yvP66+xtPiK3DSrJAW4eAI+if0b3sShyMW/Hd31Hzz+b2DLmdBOV8wgHLfLDo+
1hKo5LcZCsnx1NFVG78Yj7nc1mk1dCsGf6ncSymc5KlirUKNbDZ5cdIU1u+hhsq3F/PQAMfaf2eI
9mdVyCblcUmv3FliQDf99cOhk6sxR68sIVP441Ewf/VhH/TeZKE6RPuKDLDSdfNB2izTBIIG0ni2
6kYME8eeMHhgE5V/k/pLk52KZMRs4hf/uA43l1LaqSEaPSwSDIt1Jnu2dNucU3LTtK7zb8UhAScX
HYg6hIbfxabE+3FNfbUqvHDCU7dqkyENI9Lj5nwIiAVzfSwlUh1g/nlz/LUMFZzYyacgIUciZzXE
vXonSEPPkyazVG2LVeYMAEQa45CZT6Ddlh1xuPxDeKLj/s54oWHrYixIMKsCWN+ZlmEc6VGsst79
w8f3J4Ibqz45W31E2V3/b0I5mspWas6ELXiW3+81mV6n6VGD6PmUEbXFoc8omQfHLoKeFjUTF+3g
u+8+IQSO0FFNoNdlCrzhyGrVIDNK0xWRlm94k9ii8NwgvI1ZYhIXFUWZLputXpNVhM9Goigy4E09
4M8vkwQZA64pudl0xjmnSjurU8K4lt0eF9QBAnYslLe8FKmTuLKFTYgI0wJY4N6NvFGttI+NJtWZ
jJ2vWzC3rDwdYLiJ59lPaL8HFIuojI5DcIArkEkbPHyhz76iexdT4gW9sNerXX3Ng8Hd0F0Vqg1y
Rsg+FZHfQLnwApjwAGKLHPJYXve+ySv2g66i9vZ/tMfqicNe2NV6xy62UD9nFlU+TaDIutLPp/uJ
lQUyzmBvkHANgQNEMUyxIhoQe0x+KiUJMqt9/pC2dRpL6nojiI/jCND0zBpaCISFHD6qIIxhq1SP
1yVpzhzgV+a7ADfgodFkcu12JjBhLfzPRXiJMiXn9tLN7GTmu3HmnzmNxOCR+t5ejjldixTaF/WP
mHIciECoZlk1DS3Sm4/oo6DxNvkADETvG4AjKKkRiJcpezyyFXfdoc1P/2ptsxjLbbKbzHATJZdH
1UjneOFSDQAPsSgtJ3LrcATxxJE2n/XLP2JglQo99DsKuIL05qYDUq64uDfdiRBMsJTh7wfTFfSi
0+tPrqyFGeoWp9mytLUNRxqviTD32NPrFXKEB/rhW3rkGWzAQXnVfQIwDop7jFmOBTWzJBc/EXgY
viWUt5GM7aD9DjFj1aSZaMJU/Uo1++aUZ/03niIV7YZltpbEIN5Dy98w6w32eVO6/UU63aw/35uF
0CGgl/lVgaTghy+cbwlKRGzSCGf9M9sPC4/N0nsJJ87vwc0H1PG6/7EvvbBmbYzKEhwsMSwqHoEn
QE0xq1l09ezEcLa7LunZ69ExUoOon0BRvphzYS7dhhhNHT0v6xeIdEWRBrFKM7MEZQ2DvLaJrYI4
Mey81LvoZZpXDR4WZb1j5iGzKksyAZaj6ojwXUj5hUp0yodsnk8GUSeRUwhOwxzlAYkxbo0mTphF
4wVv09vw7xb5HdicnVA+kOLlLLKB0SB/svRWMTnJvuzO3+EM2hBcnYStq98wQAodhzAptch8pGg5
/1Q90X0Hpxw2ATdiA8VpnnIrRqHT6ivVW8/ttT30E+s7Ps6NuxIifkSpTXxu3MdNJL+PiGTULWoj
Me4eHoQLzdLHeQBYHRX8I23YpZapOuKJ0XxiKmbUo9MRLKHH8ozcYAZPqB3o9l7UWl3k5LlFw4P0
vCDI71LMgect/qKh1nkPZFOiWpcLT/WbWiDrle/MvsB5lfiiQfTc4CG0SKpJBLzKdF4sz/Zbp6pT
Enoog80UFSaa4s8I2efpx4+GufGCuR9iM+Hh+aE6Y6xc3yRmlv1cMipyDtIuU2p/npz8PraoDzkV
xldaJqom2vq9I9TZWlnHePxietMp7Q3bMSgK/U9JrLQHxkUQNxcWMGZigVlSGgW3uZt3pjowf2be
7fMn9OKicSDDSSEbZ6fOkAcL1Bh+5n111BNIhiNsHueftsXT5vrWrEqkGDN+aH6gJBnzBDsjRBt6
9aOLWLIaVP0NNYezrPY2g8GFdQNeGfGXmNd7jNNTkkf1IddfqaEJdO/ux5YT6rFvPUEauRlwg866
LqZDXfqZrk+DqEqNieOTRWlv3R9QSHkJ+F4Btx5sIHKbEsMFv9iqSy96Lnry2E01siVAojDl+Qxw
VuzitM5liyHvwialY9P3g/PtB0rl7mDYyazxqwnqOC1XApHURlt83xuCPEBiwmriKCC/N9aJO3Yv
2gOi3/PwBBR8enZz28umVrvD/VX5faX5ouJA4PAHP5t4XuFjWph4KJgx3c1m+LS/SY68beqCQtLE
yOCs2VOKrblfEkdWJO3SjX20DK4+IAX8D0OYf5zIMtgtW8HVhSuJ+ak/p19Joy5hIfjJ0HlewWs4
O0lDAV6eEEAvehBuvHG/Gl+gHdd+J0xD0OUBC9gekxVaUZSLCpiA8FPQXIxTt9/PZnf4r2TS0BJo
qGFa71SJz3uYTcbBvvcvzYkGRe8RVYaNDARJH/HYMuiQ95SEDNEVpPjp2yjkFx/R4V2ERRWzDJd9
44oDFNUnB0Ph5Au5F/SRPA5x7raBnX/GC5e0L71Z1jj/dy0QfFFWyduA5fOZQrC82YQsD80lnKYc
4TC/DuLiYjXS3ELymlmaaTBs94Ji+oWGo592S2uaSFHT/T5QEkpey2UIpYkbvdvr3PI+y+U6A7ms
QtMsHCkscaYSggNiH+siuo9YqLICYm4PWjWjnopCvI8xkKTPtZ/t0wn5MM88+2HhA2MAeIglnz6P
hlv9NWhJy3p75z8zGH7EQuTf4vQeMAAd0Sqjdg0ofOgT08FqY4DCKOGQzYWL3JVOecQ82OucMjoc
auRsUK1bM/CmSIczTAJK6xAmaL7cvUiG6phLoz3ZauDi+kIyiuCnrBsEPQMuTNMshHIX71u5RCkW
bnGLrkkBvV5h6WOWamJpLFG/BtYmOMZx1OI+gNN3mC8lEvy5JVV7XSkDSs9j001UaXWbPWALvYVo
9ORraTBF7qfElX0VqYCQn8FJvcnpUQfH7xEgkVlWtVP6stOOCtVppjeNWo1Tw4aeVe0lnwRVXDto
CxqxDxu6HVczJ6pepAcSKvHz7Y5FGzqSgrUOm0Gij1TOP4+wQowTkEHK8BPUkeZjR/kplHNE4n4R
B6UvJ03iGWcReE1enYDGXHxvDLa8ojeUUO3+q6VeLKiIi+I6GwBIJ2J5Wf3nwEfIVhsuiD1JzNxg
O1BdQ7YMfWb+rusIj0N0SkVuNX9bltzDBKax8s5ny4xX1o0QytBAy8hRCEqLseK/bFXR1IDNUHQz
IfoXh4IrbKJ74EPNChXFTzY1zx15f6wKoYHWPfCzmyijzxsuuEfYIgw5DMrm6A4bMPKUTicJwz8X
CyipWV5sw6Lxjlq2VDL3x7NK4OW9exS7THKUgNmXL/NgEEN7w5hfbBp25xgNC1aBTftzQuzJt4WA
hIqFhSA7yhhVXjGZQqMZi8ElrVRH6abosmjh3zi8hJGD51U9K/AK2WTPI2MVRQwsYa9GDLq6ZiIy
eVEYVB6c/p37Gf+rr0rf8D7XHQyFyQHtYZYLRuhW2IEvP8s3io3DfGdk1QSzwlhmJ++hV3oVdnPx
OBXsMRRJjajnvzFHFj8BFW97AU11sIcjpwcBgsVg3NEMbIepJqhqfubavOBEOnnBlPxyBNYorBKP
ThcxvT+39Bt5qG9MejTUVRs/6kP6GONzUY+aiaCCaPMEzac46dlDtEN3eZ4GkNAoXG7Jj50nE5z2
A/jAxEszYSf9yK7dciS9j7UZGWuGjAPHjMeJG4SXqmhG/2jWYv0LDJdAUxznGP8Nh2ezp13oJkEt
UN/pTQh1ADmTcXxofzF96hhTece/PQEDHnEleTLEoBWXOkyL1qINTT4XV7p5o6QuUxs7WTiaVXd2
NuWNkjCwSs1OJFbhwgQ9l9SZDyIRa80cxF9yKVcC0Tb1nPwF+bkNA7F0UjVN19+VX1j5W6ojKOaM
zG676yW5LiMTGnhXH7ay6egzCXvq8CMV0+SFbfyg8Y2tjK7h9kZUv/qNIJAb06izbiYlNk3mA2d/
koooLG2ZbVtu0YNMQvbK7ZnB7dVdy8lGaCq68RQv1CV+RuvtGxdHrr4yAIn2scYgKBeUHwrQqSob
Ob//atqA7E8I8CytH+pWSK3ksWuuCBl1A7ZEgXEH950XUL5RjoBs2bBpg69b1VojT4hPEYqVb285
reWHARaGfnl5P9j3iw4c5WV3O6isqIE63169/8UMjLCe9BfKu5bmukooZwBbOq+k6hRR/XKJngfK
7TEpZHzyPftqReL1GqmaXoU774HjhYa3VW2xSm2d5HEZoQmYwUVYDHivjpVGqBLRdSYe+d0JstL+
NjBftYoT1BIe+PWykRCRVxZ3K5adMV5HwybrV3KMxma7Lq8mMZKWteZ8C5wvGUAWsgw8NER5Gdpx
6/1I/6doSa/VfF8f41lZ4L051zRQzm6+kl3j6PdS8EL0lFKgjY7sfmmC9b6rCLRFjfNIUbaX98j1
mVCRdutBfVrdYh+08YyGwt1O8Nq11z+0vEMDSY1ctp4UbJjduad/G5+pqGCBJ6RxuWz570FjSVXj
KR/10MVa2ejlhbDeFj+ISSp9DrC2ahRZVZs0AjXhNW0CRpN0SJeoPLciGfIv/wwYV1AzZJabccoA
JYN9+VTkv1DMGnmeGIw7oxN2ULq08UDXyjuwJNpoEf5N5bReAYOJFwb7UxFRVKL+Z6xYWNRFkSV2
E9Eoy00r0XDObnEhKccrlRT+JIz9W1awWOX8ogmEkpWaBjt1nB9RcgBPWFwt9vGZu5+BLlx+rUz+
TuEeX1Nqhw4lqqW7GWqOiil9C7WmQHRDhTumVf2v7Oiypr6KrrVyhVExz8aigUVLxNvSTCmRH3/r
P+5njOzCVh6+6YQKJ284fSp6eCRqyoTuAf06DUMPFzIxW8TJMfoYdJ/JCa8MI/8mu08OfhlzP+qD
LDuf96Zk0+J/9jbn4TBO2yTf2EuGXykC9ZMt3WLUZSdY+SXaEE6KPUYwMRtF7tdaR8QkKAIE89gD
I6q9riFidRxMRteH0WKnwMV5GQwTRr/hP519wtO3NDZyI1ufrGhYDKgD1CKovmrU9PiaQ8b1FL24
rg+ZPWRaFSs/2tCQshArfrd8tvUGFg6URe3xrQ0tjbi2btTaQUAjJWaLodZFkQOQrkKnN21lAScK
As9ZYd9FDNB+aicJuaCD1j9DMalR8GKtnv6rd/gjkGXxyf1KFgdOVtXKsRrqIxL+gS4eEC3Mlh9b
I7W2AO010tZkgrfxL0WoQEwgS7GhNSlEoLCSHhsuw83VjYHk2zdF8bw6qv8S4Cd4s0X0y1Lb+ZCG
vq9/XBACnZJuqnnXsWbooEMojkPy2QvInkIs9RsEd42VroXvfCm98DVbQXQoZGBoAMlxocrKcAjN
+NlyW3Nc/JP/RKfF7Zu3K9FrVVNCRTU7JkeTWn4IMsws2QZJRi46+O3rvf9s7q6/S0R1k/rzK3Rc
/bIe67FtN39mDiQiMdjpmXhraUtdghfltgHFNKour80Nub5urKa2ccrt4x64ku97ENruAdBuSBbn
5ka1eEcBxgh8dUQFViJpvgDronpPo4SAJrF354Gs6aSaKZ2HwjaxV04T4d6Bm+RbmJ+cVXsNJj4h
/BNrSXdwM6UMo3Apa86WvROaw6Vok1j61qQHMH2NwUOg7yqCKYFWOxafb9T93k+FiaX74Y+gsRvf
utodVnCv66eLhyMZSJj9mSWNh6y7NRlY51dw08tP3prTipowMoQqwNTVJEgxBgNP71Ja3MIdAo6o
j9h81WHdwh81Njk1oWWzCuve4A697tQm4csZ8118pkgOYPTuTufijzzOunMbp8rs4mWM5m+Xl78o
tZYNye+jq7ZHyOUhZDeoRvlOUHOWdmu7XzDttmvxxC5HpI2uzdEpBkZdT0isgYvqZbrYr9oryx/n
YlRjGOoMRucqh8kezli24ZfSZJiF1qYmIRMFZyqtIEUb3uTHXU8l0tPTx9/RrSkzhgjbfYOuQRIW
HOWoB3WH9z/65ZGNv71Qxw6NQnxCdbN2eM2TQ/JLGrl7fLMqyDyRkuhD+v5XgWilE86/TzGmZz2W
Viw4N/AjnaWW263PzuoW13dqvDhKIBXeex2iRwzNLS7ktBO5pK3Vz1W1CaFoKqUGljOxC8YOLnuc
c1UPf0l3kJNl9vTe+gIFv9tzjAyVR25eoTUdUlSiyYo6S0Pc+Jt2rtIFsSDuFnYlZLl0QkW2jpup
9dm3i+NSrVHsIcqEwf2jkEs0WWJqiFknX2vOOw9X5JdaVYxFSiv6MivqKusClAmZFRclchSk62lM
CHcXk3x8/dsYf5EVDoiDCE2ubjw4z/qACL3OgjafOyyjQAh5IppSgPYWcguafGftDU9+uFTG0V83
KMPBFLoLg/EbhSY3P+cysOAeppUu6e2bGnjj6KX6A253J8uGpfSql+Y8jn3NKbSAuZdR9nLi/yra
ezqeauMMuTuL86J4RLYtmU/P5YDV1WqjXg9Zampg7Kg7miVKpNJRSeMOsGSfv6x+IrrIOQdn+PSO
ZCTIApZlXWU0Bw6sDbEr6p73s27fl9FHKnd9ngolR2CdqJ8pBndfiwfNdZSYUIiLC4Q9IezAXrYt
syt2aY08nN01f7DF/7iOwphh3f1K0CsLowC9OZ0+UogMIk9jSXCxG3EYSQEmrqi500hUSNk5FSVo
CvSDqeJfBw9Nup5xTZPHoNJZ5RSK7khMiQDb/f9ibjdNHNvVVL3SZ2s4Q872OJve0G7RJPAyEDaS
1q1pep+uMyD+QLpaUb8tfgvhAJZfdpPfkLzuG+NJ0gHGbOiojWCF34eED/uE5tsDNtSlMuweYzyZ
OyF6hiEWhpS//vMvlvGVWzLcY0RT+IoER1JBFvh8ImhU69EVrHgPXCSTTD+CQe+nIvgqeD1vc5I4
9gC1FfwDSef8MAXqpvpX/zelFCTXKm9sgs6f5booNM5KXwttKIX0Atinqg+Xa8QhSL8d11IyVuqt
c18HbNVNoIakeCDvhlgiudqoKMwMkI1GrWZGQ/paO16VAPcLOgCXogcGjkuaaQMp4SAuGIqBg37f
AaP93Iyhw+cDHhjIxbX08L47c7fN88OzeSlroOP4coMfW0SFz63By/JgFVI2YLkuzSJSnfytgHfo
1+EP8yHzYLD/qK7MOp3DPeKStLdJ3xfyWviAINGKS8zBpWlPNbJNHylOof0rDdUtvl7DSYAgurM8
8he9BEEtLSuVU7/valQuCKmbVmEs/NRkcMyhRdk7f4KLBBZcsmJNeT8WWS3sYCdHU441jHBS9ahP
CXkXqpNhdP4s68Ve3nSUZAUnNV0UdwypxGTYND8zftAurH3d323tt4KrXSm13CfgAMbCUiOGjwBg
YgjCMbpQVVCl/cVBH8WJPZkWvRAc3jSBvEya+8KgWr7LlMNtrzmMj5JfeIxxWqLo8CIqNK+O7kyV
VXDng7qIKwTyv3nRXAwsw25gVu8jowvq/y5TLrgDJdhHncQmDS0oYjk3VXnWp46Nw/y1xvoEhT/C
GCADbK2CwdudTyS+A4o90Qy/en8UJFEjlqxj1IqPlzabRiYWFc2MAR0HlbGU217q/46E7Z5F3V9H
6UwlqCxZpiwWfSYXNMgoAjfK1neiLEbh0y8WTBysgU2hdJhPwnrJKu8WiaW36rZRssRYy8twGPmf
rZyi5H/v7nBCeCc/RVGWdkzhGBJmHaLc/H+qgKwQDSIHF91m38KqzJtIv87tZxFvw+e8djzKteln
AanAzgRAI7bre0VzaXZ5ZVYe/qucOiPHyRCUGoZns+CoPC4wzll1SM3vnT5Hs4H2zCuEmINTQZfi
qKWGAn3lnSLnjRMhT/L54eRb8rHX/OTryH4fGEOoCWkPJgB00FB0lFkY0RTbK22H5hclzilRGcIy
RgO5cIoqHJ/TtUU3xekmjRe7diTX+kd2YI9Wb6GdIN4brA3SQKOIKwqeKADRehWn9u8KrrVmfZnW
L402uh3MqDIR7JVhw2f9WRQ/zaYN+VRLeiCxiLcoG0Rth8VfxFlyUCYTYZTj+nLnF3cyVpca89QE
Hz5WCkadM8N2Kz5sGdHyZBx1+nYVRO6k30Xs9EEWIK3rF/YWdPr6h/+A/EKXeCH8camPWymHb5YX
oB8c/oQCoPw15UJncbm18SZValpWleRBXIDyQkkVAhrMlJE07KOynziMCMCtdrjWUgdPO6ngbgne
ulbebZ1O2xPX8kvt6WicTdicn5TkK2GHZf9uKcVpHxCDLsFl5Ceo2lq9IJINAzXCiyRVIXvf6wXd
lX0d9PU3DzY1EWtmsABAsdJS4cvaqbmMikG3wOwqlr3GXgtlOui9sMFcYicP4xJnhT6hJEZKLdav
U6e94v8Ud6peseHB5dt0m5mE0vLI8+ZHrjyC48DWUElKFeb439Y6tHNDo2/rIiJ0by6Ed731UwXG
tEdTRfnZNzzpEOjVTHDywoTxi5biUlKmZVTelnE1H9SKUc0H2bgyOUZ/OM3lZzsj4VkjQZhemLui
CB+4ajIkHIxQzWWLbItpXP0OVjD9duf45dtQkafUfWm+QPcU2RX0No6P335Ejn0oOMuWsdDWh4e1
QoD84wlq7Z5b9ydmk+cPmvrXbHLQwCTwFOr6VSYZ7tJSD94g+hG+NOp8mr4QUmz7aCKLsBFmmqph
LwZ9dZ/qgJtUn6z7I7G4qiBqPUau33+sc0ZUXDWlUdVldGcQXaN/rPEIuP7/EPQ+Ilz6F7OtNTZK
p/HcZQTUOuxYNznO1vFsOzQyvW4LOOZnOZkQBen/oTi2zM++YvJchiCxpd8WNXI79/174tWACHqO
N36AaAcHbPKv5PElocV1rNgQiLdLFe+/mjOngOoeTGfXjqaLTnIyFgl+/8srrOZSvsTIeuL6yJ6L
T/FgSPpi83UQrVMPji3iPNAfYD+2qOgvmLTaRiyVixTToyjdGwGx4N8v5IRfz8tEqb0z8UoPzWcW
aXpXiiz/N5AtxoOxj+qjXEMXQln82Llyo3b1+pL00X4Gf0epxBcxqeZwh5e5Cckt0K2SvLo6rmpg
/UwX86M+jWPSSuI9X0Zq7g0aDu+Y4L1+wB0YLvPngwILdLQiHXN03YijU6Bs9QAmJecyzf9iTShi
TGcTG8VEx8p3EwyqmLz1H9JwudNvOJDWWyGVYuBFIMAeaA95o5sgf22kyet3QxtZtPRq5YJ6FqAh
QFBk523lLpJMkckGoHncuaq0KKYUig0Zd8eV9YMTKkfCsjrcJ9S0+0waLLc/DsM5PJ36hb1xVotg
1faPTtbDT3Ea4akpWn9f1mcrCYkI3I+nIdLcZws4dfjti0YLGXThTiCZ8cs+Z/N7MMi2uoONEgcd
6IQ4fkHqsp7oWjaGpYBMh4gINkFHtXWZlZjeiFqgxg+JDLG8ARS+Cqg00L2Y/mcHQkKh3/fm4Q5i
Q7RjhMf02ZdeQdwJk4S/ECBLfz6SS/64/G/cv5ucNStp11LGF02VXnlCJG481JgLxeW93aIJny9+
78HfbG4+6IZRpJ0sZeqoSs3K8kSE7wIt0OFr6cTum05p7PgA7upWifJsiU/YHrX4B/FzcMN+wNuw
+kplLNJTULrYvAXeSvf7wUl1CsHQkUcNXqTEK3QgJw23Eof5J/trIVX3sX5RVp0+CAgpoywO+0gt
erMQAY57OSiR16hYNqTJ029xTs4b3wU+8KQr3whDXar6FP+6PmlfJngADWZWmkr9JI91e1jCIdsP
ecrnBjbdwAghwDnRtCQyrtnUCIx0QR6c0aBqqIorQpTb+iWyLdRgqq2W104Mf29ktsicdOGcMAsd
YDX04mV8uoy5J94nRChqesWfSFnVGeWc8vSMj5kt/mF9445hl/ZbQ3dzgYQQiCoYauSxj3fdWiab
S8IYrDi3g2MvkRljumMcJ70Pu979kUOpwYj5xtOuIi67KLysKkJkZxZLVbdswLVVQrMIldMl1NHW
HDbXFYECc7dQTrM+xGbGqgyFWyIkpqsEXQlG4sk5G8rKEI+acWM4Ccu8GXcD0JPWWebkwaAc2Pei
EK24++kZj5Rj3vYVGCNCQI0AIb3byE1O5O5c7FmeK+aI1R6nWNSmnD88Kf6Pad4fj6+pvlRXpzrV
dbZK7yT69xNOJ1waJgrSOtgDl4yVhNT/5qnKYCR4R7TIAZYpHv/IEhqh7FeIdETI6ST3x/ofZkTs
nVywky3hN3XQgmR25HkiUFDXI07tXMpNxu5szTEsuPpKTtHzAfFOxzcB4trCRO5WWX9ErZ+AcIz1
PGJfUVRxxZwvIATQFRVgSzE4EF1E2b2qT1+GQbtTK+avXSCAsUIBlNaF69mIcThaXUy4Uy0Wr68q
7qYYuN+iO1WzJleNObW8HYDgOcFANziGF3QLHHZG21Mhdh1dDookbuyTe/pM2qTUvyXKaP5Yq5kK
IDeJ0Ri2KTvf1ocxx7EnmP0Y8DuLKeTSqxM1cQjJp/a5MIQzzA6ouTNLdI2Ud15vS+zxjYWf1Vtc
xQ4q4RTvAABGsgwzuzxej88Q0xTeNslpSB7ZV5xN2jYt1qRjLAScCSSn0PuJBAfUXIl9eecrHfRR
8BPbQPwIbuY3aDFJziqxMBpQzLzxPz+jCkKumTBH7C8qaohGjn9tsmrWtgQYp7Nr3pyJ2ogcu+2V
DJLxvB1vZvR9aDKtR6b+FOsNrGZbHtGz2sNNaQIsu1WNUBxrF5+xKljnMuQMljD623Jq89h7R8N3
lvuI9K9FzXHpVHqqZY5toBwecjXewbwuNQlRsxbOtJYXH3b3HnhcD8cMs76wASsDQH0phTt+BURq
WrLfMeJqAsLRvykvc/BLVvJ+PQYOeyJJ+UVkXHap2VoKD8tYhj5I0wJvWIrl4F4XD3BcCvKuaUbc
VvDyNgAT3ifenABBG4Xo9UxOS9bIYyBzrV1/25+4h4upVLZPe+yaPyriv7iBO1Yz+/c4bR42KzM8
01MiE5OBrouf+axebshSndTx0508f9lZWhKmeL8za35UgUSitefKPetx7neI8QNFMgIf8lhUNjR+
dGPCsaWiT+IDDmpx1V+/T7S42DSDwoVZLJ7vURK6Qasw0QkFdm0mKWKlA/kbxL3H5BSAeT5sM9Au
vIwZs7TaI4sOuWRAtD8HqCPdpi+GG7apLmKPYVOXGPFoOF5gIGsmGaeFBkjAK7PLKjJoFEYRRJVx
EnMtUDE6XbGpYPFqKdDsNpqEgLwPh2tEk07LFfH36amOipwUP++qcIsc+V94CVuDTY4QkOLhlyLX
CY/1/qx+6MjqcTPmHHO8H/kvI52ejD/5yIB6HinTNw8QcsHyUeNYsI9JDlJMwe+RkKZwVmBcF0X8
T0fTlrDmWd1tdF9+zQOuwizurcnv+u8L/gIEMEb29Mgx0f09gPk4Uvus9hptge8ZTxLJ7BFqqetK
pR7ydxaOteBOsVgn5dkssHziI38xy5Vp+/61KjfrcY8M9iMSrG2QBlVbwTMt2Whk0DzIY/N7pR4M
XBHYIAYFbRjmpZXRcT35ji8FNE44Z7ZicLnZsifrnWRiufjMdtiJDXFglzAcWS/2xQHCDcPX6r0x
TqtshMO9hHnnkKIMV7ln2Pk++Jqc/+8oeMlrtaq0Nv3WBqZy+nQkMjdNlFLhA8SOBVW/U8AEvaib
L4FRpBLt4WAZ1580EYIIdWkGYmihwjSUPisnC4YsDufswpiGCSRTBn74GxWlwwCWwxkbgwR2m5xo
VdKwAfOeL+ZPv9l/Z1mt/9+Dldq44MBx7huKFa8NVV/VGdCNJhSOXhgcAtqO+3kNoJJXMfCxyKjG
D8tnxBhAv3+bHhlYFEy8PGmTMLWZXsp3UoJSSD+R5GhA1Qwn/8cTcWrRoq4VP7EqlVVIuFGr5hqn
ytnh9lHYiSuvoaIt19ey11kCzJbHYXnYQLf3GAnUT15zUfTiWsiyUUBBLN3hVCqjFgOWoylXVuzI
DK2mQzAXcChxcAp0+FL5GBwSklCrtAEdx8S1gc2XtWOHIQyZcmh4jOJr3V3kL9CYC8GsqKLKE/rt
YB69Qb1F4iTPL9n5ulgfv47B/Z8ZA8pYURBfND8Ap8jwrbWQH/qsENAFW4ThVfdb3vYfFbdb7Z2v
GYcSxvAFTQlFM9eHx2q8Qz/FBVbKfW3sKKq+GEy42DkOXw8h8xwbOuyXZ75cqD2O8eZTGfR5pOaX
NOn6PTD2dC+EJyueiqDhAZzEudnWORkK6oTkRY207CGM0faeGGgkv7l8V7MFqjBNNSv5703w0Peq
2L1OpcBI27jK9rlQCuJOtZTp9ey6yeYXv0pEnr3y3R7DUN82LTno0BTodemn0Cx3jDKDZL0LxNkB
XyP8zKbE0rv+7xGt3+Q3Pq+5Elbu6NNXo0uVt4wag+QWxatc9MRkyhGwE8q8JjxwXc2e2thp1J7J
K77/6J5++5jC8H8XLawFMZb8t4cnUm0MyebRFFQBA9bHWoHoHyOk9x55kvEdO2CfTdIbrESuDJP0
79BHLp7EyevwZwv032YV50dzVoscuw4JmxA7ZP3NRe9ny5Ec4SMzpENmn62WvNiGl9hDvRTa+Cgn
/3XAzhFlOVeGym9nkE4XqwBYX2aesO7b/6jraxsOlcGDOJ3XDTYWIzYdQ6aM5NSM59igqW+Lkc9r
pm2/37ShAYdRRGRVtLsPSVXtgdxFI/P8i+gILqTRcf4axPQxGRUMH3VZYuIeDzJQKl2s1U2RpHKx
n4p7ijpKi7KVRUJMMaC/mjFk+RWTbGRm9JeUdeCMTIhSPidpNpAc70r7Chc9PYwuIiwvMCWri2Zx
WDIwQqBiskkHDta/NZwwRaq1xFjHXvPOW+/3VkVXNvVtFxc4Yy8IfL5Qc/Ni48866DaZXzb/9D2C
R8LjelGTg/ka2Cq0cWfgXzaRVG0+dnr93KPegBTzj/c43+63ttH+xWAS0WVI1/5yc+XkYJnPHcl7
xb2WIOO+ds/NPzwgHbdwYywR4/wrJ+Km2pA2nX9b0Q4OdELS0476WEDAz2myVT4bWKeuComLYoaC
GYrxvVa7wts+NazNdVGwOj4qFJWvyUxzo3R83crkXbkBRIyratyBM5dZhKaPllOehro8OvUHWus8
JJ++06WXkLzhDK5oJYokalXXdSbxyUMQTB/SKOHCLPSe9YfceFFB7GYKh8qVVouVNayz1ewgI7cE
hk9BsI1xZ3qjBE4CiWu+hrbaJWLJqxntkA8BpTfVbZEh7oyp/w79OhjtDUxLCh0oZKZTBGUfc95l
jSK3YEHfej+HB116urvH2IZID7zI716I/ToJlAq4aBqTkuxngu6W0p//NU+zv4fSpy1TftaIcuTK
2pxqnEJauO1SlCvZo15mdbvuMTK7mWpfbghb6g1LQIenMCxLvFzCnhGfgemj3TF21Fti/RVgAKYV
FyLR7SFz3eaXqOdHNqyNr7E8fXzx9cTGpJ44ZP7Wwy6wrHx6UroMmnqj4XwR2/aiaRbtMW+zXZ8H
gtk6aEK+Dvhw8m9CtrG/IAXlIisFfIrEehRbNlF9topmKcFA7g9vsc3Zs2Ckz8jJRvo+EJUKmVsr
oTj7HxsJz5ogC2iaeUKVURl8DhaEGxfveKjBTHmZ5p9stoIsZfnp286SoUWVI5pUrPCl25DXZKyu
+FTfLw6oqjb9wkE0NLK34oopg1W4gCu23S1HN5Gbq1647uYEUongk+93RWqh2w9SBl6rj1vQmu3l
oOBKlrkuMXgf2AgovPP6Lf0cx4NtzFsvs0+1vmLgar0a+aRxtgxWmjjfUD5XV6xq9d2MglGybSl6
vFLLrn6OoZ0rhFgrn4SSHb5m3cwpHslBlBPEHFfsK8iycw/uzVCjWw4cX9dU1IH/ILjQfHn71U2/
Rxx3y9h7NYPyti0i/E4ir/vy992gysl1kjKnrJ/kVJBnPwTUAdNidj1ED2XOnrygPbmEQz21Rsef
fLj5u4syWRVBrF9nHSGWmsUxFxgp9KE4WD/L8pe4ittJeeKzkVUOXYj2judN1BGKKXj4526DFsz7
qmhGAHZaIaZCxBIZSOyywSUL0iNXJA8XfGmayqaHe7G7DcPtgLIVeesuJTgXtKre6Rj1W7UdB+/d
qIIniWw2Hhe0d3XGNBGHI1XhbhRLpz1sdDuzyYytkJqrn8QGRevfusxyjpT85Gr3kGUoulLAqlcW
MFft+qYuN52xnfYo5FC7BguDsJuyhuN45nU8q8zZixx/HGv3cOtUPMjwAZxXngGb/j0WogFN3VOI
GUNTSDgW8/DgFrpyUbR+q+ZGDBJEi0trPyY4/0uRF3Ew/9uEZuYT+tSA7ftp4aE/MEdItMPAQ/9s
m0/K9S8NiyGQw52edS9Oyi2jKlOw3JB2UA5ayzSzBFmGAD8tz3GCZI6/kYkZZz88pgXaXmz8spBM
eybVTmkX3/5fZMf1vhiZBF8tBrIyfJYDdKUI/p6ZC4OI8k9kPkRi17OcIk0OZIFlAnRDewQrULAo
20zTyTt4n+l+HYALMWoYc/SzYAwwaRXChcrsEKr1KfNTJ2Dl2j6o0840P0lwjTYdJ4GeHHzA7W1Y
FmrBgWAt5g4YzuqUbE0K/F7dtyQ6nvcMJAYsNSwukVCZxL7j4QWvbdNhHuCRIYOjyWLsnAs+XY+i
RTZmAudtc/Tb0lKWvEcKO75+s0Ug1UUMBJoGSXNIfsgBCKZ/VFe7jVetFOrUP7GxdS/l9/HKUpLU
jaTqamHpkb8SBIK/qMZL9ilDcJ1nbtFzdJXiqiRqLyEOMw52niPWVbju6PiL0AgVgnUj7vp5hDpH
emUdneEopkCQi8Jtvc/8qjk9OQAZ+N5kXxtk7Ax9DYyrfcV+jn9FyZyepjStO9pnFGsiKI6syiis
sbvQL+FiVbsqU/GBV+6nTvizczDyXS2ACKcn3o69Yxw8GhBeks2VpJjvmqdBWNgXza91BDqZLqRM
w6u6HdmHI7ocJa5VFXvdqe356RhSTB4LvzLtyf2rWUuCKpq/xP+vZPZ3Jhgil4bWjpC8s7WWZPji
wdKWPRMAxXy/CZ7Rn1y+CuYxpfrfNTTvDMnnmsggl6kMcBP3PN35Yk6RitIRagVQ9jQRbMRRsNmZ
a7D0ASGo+Vbghmw6mmuu/IFMw65WNv/uiTnrcPF2cX7ZuEzEiAgAenRp/5uvEd2SWlgkAxvR5kNE
Mj59ZPUJVvFIOtNz16OrJ5LH/yN30YOMNN5KexKMhilE+RkNOZbPe5iKmXC2g742NXKpNdegmXdT
i1/qeZkcguCX4WhsbtzqKUoaHoq8MZgVfMaMs5DBBYUxiiE6B/SViRK3RIu8MertCH/tZp0jfIwR
RihDLIPY7PFKc932e8/6PRlgbo1WHKNzvF6ZgS/MjYLya/WYAfCY54uxW9F/TTKGBc30R6KD/08k
rBGpvxJhZnZ9Jx0Cpc8262EO6x7EJqBtFC7es12DYVVxEt6lWM+/Pw7as7G42r7szEVCiieAuAaF
sHVw5jIPgG0ELv3ToscOOw7ziO6ZnvgU7f2A+HVZKCkePPHj42w2NZx7mU0E8bZEM8/vtfvxiK3l
psvX4XwwnfIgOIxVY0BuBQUWkMgowiL09MVRWEcBc5yMXLT6AuKD57M2naHyAtfuT3jPP8R/+FN5
oAjEZmmt7jF7luJ8AfYqaCFaVdWYsHJqukMdBaK/SC5HkvCiaaUwiuN3nR0p3qyZNsZAhWy8ZkUl
B58KcIrkjChiPrrdyZljzMXbO49TfRX9xKdaKGYYjyuOCVLwZAA7b+TqTEtYC5AinOXB9NdZrNa4
FBI6zAm/tbypaosGNTRJ0qO54fTWuXnFPNP4nvaSUU+OOR72M4KsqScuCEMuKapNxF7y7uUiz6Am
VNItG1GiW6hcU/lUnOxt+C7eXM6+mz71vjNU/9J/1x8cMnTOYWoEiCqnOiycbBibOzGPg34JLguX
lG55crOlAVDujwfHOC834rPrXv4gXjKF5xTOBhqcz/HiESlbOgJKe3ExgiXbd6sJIX2m0NVRUCWl
x+7c/LXeWwaVf6AG5Ayy+5NNIA1bJTrthHdn+0OOrfaDs8qydQzz3cqubq3QFnTsX7tLPN10Hmlb
EPNhM8mO8SlIfvTY4L2d0C+oqZWxsH5DO4HTYJzExIz/oaO7ysB/Kj9EXjjWs7MAQguKSQYQYuU7
zzznfrGw6repZJ9ZdDaIf1sUIfAk6l+NzcihBcQt+u3Jj2arON3PkR1HUQTCqYalg0nsbMN48b8j
f1FADwQInF/S6wNvyoFwQWfWAQqLbeBISIqB6fyBXnaAR8BC8JISrTYcfoAgNgy4EcoVI1ej6pTB
DvAOAi0mv7XqM6fEvC9Jf7KSgnbZ5Kx6JsM1hHoowSj+/XP8gFEXWwAoxMTizQr1FqqQ7PeCZaGz
MwQFpX2s50x5Hd4DnEc23Vp0csqAD2WvYMivHCtpo5jmHaDd50stuNAonu+X4nYd5CUZBpO8UptW
FDztN8TITi8qMMxRajICzkgDzp9b68wiSjvVQ2uKXfJT2INErPX0uRsovkDgqnZuQrdzH1lmYXQS
eQiQm5VXy4cxxQXKCC1/n9AWxRFf0RE+AkaF670DxLqZMFt4MEnuwTtw7dNsfiupRgoShfr6uo6T
f863lFkiTH69qKXOgR3maaG7E7ZbQJ33pyUwjWUtJEtSW8cXjUtt/QslYqiDVJdgeOEgRQAT1aZ9
ff/42fIPgJCzieW+mRVUDupuyxOPu3p/334MYQPF9pE94ymJbABPInJr3qFAReHkr9A3Hh6ikGqA
Df7hzK6J8o8jEjWMGzX/2O5LJHkWUTP8iwIxM1bBnDOnLWjcEFf4bW56wQCwP39n+8BmIifg40pe
JIp+QL5/7NrADDtwc6bfc+JvYuX22IHC3afKLBANOMKsB0j53YKoit+UtIyC7iy96SEjFgK5Nvs+
jGqV0ifFixM6rFlN0t55glDFTXOzh0Lvk8xZxnJ14fL/wgWhU8cP2koALkm36B1YPXDrxrfBcSC+
LECPJhM0gm4kG3Z9QpX2Ek9zlLjr9CwHa5avEK0ZVZEzmNkBqd+mZs9pbOWffG13Ny/qsqtzhB0q
jyn9XbDbhsGiD1fETMD6IC2KyhLKLV+E/wmURJIO5arak94YlBD7nvOfPYfvRH0UnXrI/Ia+pnjx
tgsrNlMicrS6w9JMy6Qc7Z0e7PmeP9tCPmdIJTfEp+PGhVnsnNi5py3PznjN+V8xgkzp0kcHBZ4u
Zo0Zygedxrb3VvQzx/g47XZDoD0D+PtvmNs63S5tggKOBB1N6youKSacPrSW3KP6Fuagg2HOpIy8
2zbMHkfZfprMGO7DkojkvObBAMx92IPBeapK4Fq+9wcZZHuxug/27H4cmoIF+vPGNmx+4BpSVSTu
R20+aELGZCfcYKg1UKHb02DQ1XX2qQDn6li8edWbxpwb/7gR59rSNkQcldUqFh9oeGsXQCihU3Xb
w+TrI7xePmWN/SExIcZuiRsnJvn0R4mW6iJPrPCqc88GNpHIbwhpVGTYrPf5P5YUeghFXytDD0t1
8ZKywe+bbwoa2oNJJRyiLQjegApP3fMnyvkk7U5fxNCmLGQT7DbHCjjLjUfx4Nu6Kt2hx0dueWWn
baegrFsEh2Rec9sOTcbCbPCL5L2g27Dfmz/RUYNJOLAndKP4mpaikZ0WbeGhsPm4DcJ0F+wGwtqN
nWmpQEVrxNNEVJDzkjw8sUYoO6mg6rBwKf44OC3RFn5COLBTlFQtSvjuOwZWfpBL+T0QxVdlVnTi
ZtnIdRbpmydPjBXmoQY78LWPMFuLLLsOvUzRySMiICaz20JR66J5oQQYQmoJYo/DK1QFqp/sjMJ7
20Gmp95IW0sqgvlGTmnmWOAy9o2RkqMI19O+5WuUVPgP/cSjJuu4MJp6WuBvn9bv70f98DXaBxHU
4UQAJwstgd0rlM5oxy0PSi0aYlxMrr7lbbb42sZjiB9iPrDfIFUyzXGz51hTLSW6T7aV76Z9wZBE
hVwPeFfNtneUynDVACb+QORV7xNlHq+zVOqi9qWmw0hptgNueAEvd2w25yNVdzJ999jKqoyk4aXc
RHhslAJtqB8Yav3RO6RxcTjp4KQ590OgBhYq2AQGU05Nb4oJZOKmt6IhE7nJkAqKjqo2t9Z8ilfA
1V0Hir5QVZzbLCW6x+mJGDD1z4/HbROv//NJCsJqqNPlN8vAgiTszR2FFJ5hOvIeqa9ME8HHGG8T
LF2yZXgfprKKQxsaKozz1uHthdRzT0WPFaUW5XZ+KKFi8WMQ9TKA91hIL1BdbcgvrdDuY9UnnLKR
NNlK9ZMcFk5ggJAjZdyEyWQ1Da1Jf1N+t2bU3Ezo9dEzPa406yehdyWnVl+kgH+oylKd+EiecKCh
Uwp3yJtpLyrO97t+sDDUUMReQwD07CZurIAu06dTB7YzPp36Utl77+BibpVz4LLsovR1axbyhKij
wFqaclpROl7+WUM8J+bw1uk8pyP6qOeHg0bHSZpuo5vBGYtyOSQmzYfNaEBLHnr9iXAqvOpWIxrf
kerMSm4E4f7lANVgez6crC3meGl/lt+wceAYTP5kJp2lHsqY5alBApL1wZPSLaeZpEdNDmDadl8w
xYfU5E+jvj6h+6+VK2j8Sa4914iWVJ5Kbly7ayTcNk4eNoZ213eMhaE3AfNcTSXC3AKLRZ3Srgk7
WIYoKoaWOngZzdqO7RrYUKUXLJxJ0XFCOWbyeMyMLLd0m95IA1QuKxln0RMnSsv6gB6PFPB9Wais
OeK5ydFk+/ySPhWPlw/nQ3zs44cGx2Fx9WWxj82sdsjwx4JXyajjy41dZ1jI1jrtBZTSUSbFYUJY
5etsN3QTXkTaLCI4zpX/NwpyDZ+bUD98Tmd1BGZM74su5q123AFYiVzW9jolJI1lEsAfztwig0BB
1ufNWhGhVnTv4tRHrTtyZ6A0HfZBNPhLuruS4e0zNWpeRMyQvIh+4XbBFzZxzOvO9Er0GIAmCBFi
EOP/7hJsVxzQDMRltlG7s+GJUl/SpO8Ts/0j7VmuJpQ5bM5cxj+yN+Obd4MWn2ATBP8qYF9PseTe
QZkTiVKxZj1WpYi6siGMcry7Oh/MXWbex3ajZoEYNdRCAjCMDri8jn71MePc+daSHHYj1fLFdJ6i
Ih3ewGYiHLAhK+bcJZ6qvP8Xp1PInB9GLDsYoJoY6DkzyIJ5GTsnPY5xc7rdM4tuDoFUItEkMWgL
1M4t8nevbfRO5HeLsr96zrR8NDCD1ikU82vDEHFJOcKxIsUyKsBXWkKmFkFp97AskoGQfPW5HJsG
W2lO07tZlnRpTuXP3QNXnrKpZGjhxnYp/CISpZXHyDtNeMJuehQHSM9XLhQyC/49np9Wj4ykAImO
ytq6DliXMVGnAM1DO3Wd7w0hEH6LiugFmL60WpaiM++lwStnCt1jc2NloL5t0aO3YZEo9/FQZgdC
9KbfRF0lok8GVEjAK45b9s/hoaF7FQNlaeBILmdnI19TP0D8qLUXLVvE6HzvTAbWgskUCuBdTZbX
/J0mZRwJf6rOa66iLIwJmmQSfuWFVk31i8mWDpewlzdEIwhpTbsi2sIQ7TDyBTfBEC+8tc+ZJi2l
jnvW9wou97utnTT/vE2tKNH1TTaUKKmmeimkozPk2sMyYAn7Z8bSuPhOYpwp23+tbN0WeuQy+ck9
YlpwK0BBI9GvhlunrfMOlorXDr1CXEpeIXx0+M2tyBM4nINdyroDdd8XDYDUYT3LS+NxOG9VCtHV
0UhLactXmpzY+/8RgdNDFrsdV38y8dLWMXsnas6/xJTjhPeIz32CeCjqLxC+Tc19mZ/LRnqksW5l
JSnQB35pro0PX7h9XpLYV89nZezle5j5vuEvfK/55GfV/S+dkDO88sR0G5OrNF9g1fRtuct+AlV3
xD+i0Wnxk+gNWzJ573RfllOh/6xbfBg/39/ogCSNnpEoJhTeRyjasqwsMwmnylUGqPkRPHAxawVA
RPR91YvYtY6PZ1DEBBZtBNVqr2hv82h2c2Kkh4nVM8bYXKGDOZiKg5Qg3bnKBXioqlNFK9Xhqtrl
WIsS/vLyLlPnz1zOjim8aDIEfVBd7sbIyHFX/VCy7VETOIKjo1E7qqTdX+xRoCzUr6sntKTDqXYN
cFG2FLhJLbBFtS/6luCLz6R1BwjMOo4QSM0HHLdTlwjtLOHvccDdS+td4DMDvQw2gE2qGQdMsFoQ
TBb1Yaf5tUcueDIAgUD4U6jwNEto17gGeTbp+vc+EUA8n1TYsWixnvRAqbin8C5fpbxpF3Wf3tYP
7N0e7ngeouS9SgrWC7BrTc8iAnIHtKN09X7uEkPwwGJ/Nd/DDY+fREK8NeA6De/oLOr3L/gu16uC
OtA8uHcgC1294NR1iFt2xmAO6Mt0iRtd6l9j3VkMKjmhxuIKSXBPw62TnhizfFz/c72emlXgYCbK
f/gfVeNLk+StZjDvd+/7RR/MlC3avupmegQ0DhIN4meRXgHjqAUiIkqyVopEKYbVO5feG2p4B2GH
1+sIfx9z8M6I9ILd0a9o7dFPeKpAaa9zBZ8iLFYvCb/lBxOYYxGZSDfE+XVZcXYRarIdYOaufPxW
/eR8kcee72r+Egesp5aUW0itCGdGhUcfud3sum2/9PaDaaajFUlyCs6IAAG5KtkEBvYgTIvBMFyF
hMQKvO1EWJnO2Lyux3Jn2rQrM3GXgLPRln9nv3aNOGfjVIfiRROTBZfOhDpSNQlyB6hGbFqVxlv+
vnLRjqqi+Uu88ckxixQuOY6Du3gtPAmNQP0nFYZlHnFHSKwlXBkn4K7Aesn8/5ZVBNLy5M9RuIre
R+vwsQlYtbTEhSWnkA/OBVyxaKtlmFnyL5RpkC4ecnqelg5JV7uCfh2XIJ4UDB5TjnxT8nPxm4yb
nHSaYi4qDNJAgxLkqGf9E3R5y9SgmHrLXv0qAyoDTjuRv3eZPXLbaNaLbcps1V6fzjCDwJwr4c/L
fWTmm6tI8SrMTUmVJ/WQmthJ1f/ULQDvtiLkE//9o890Sp9Ev7zHVwPyJd1Io2uxr5ladiHBs1Yh
sEpUYEERwL2DSbR66kub2eNSJP9to3cxXfW/CvHc/MEVc+Ij9v5TEmTWcqER1pfkJ3ohHovoLd07
B8yBNsjMxdkR2bmegy3YuRn5l6tbV82ktKYPT5xDFe/sR7YHZkp+5o/VwcBGO+biiWNn/Zy1BCU2
72lKiOAxObfBER/T09VOW8cdk4LR6d5nHfvxI+gzSTzLzUshNRNgfNEQ/RLFGH7zcQiSjAmJ9CNb
Ld8xZxWgZyp8OawetgWLdEnfHKgRzE6/FbgPA9Gi7zPAgpZbODWziqBml6iMp1TkznPRM1hBDWq+
YCYMRz+qSJvBKdbBdGenF6IA74SiHjX5ngcY2B4roj6HxCNS5f6HdLwvlhOlFcKqIssKwmdLMCe5
f2kt6SQXtIVFSwMOZMRUbhMPUCWpuyt9o9wWtC6KtdK8vGRIZKAT+ZccZ35IrCy1rC6TN9ws6K9l
nNNk4CZc2faf38lAL22WC8tdJ3ePYOYasg1TT5u1BU96C3CPfVBOo06iKQpf/2buaM3xLcZF/NrX
skcG1zB0LD61jp4MCS9DWcGOPFZ6+58jmX9uCOwV5p0l7qH22df+Mn4O+v9rBD8vtf7VW6+ie8YI
DV/7yPv6bDT2H6a+UmwpVSbQewbPqnRPRx6Crj6R6n7O/DHPa4rgaLocKnnYXirFM0FxQswbhxsB
uYeEHwZhVJaVCwq4eOzuYgFf5wkE1As9FlatIDi5GF+ksyHbbwktBXu8tge1H78YGzGNmzDGy/VR
mZGSPvZmPIQ7kR8OYG5Gjfuhq5FrbAVagHQ0x6Yw8h2KlMogmqOZDKxM53LVpNQHuH8V5IJ9JNzM
+k3AakgMv1NVcWfB6/EjAOeEujdfqOQtAsdgm3Ro9SvLO9HA1hv+4Ju/FD5Hv3vxsylg3x5CJODL
9gmnvD6xS51YwG0m+FOXMggfBCysvs+Cq5kHztlAg43oLP3GYFujYfzSYJw7+o/Z/P5OOFv+sr8Q
HtpBzFtx3crmzwoXnqrf0d3a5seibQ3czH7wVQBSP/vLjlm5CaEr5oXfKEs+AlsS/ey0ZgceWuco
dGeziDBO9b47gkybX0ldg3Ck48fHCqtLepbPoJW7UdPPu7P7IQ6d//o7GjRZdg1QxskgYN9ilFHY
vwEPyLteh3S5dDkXOnWr0+8zuEDP1TZuLzDLQ7E6F/G8T99mETnij+ba9GOc5lJ+6fIH7IlWsn/p
pKMl5/wLy02Bz+MhmtDJ6M7ZpUcdkmNMiP+jbolx45nFGz0xyKWDF0dVASni5rCPJ7LiBUwrsObZ
8UOIlX1gSFGeqdftJQd1GA5gG2yyYrI+cZzkS3mKOGPir9GPEzlFcLQV0pweiIDWxU3YZdiyBIR0
TVhYTvWyhg6hQzZedAD7KSWR3Kyc4yK+UICFJBtgR1hSZXLjFZZNHdKdTD4DVWEJU9Zf85XFmcar
DSsQd/Hdy1/3yr5EJfAeMvG+LE1I9It/plGVvq11br6aHgH1bLA6QkU3ZaylTUROaes2/KJwPeTR
h7Uy+a0SQhWFhj73eVabkHZWpp7J1+3EosBTPo660b/PgoKKMV+t5d2unurnld3OyLGzbony6DlX
tiwFLRp6Osimc9uwE/Jf6w0KJMcP0iF5V+P0hdJDix7zhunlS2hDUvLcQHujuMah0At5Atel+rO5
EDPy1EgK/x9Ej9TsLvRpcJ1v28fEF7T40vq7+TMTsGDojRPde5EKIYw4sUF7WvITTmiX5wtQgzT8
B5QVKqQgvc+9oz1/qbvlRDXtVXanbtimGPq1WfXI9vyXHFz45U8Yb+ghjV6/ltXK2VuYKxKBxjr6
qyELoSAEF27EMiOe//Xh0gnRFqcDDH/ZQTMilJaPpg0DYlDooS57NLR8Vt5BwLQ/VtUGCZowgzM9
uNnXPhuNJOq1RFlLNBsWrOOI0xUPQig0fchyGVsvysgE8aDpA7FpmUXqkeavwb98FdSQ5zpmd/9k
J4I/AGsUTcIIBPOkQ91RGkDoNhxYbM5k00OKRfCvhw31Gn9pfAuP2ljhHwGIjpUPgYyyQEbVMlsw
H281e7iuyW7/8IgF5e/Ek49/GN0Dy8BQqIwzdBf6lsqB2jBn7d1Us0GPIzTa7LWHMMmh6Sy2ICwc
DfzwcSDHRI9IC2miBxcmLuB02+rBxRB6H7l1arp1M3yye3Lk9+5Uw7ZfZ1dF14Z82csn1BOwRxXq
9wRvECOhfiRtt/hL1aobYTdODP2Ae0W8cINODOOyt5S4KB7D1JE4UcLHIvpLxv6fMMBsHTxXP5BY
8CUJsYHOvX9OS7QD9Ef/nuLmvKWjvuHwMpqNMDACQQ81HJ1fAemr/Mif9zF0sYBQ3jklHsW0OrEq
iRYIM7lCyaDqTgF9AP8A7Fk9S6X7Ejhew7J5bvPMh4P/khtEVFj5MOF4Vq4KptliRQrNoU2GrTgy
SjXqRWD6DnM2poedaCV9+PXU4Tmbzu13X+nFLNfT0C0oaMuW5DpJDKGnvYhwnJyzKObuont7DkG7
KMI7uvyQzS5SFmoAl87M8xMVcq9dNrIiraZbLrM7byRjacAyecz7oTzddPm0OBu5LE5TymZHiom2
JLHTrshR/WApq6rxwXk9KEfQLesEvbvECdJ0m4lQ5x2mqzGfMxwF2bFJPYeuwkK3sY+gRpq4p1BI
gG0JRgXr3ncK+9UKz13Zk3CbGKk6bzpePCa3KVkEWFgJ556Mx8nlqRy7cwPpk4wzETGeAfbGIhwf
qr2ju0av+6q5zmrcqX68Zx/L8uboHWjqdqCcVJJdulDENeAzjfA7QlW2dZL6T6Gmmdftrkcf7XEY
zxDpym7YOhKBgjsApi7j4+e9bueyKB4CGkXH9t4YE94VAJ4sCeZCjWD+KJneQ+IrrJNh2fmj/ShP
hpQS1E+dXXWibBxcbV0ddeK2AjXkQGnMP4YA52Gk78W8BmjiPIOkMMwIRwwQ5O1pexNcq+NnIoim
9ptd4oxF4p7sCLY9GiIC4mSCGKJgfmtx/j3/NIOfYYBsNaA5KIRNbg9MJkG9QEpI3nT268WHWPm0
3vwRozLXLtGhQDZUqSWebviOdqVFSenHtPfbUiYyEx9iSMNjGClHMNxVKEFI4OcXjRRnBF4faa0Y
WOdMang3RXiraJIRuTmRz0kq7+dTnK/vuBEg7hzsY4M9pSE9QIb88Y0vI4gvHmikmAZuj6COawQ9
D7s+U0wdikXTZG5b59YccYHpusG8fM+sDkbND7sBdQvzF7+mGaXgGr8AmaZDOUtU39dTMsniZtdK
wktVVnjAHP2bAQDTF2/93fXCkGxRZvBz0WRXNlZnEu6HR2YiXTuLcHVQctwDi9qKhSv2EBlLNR+L
WidC8cnDmP7j98/lplP6skcrD7njABaiiMKIsK8C0K1IksPiUKfZFw79qum8PNnGAzgPcudSxzar
/ZpeotT6vqxdXfSFDn1qNcd53XUsR4X5Yw/sJYAm0Drbd3t2hs5K178qD3ekZlzhDt+0G7rtLUu4
CRTcXbNgVwtTYe8Ydo56hqtRKVUHWc/y7T0y/9cNLY6BSCd4nsC301ojb6mPnYjGC7DqA6VwE2Xj
uuLb2FawUa+awTqaLXmfnzUnTVmv1Re3eCQv/8u7l39HP9j8FEf+QoASgzffgc2+xtvVQRpntXnn
OSdO/pO7NiRvaPtLEDgCPjPrJ2Ru9viFv9ffMAw57yXYVpmySOoRVXLujg/sPEyRG9q6ggF7r6jr
SMEVVHxhqK3OeeDqb8AX+R2gq6aYayc1EWkzMS9QH4JN6/mRyoRwyBWi9i2WMOvWtEP22CG7Icvj
IDDkLESrM0p1yaHJujXcA5SHGejH4rnGij7N50/K8J3MFHuJWvIlUUPW7oV1nrxdloFnjEUbZxbT
a1vacxLNwHtU+Ze4elQTl+8sc0SXU6gyDtI+lrx2IcIm7xVYvT/K7iuwDqWCIfxKtO244VqG/DSF
oWrAwYA7DRnjWRBw/UMstKTJ3yAhd+j34h2QpobV0AKZm+88jdZsQuLD/uduvmJgCdDVeyxzey7i
PcfYm26mEf34zGFUbAhXK39p0ykTlsiLsflJf+lVVH0JaTQ5WU4mXmOvj2Y3uCHiaFy1akWV/AL/
tHuC7SqHedzYkvFB/Viy88rSLZ1XaLo5N+gBVV5Nz9yGTmyl23xNB+334RwJ27u2CASg/pra7vfn
N9a+Rd/52r/S430YpJYjo/TR4mkAdN1Sql56JNhm66TiGlzzEUO4oralSCk4MxmPeeQdFFYF4Gri
T/sKDdvJ4TOsaFU+iOne4jb19U3EQoe14rCtWd/LitW58bigLE0t5NQPn1XUDc4t9O1G/HyOuJ2r
UglZq1PyTXwxA1gv/DCc1TJVbFP+c1HNFPuMW8tQd1SdKAsGo4LXtpoZPwsGcOkAfn5qcHRXVANp
J+xNVftOT8D2kNRfgss9iondr6gUZZdWjislM+pDXc6IiSA0xo1VZnJ0LaEjDymzYL7lPSyrGj5u
fbZy7oP6/zbVliE10Fmg85UlzPGnAAKwgMGjze+RZZb4ng8PH9rKTSf+DoRQV+atpA5DrqHFq9Ws
8CM5JDaFC0nvkgH9ik3XyNBo/YV+de4oDT4uvwxQGBLc6CvZtSz/qZD3Sjqy3vSxc82dpGsY6mQD
/28dDV1Pz3XC59ZsHrYx7wnQdprw3WUPybYCDtdyFhutfrG48zr6DSWWDzpYgkQC/GkysKb8bq/q
InfCWHI9EM5lo8KnG06wV3oLiqpNoDPb6ZdPPJiCxJ/Z2YOP5f6b0+DnJkVfcDvytI3JurYZ98ip
XUJrzbx8LArBSs1/TyJIkNDbMaaCmNNR9j/zMPCIdNTVHP4hBA7XbFhHyNMSIa7LAGjVhWfAC2FL
QtU5UyZZ4ZWROoQid3Ak/7IEAuLyFL3C3JXvAds+e4U3FmC4XWmr/8kTLFt5heY2Gtw3sKfZXqbd
SlBPHwuNXY15wZ0j6Dgk4v/rDMyOrO5eRvH0RsW7aQzPREwXRcvI/m4KbWJFTboKW/qjNUh4Ji1n
BQPd8+aweBG6PNJBvB+g9cyszid8dIrY6eAxKkAicPz/lRB9ht/8XSolW2gRqkG2cxv0tARhHHyO
N3G/kcTD1lL5Tq47GAQ8CX+J3LM3SRcUxjj+nz1UgzAKehoAzG3Kez6ABGPIlkY3tBg4QvBzAETl
7PNWEviOZ3Owij1uNELCjacnXg1TVHvPXG8Qc6EvHhAHWsbjDk+vQYHUETL0RfT1rH2S1gwqqnlR
byvaDrZPf6fBlf9/yg1r15MSuW+Dvgj13Gp+BSAjLMApeiTIKXO2z0rUGZm/P5TsvwzLpaZ4Cf6c
3hb+KCX/1pxmFX1p3A+6b202j3XUdzGgALEWrm2dTxnrreXMmvUhvXnq51sn13JeX4RWsHzyC0yq
/5SttuxhSEkL3TmRRsaYFOHfo9TM7I2MzIukCdvXvWzv2huuvtVFtaxzlrQCx8u8qC8K1WdGe4aq
GgaZlVaSnEnAfpNBfOcfipgo/5M5FYD5GLmYa0Hp/fR1km38B2EfgVISPEO6aWqiqS+mq053Ycp7
OZNHZ1zBac3Yq/Sd7FEgA6G8198TBa5LhPqYwGpNNPJIpybHlsioM3XzLcoUsvXg6lcDuU7Mwrp/
yejkqjAJkLhpjF0/TdnPzFdqYmn4L3Uvo5lnv0Ie/Jyf11PAAMuZbT71qcxkbIhm8XgSbPx30+Ng
G+xAlxv5dPYObGFIUQJlzvHC4hbl6fJxKwPz+2Q/N1LrbdnG/89gTzAlAeBaILl9najhiwkA/wbQ
Qzu6QQt6emEqqH2wYc7G52bIOdMhkbRqzfOp1jAWb8zEHXOw7SkN0iId/1NHOxLIkv/MZcM8wRB7
pHnWGbtP68WVVf63G6fMxqlPJSLZeKHE3F3d47MrvtHpztNyanIDfv7a9Y3TyqUQ7Ah1xQVwUSOk
Qw9abj2xAm8K5uxsx/5c821t+pboql3Zta4++X+3KclmjHPuP5n6KCIdA0Gp9NUb0TwjqSO8+62N
chp1tXd9OJX/iSNzNip+kvvG2qchYwTZ6ilBynPFdqYC9zw/MQgW9AuiGt2sJyVI9Nzb22NIwQZM
h2ZWbIa15t9WGYGfl5v/OzNmSuSP9wZuU2xzDF2bXi1o1S31arzHlblNifVWhkYEV/tcH7TSn5BK
hqg8oBuMYR4/aXUdFOLX9wnvImABfs8lzWL2cVtfze5SqKmA5JN9G2T9upjTj+EuHQW6XMI2MmzC
88tOgRhosdotQCi8YkNBN5HkaSjZTpk/2hAcP7teCPgn2EBr5BQxPbqikifcmGpSgXun3HMd26nz
3OlgTlEyENDmGrqxUgPfQi7q0D1IzlXuP6DotPzIqAEPvjvX84nRmMU/DVzeG+RXq5dqpRBbGAXW
2muZG/i5AxHPWIdXPxPQzxHPJ3g5m6LD8O0+k/1hUeYNCIxwlm4nq6pTKqionq627/E2v0do3Vms
bN/5tMA5QLe1NNqSIYPHn218eZqRsFWrrNDrIvate/82UjFpCx9JbsmA0UqXvFVa0aOHQ5E9FTM2
bxLAID8j4FUa5ewN9bjcPqrnXCB3PteXtFSaLqqhx3wIY/m797a82ymL39+/tUwdaZvLe5gHavQg
Few+Q90s36sSusnmMO8oozyHCi6Ejy6SY10wHsied4fPCQ6eErCSfWlPGM8/imKBnG48xlqzjhHH
qU0WHOxkxr9t+f0nyJGcEPGLkEqfRlp8zt4EgSqc0WQ6kTCSbwcbTpR98EUVYvTpfjdCrdQWKTqZ
3BWtJt0B8eDC1LAk9CbmStTZqLyNNSMlM9sxHHCa0VRdG8xXSfLPqqiwaBGX7nt/vUA+SlhA1gTg
++p6yq5J9iU3OMxXAFHNNsKXWJt5JOo5ho1B/9rPB3e2aTKKuqZxxwfLCwDYcZlGSzW+Jk8gvl+w
F5Xl8LigwWWfPQLuDYrk83+FNl59Ke3ulTU3CHaIYVHsQ72hX45/1moxmfIjsG/PVwsFNayShIHG
K0aF7Jzfq/gpIFVuaTbXrBK3bIMMdJwxsWp2hxO95TYJyAQQQXHSYeNbDbj9PW0S+jGzuhVYfZXJ
TR47gDdgN9tSCcU5I+uJiHZTZDfkirelcV/z+JSk9Wb9ovicfXvZkPE/mQw7Jn0WmRMjfjCl0mzo
pVqs5j+QD5kHq3J4uOChkx6eQbSuQ1pVyWqhKLmcOhO7I0Asgu7DBA+qHAKISc6xsHvGs6S2FWHv
a+o63eJCZ7iM8LwnRAULMxaepFCtVTOkpUPhMeRQLQaDnqChRC87YQgvsmge5r9lMqPbiav5VjI+
T6EMkNw+1KKpNr5wTxr9iB3ikTsGUpkZLq03YGk8p83toZoEMCbGGeuqMAxJEE/CfsuiHj9H90Pn
271qbZVav+8xI2Ort8GSX7Aka48lqMRrhF0ogWBNDD+3WU6RRucNqvZMSOdHAydvdD0WCZ7/BIYg
tqUwn8/6DAX6IyXiErWakWyVuoAo7d2yir+/LUWmnn5roxcCRbYEldH/pft+OuBLnXYgFhn/UNHg
wFKFC1lLXjFKqPW+6VhSQ7Z8qNXB0vISUCcdqQ2DKxYZ6z3yIXQSvhwtZWr34jMO7IHOgsIbniHn
tjoo8yPH3HKpMu+Y878xraNqeJbP2zwViWQ2bTYQ+ds3T7+QMEVPR9T0gqJbCDVWf3YIobFkpPY9
uNZ6lkVETWzWTmHPqe9ZP0Iwc2f8xmut3BgHw3QbjjEX6ULewsFb1CP+6YI6ZSd0isI+hI9IJh0/
ms/sb3HBpcD0UpFUXL+iAdxMIAU+IlJfx5j9qbZDoyRNOkQ7Yz7HG25ExFlYHzhUVQeVwT9PCttC
xkecEMwhXGfVG843uw5qE6pES1LKDGdgAo8Km88ZKo91jLqtqlRfQLAz+83oq9WqprIXqyWv77SY
XUBNS1ckPIlMldqe8vd4OQrNxyRC4IFQA0ZbB/bAZhLfS9q22XzU3OMm4dedV4lUU2t51O8XIVB2
mLRA5V0laF1GNdHYrw5jLF+8wOqoVQ1/fZIUyZjCsF7WPZ9d09O9nLaqP+BMPebyA3xh+txaNP0W
/sUhm5nnAg+7zEl7bIC0XAZOUrDsKrhgrqnnr3aG8WBLxQjdTkJodlH9ZvputHxOgbcePqCasVkC
Orlz9RWyQh9YIpcJCnUSnXC2a8r0Ufj9CE2ICAs5/awG2p6BIqOpUgE4nKbnw8Oghcw38K3x41+i
qlSr4WKOS7h/9Qljf5bKdjgZfz886qh/P4loFmXF71jeUT79JILKp29SJlKG8z9bVosTlpYK0fLe
XMfrA/OcCy+72F874KSzOROCflBhpO0V1vmlbDKq8LdT1R9AYKFtni/UoYCGHUCdNwQBA5UkLnmt
SP1UIQajeQ5Ox3F5uE1t8jTtvXlgmBZRzT8ZpODnsvRu1m65FKgSBECYuELLXOrVBbzgnUcsPf5v
2VK/m3VlQGk8HAjTDq0mf4aod85WsWye7wb8y2TjN4syZsigv1At42Y4tALlwVTUd/oIbFu2vjBW
bmI64nfet0gGmLApojGWCqMF+uhoo39+ip6mAQDVIMBkXDHFB+B7IOJ4NtOxiuxjVr38lgzaY3QV
lSWIcJRyUz/QiHG25/sWnq0Oav+cz6UPPHvLOBzCiaW8vVlgTU9YaHQFeqDxv+1rvyFHvEJ4GZfy
SI8TSAVphDCS1SB1fZORunEvDbSSbXG2JFY1UHc9JqSh8blGckFY9yl7jqXgGKFcZeFNe/FReFG9
BNe+qEBfkD/s1nXJNVkqjs67dvIj0vqnIGFdFYOamRfvD9Ev+miuQC8sbNKfsCk7j810fOZjpTTd
F9mDngapcQO13JMYTAWxBbk1H6AAhpjO7IvWdnMk2EeKBalu1r3asRLuu1Q9W3xQQPrUS+Ui4Ckh
mGDUeCGr88uVMRzzYPulNiQjfY2YpHVJLIsMO3HcpFe4ZjQu/lKoOVks4bXxlOBODONbqhmMq2UH
pMxV4j1ix/mFdp8sJCBc5eEmjNdxVNND3bkq9rGpy2au//OAOej4gNiOyMO02VijKRbGAjtLTiSV
xueqg87WDCOOrgfuoktq7Fd4tuKB/FAOmrbJ25q/Qyf1yI0DPI78q5Fwo0fwOiMsg5uWP3UvwYDr
mb1pXooTnZ48ze5vepDwGhulriQMzPDxHiXacGAu4iiatCgkKXO+H+ex7U39gzgaw3SqiIsvmjJU
sIIe0bytwlLq+CnxAtjY8Ydl0KalvgVokH/XzA+TLoDqj2kac2OCEeitM7xdcr1PY1Q2jDgoKQ1n
bWuvrJZOk5+k8Cw77Yif84UmyJGOAmsmyDtAHpQte3xLdpdA8I54iVUG2ut88dOiQKlhdNAGcfKN
hOLcDZSIBUMzJ92Zv2LrieH3JfPrBYf2HafbOPpxEfMJrfkJRX+l04lvT8uxBvyh6gj2jNhuB+hi
R4Qpd0D5mkkQ2YeOZtE5YQUOBKblSRAjVDA7SIMZQTr2hNFSeszxLvSu7tyvmaiFs/KQx8JAJoFk
qqWNzUzDz+J1QItZXaRb49SFUe1vRrf7fI+KXD5+jF/u9Ie3Kyldeowhs6GerBANdfSoh/bWVlRW
h4rlyKPFXa4/1DNKxofKyW+kzfAqKEb36SNzPc35KBA3PWJRWR/Kbh70KmWYEaWlrPJXLbzmuZPs
Ecb2mXp4KrvBUVTZ1gyyHL2WdS+th5mf4280oZVespbtE+6vx8kHx+OqGWJQa+FwYFknLEbZuxyv
YH7v2jYfyK9j8DhFzh8+kEwtbK49N83wdBTKyb8Z31sM0Pc4UZEO4HgQR8+iyEUY/UFj2eCMgcjd
GiYs1tGvA3dbHrTXoljXoyGTGZgCIKHjNtG2fJ9wzm5+8SkXLb/4XJrXik69fKwB3DKRvBNXyAbJ
LtHDbHBEfkXQ0XEDacgXMbA2O2ng2Cdaw2w1nifPiUsNCHQCT/a5sZjjrtFhFvop85U0UbIIymkh
CCnzaZi+CulACmX3QrJjXJeyjpcKFC/jrgP3SZayL7TDBTjTPfvCLyyjnihUwJQGZiwgZz7cak9C
kSnS+EO5zCLyZ7lD5DHc32XToArpR8RX4XLTaWwOgUJtx4fggZVyF5QNLOS8WUvh9iJ0SYinwbyr
9E00jeBezA5vDMixN2+e8/Gxjf1dj17ftnXlXd36dGZOWIRL3Poy0Kccvi3xUXIobHK/Iff1ikRz
gA0kaq99bShkiTqFsBcW7Mh7G1aGYFNH/lCikWwW6NOWAXFLThDb80KME5xS57EcbDN14fayInvM
vjyGatGJr2fky5BnR7JFdZUgPrGHAB/T9SFPnnQCS+q8yLDoCVZtZs7yNixTDJI/798Nva7YDhMu
q8gZSQSaRIoT6jHTibcRtEOcNGfL/TM55taGfPbNx3fu5v99DMNqZq1DDF7+1FsbFoNlaMuSool9
tz0KYC8AjDKjDslBwO0/RriC+G3Ol7Z8mYtukorLCazMQQawT9p3HI8pNDlR2w/pJW0g6AB6WwYo
IkYtEksEcINra9O32S4nTrqXIZZX6ZU6AB9bjzOM4BrXO9D3ma02e0usCMjjF9zUonWNzM/fMIe0
dkSpuQMl+Yxk6n6CJyX/do/p9+W/VoegV0Tbz/nSR4SDKczh1h5cucX8miBca8nPkla0D00GjxYK
YnCd81YWjAKqo7BC3jbBvDegS1srpzDCm2EljNr8LvbQDMV7dW6+9Cz09K90Z/71q9MfiNraIa6t
exXdWW+c2o3Ms7o9B29wpLQ1ia609GBtAZ1ALOgFsSYWeXXeynj8vsWM+IGWaGAYkBEkCzACRxzZ
eew2qAe3oMRoUpaafNA/tOIf4k3aaAGun4bcEHHCL4ctMSKfIlYfXVRumcqOiMdB863rWlglcoZi
VGYryWVcrplWHaOT35ESEZqM2GV4uI9k0DFB5l5nh2Prrhi8wlqWUU3ON94Gi2ZmujblIz93zv6n
mOXhjDnqeByYgTnVzXiEbZg5X2he0PY1CW2W3DEFJEglycanuW+PH2VNE5Bc9v0GZE95iK1e/s4U
r6nnvXZIF4uJNLCoJ5N6OCljRAUrQdO/sOWtWRXL+K6TXMau8fpaVHFgGTEi8qPqwd/IklcxrCjd
ABXwGlVy10leMnkOMNH5aK+Bmf9bVLwjkdyTBkY6X2k5t9W+gOBuzECjLBZmf2nHiJh19XROrnf3
YVvYYvqTCvS5FolaNttq8gfWdO0UCpDZWNEdx+yRDrCaJM3Pg2yauu5fpg4k2iFINAM0SfU0n2vR
Vd5r9WHvGX70UCpYP7mKDR5DNsE13NTliEsqVfM/mbUouHOxw7VakZejZkpP/5PbRAVMeaxPU/r7
4gE6G4LF+ekBdNCKsctg23aGDeBOQrgG7oFVJUMlFX2htThQTfv2T9YvBP+CA1pKfIqrD6uDo3PR
O/ygxkSIAujOUp7+qNze/s4NeiUDRphPWuPI4myPqIHcDQ7cMPagqfe6Gm1N1IP2T7rjS69d9E5C
Cem8i5pgd3dtzVP7N1yONYtayNLZZ2mcQ54Lk9RCgm+yOBU+txSR7KJEKAU1pE9hpgB6LweZRfob
CPrfaG+OrzZFtmnRfnNgHxJArDuA0eD5EZBl+ZL5lzC2BjPRLV41/SuOxHvrtFWJwZjK3vgWQ8FE
RzoVgXWoE6vFpIp2agFogVblHBe/js/DFxnQ3L/3TrNu9rAraIbdeK5x/UJFxSWb54Zy0RsI6JFC
5G1gxTc5EFtazxxP6klUBHUbRaCHIH/SZKg6xLthxSdFK8Pct2oNNYp9ZLS6rdDyPPJYY1EqKm7G
/0lESdUty3wZHG1fsORgrWW83+vIrXHpFL+3wLbk/vhHT1D0l5PWw6H42nJEHy/448Zg/nX9YI/c
FY9UWnCcRJmVTr7RSKnkaJbMLgIXk0fLFv+mIOr7Pq1LnbmlLBDeiiAymdzl6bM4bF9PmXVZz2Ek
yYL5O9Fi2Nd90O91fDu5q5mdu2xdwErmvkROrsI20WqInfeUZ6i1HtBQTJrPs0tf+3SypBu8xfW+
ToNnv2ItlKzG1ZVxxs7Xq+j5jTz01LK307yBeylBH6BWz/btARKLrweNwyO2Wv2uHxwnq28/kRbr
/bdOqCvQtKHTEAnUXEqJNoE6JIM4+mX0Au0NmBKb6AlTdUbyu4WhzdyEPoe6gi4XPyrZ7kH0C4MK
q1kr4CQYroVgDc7v0YsJNzwe0I/c/GJh63yrPOFVmwzvnRIRpF2zTzAdZRHTmtt1fZVMN2tOI5ry
Z3yDg8oPxGuQsYf6Q89XrqjeTthC1iHUV6Aii5KqpEY5D6WpdDgW2lp1690Be4lBXmS71gSl3s13
IjlirZf1M9V6KSx81IuMKdx7Z9meVzuA8VyiVJTtWgfTzBFifEimFRxYKtRXhzvGt09mexW99ngW
yk0YPoL0bf0BtocZbJLHZnqJP9WTsGLONTaCjm/RxCZPoeCxuwM1NeSp9LfSgnrG7KgnKqNxygg4
3L5rgKpxYAQ1ICR/4RtSm8ZCzI91NqMPwvTz/2f/TPDSAdfIrUvgm5E9OBPjtSHtDm+Q+kscJsnz
kXjFOLzsXJL0ZCw3VdMBzUYD8x3/nQt4fYiDbLLuZidUvb27JA6xUYTevJP49c1ctJdGUlHIA6x8
Wcn22o9B9Q/sCtpYSHsgAIuFQLiHVqkl34v1qKBhwoZDrjZtX+a0XJVNEx1uVfHjFDsEy5tDbdRI
EgZAU84TSwO0P/x+teq0MN2tLlzZqaW9G9EyyWkkl+Byp3ge1t2vrCDTN+PRwEVBWquuw0Uq6omX
KMHC/4ZPgGP9iCW1IYbUIb53vRw4Qeiw2i6sDvBOgO1fKgJZ9z+5aLLc8vweHwcslHelSq6yqKdk
k16sBnjujl3vVK8lC6gQ6VzI2L/NCmGroQR91QM/re5kpa8NRnZJCujolqTk79gjsMqyqbqGPh61
7RcreFLAR7qWumzK2I7r1UoaLvopWI2/utM8k7JHsOKTulIiVJIV5xcZPOMhPrsdscgoRTUENV0J
zSRKdNryDVQGOB8CmxIj9AI9ZAtErA2zgoYW60uKbgfBUYaH65XzIFsqi83YkUtDbPyNcTQRm/nn
Pfaj+/lH7qUZKtnnWFsXRZM4iRBFJmJcsPjuCHuNuoXJRvak0SdQZ/bQZJ9gnhtxmQZ4wX7uAHu9
CutPr855KSRPGdmxwzIJjnQSbHwg6jIo/wmQ4mk676CZKdb41v0U3CdMhJMUoXsTtqSarBBGQfRw
+pPW4YStUWAn6qSdpfnZq/+p3n0u34GbRDR5OhO/976HBjMZOPKypsML5rRGajLq6jaXcJjrbKh0
nK0jsooqenf7+/KnJyTwxdqGUgenTOVCdm5sjlqM0dSjQwA/tmBuH4WTx2KIQesJALeRrlygAhfa
MxUTVog83b57rsVeVuuoPiknJLORu8i++sH3KNXb1rZw/RV89tNnL78FlJzWsSbgB6GeLJJiECGr
Kg2TSiuGE9ScHCtkqatmiXyWFrreIjzYLGtPp7r45Xgrbx+cxtquGBvv9Kkl9xag71NzM579bFGT
e7tdk4OmPVGwJlkAU7/EaOeQiaaZMI5qSfvmvuODzKpZATiU4Y0HZxasbRGWR3Um2s4JuCIvtoEG
809wMHt42LIqVYJpoBe4cLI5GK1fyqG0j7KD9nUIeDXXiHJnnCX+7attojikmEYIAT1+i8Qgo/B+
55yhmOPh8rz5yAHun2h61F9rMmwRDdzlx8CevRMtmdcFR23d4IcdYcT0TW3VbAv64B/imiym9CWK
Re02HviPXrZPDoAltHgS5aLhA+Qi/N1s4/L5ezyYd0ASnypa+DvJtV3RJ56n+YvxB1wRlVbJxPYJ
dy2jNA07JuJdAsvnzQH7wFQ0ONfTiubZU1bDxs87C1OPiftGjGr0iDMeoiAtlDWNMKchFm0la82r
XDm27Nh/DYBhABOKBsBACZJe1a/yZqg9XymdPAig/t/49Kg1Qj5Dx66dltnXYdM8XhPma3PfM1c9
TBDWP3AbINgpO+sQIPkgAaUnraIobMxCDnNV1fnToHpj/gVFRP9IzX9eOcnp2HpBMSbU8fwzBzCn
zFWV3izjZOI85GpNwOPXghCXmliZmJSf8PHnPzu14oz6s8I9ZzxIfH+j4XrH6BO5Q/bwXYUcsx/J
82tjnDQc7woZf+zdJDODmRPpRmaqmq/6idc+1lbiiuw+i9zlSJqTzRo1C+dbsTR+H1OHCXcpymva
aH1fzJ8fB/koHYrHXInLqPJdNYcivI9H6DzjBwwLpUCHUsaeddJ/GwV/70IjDa8l6jhKqWKO5f+V
5zS48NQvvI+tVQRURjVvhGkQrYD1tEHJFTedojRJHQ3aPrLwERR8j14c93S5x+X24zFxocQ/dji+
rgr1cm0h2ucq6aoDOiHjP5EeYfsSbGpUfmwzNDkSvcZL2GYk8RVsLQE0JmeTdIQhgMJkG2pl3kPi
uqvHiXsop1/4srsKSfNw3KKrs//C70OUq8CGl/pbiEY6n4n7NelAN1Uz6dMPzYhOvcfCxWYzswUy
e2lwBBrgMeO0BcMSxsrFFQVVY0KNYnKW1v2Px9Imv6VNRcNcMo7acxchEe+N4eFgA8rN3BsJHAJJ
GYaPz1PgnML9Z4qcNMQqFmAPT1zoKp1ZSlsFJWGrUhQhVKS3Yb8qbk7GVbZiYbzF8ZBZB74+s/3E
fc3EhTbgMs8C3wnNZOmDh3LqKDkuA+nzEp+alc6RZvNjZkdFaM3v+c2F8gSI3eNPLHFsDjJC9gb5
NxOH+dEgb1KBJQr0D5o9ZvqePch0lqMT0OUz1tbI/M+3cBKUD0OX7AE8Lg9lOk8WV36uaGbPUX3K
BvvMU+yX1ROF5OmSSD+RE/Y1Wwh/rjoBqbdnBBJ2pbm9jHc20oyeMAHnA1RkeWlXgBO9/bZq2qg+
adUdDrqiCgz4HWTAZb0flCf4SgN2cqydMbkonktSTQWq2XIzIBMeVPn0gfh826T4mPhmmAY0WnE5
ZqnlsN8+q2vvAtoWJAWzXA6sJgn7kAOy1K4A5VInMDtSYnPS75Dx24bXrc0MbAXBLEeJgfzJ5QN+
nl54h8e7qOdCqFkQYJXHxl2XrIiDyRUZAY6/xxK7isno9zIll3ug7h11EVBQzT2dfFv237pX+iFC
kD0zPah56wdDN7KBJNgKo982NP+dF1cEoc5FhbbGFSbLvZZMRYjLtHfug7QujnGGo+QFOj0mDPAt
yoHvzKTKqw9VvWfdA3SkU57bf1mlhShzjO+B/wQab0E8J9hKV/Aaun0EwhTMd6/itkb9CCDdVw1E
YPXpDwwM4Gte44XP6KbAt14iWKgvSIMcLwHQtCMkq5OJaW7vkSly5RgHkb1upaErWmsHYhXjxV97
PY0keEMaJ95B8QJgjj0RxjKFsLJaoCyj0Xjq7NyH+cDUX7zWHQt0y3cBISWEzyzUElasu/Zjgngt
h9KxcpdbAlXTi0n4QyJlQLGMfrC/6A1nj5hCYi5uVKbTLPptvEIO2EVURlji4jaH2OF3+S8Jbp5l
fvnePJFFOcbITQ3P17UA9Rv/h7dtP+XFFRHlN0ptrruNPaJlb1rMz50h9f6+MY2qWNpDGjE5QuAF
SgpULdEUWQ5gfhdSQ8+PwN6DKjso7jQMvU64xtXPs7rxnrQI/8I+p9ORyUnizzcKsEMdHooClmP4
hsb9UFd45qaG/knD3ZpM9PQPB8fODjTCS8PEoXcAUApMcENTZXIchlkOmqaMGEAMbP7VsZslxoI1
pSBeOFzt1Hej7cDsxHDeQti9GtCjPCM/y5O7YlrYa5WC0R2M6AmBoodsWQfghJ0I+nRR5guVjcN9
6nSL6Gyl9AdI07SwMkiQ+hfPux10xtD64HoEOi3/pLv6QCI41bdadPuzmUdQgKo37u6/g5MlJhDe
ficKGyNXkgFNquppxMhrtd+Jud8DvtBO34sIFkSL+fQhUt78iWflplZtH8exl2ef9qJOHj9Z9CpI
iVHPq/mbDXkTtGmbXsUzPxOyV9Px6AzcOmF1vU8QqFaeBFfZr0CDX0e+EEh3/wQ//yHH7l85AdDH
9vly01jyLu/v9+d8C7CM6FfNwhQ+QFuxn0xraFQSZSN2bwkSliiOvHdQPGAEd9TmQ6KfMGDRdYO6
dpth6LDG902k2SGdbqKm6IX9XIGySVzQaJ2lYDu+z7/TOy/N/sxNIxSSFJ6PeeZUMDMT9TbDU76A
7XG2GiUM0UtvPCARZorl9XyAEf7EYleI24MwWQKbjv/AzCi8LS0RyUi3Fg4J0r6d7f56/RmuE5Jh
N2EhaIYxzwrg9+y2VmrJ69gagHfxqcarE4mim6hvk0tdchCB8+VaZn3trxycGfFM03JkPIf6TYuf
uQsfFWUrOr5867aD9BuyqylVK3dGJXDae366Dt5RlXC3Z31EUr/3FxhmUY4fyzD3mK9pYpBMsIe/
DFVeAXYVquZ3TfLdCmMEFhVczrJsSOEvQw5HFdOIZIF7AYQkOu3A7Ne3D3Mkysg5RmmM9rRkx5U6
TYhJ2R8L4TN61Ime7SX+jGSQWuIrzNS9AAUjnmcdBojMOr/83Bars9lZrzq24UVYm1SuScZTvGTd
Wvf6BtqnM0gnAQLP9N53ijTIu4KKp/rb874MoS7pLKftqf0Cdl/yjm1E/ts5gaR30V8w242fhanR
FrTjzMDr3rFQZfx0/nqon4wwzM92UregO3RU4cyh9Cw2r7PbK7HD5Vq/xZJqkVfELJJPIuAuLcBO
Y5LtWyJi8mA64f4rUw1OJv4iwVc0EUMHBP00rDmCY6+6yhVhwMRKnKKqRFA/OKN9xAzuPeRLoupe
3ur/vRwNr9wwPP20cqK9V91nCCIAwknoC7JJZEc5ZySkdxh5i6khbgMhdfb8bWeQAXzP5XfbTCuc
27xPx49aIXX3WsjqJGLYMCOUTuvW72MaEl/WBB6hgCh17Bug3wyX08otPGvLA9XRdOX79DDe+ZiW
rMqDcbH/O7BIo/WXq6iIOREbx7/isqsntaSZPwLe2t0YAXzlaelqs3zbPZ+rbwkwldJRBZiA5WUc
snmHNqjZve7WIFgieD4raAlxdPajFlsSjthc3F+ujpKVsdRrH+bAVgx/JhiB9CnPU8LN83iCSIOS
N73F+qsjO1GlO0wEPNS/osmBFFJd0pHvkFh5DKjm906rKJFg1JOnJm67qHsaZxJpesAZiYk8kf7N
iCjxgQmieDDp3lxMdiaSBT93DjZy+5MvjWgKiljZ1eAzZvMcBpmotCiuYLnf354LB7GL1p8g5Hxs
ovJPfqu18IA53O6cD8znm/kxmV0jrfBBJYpD+p4jqSDiVJCTZkWpwWeR+grWPgaEhCOdKrfPx55f
MOsL9qfjfNmULqsI7qmPb+NuOyzK8COyJxM/My5duyvVFRqETDcnU6+qO6Gb/pqwZ/D5pvzuRfMG
ygLAyMnrs0Dj5FaMhXgdezdN7Z0KlQXXqmL7REGPPmYSAoLpv3jUE3R35DVlj2W56PFX6LeV5gxW
NF8bDRIYPc8fXrp0PHwHoKvEKziBA+PS3+1HPzqBg9NhN6KTAJNuaSkbmsuPsthycsv/gXlYDYbx
MCcODiTQf7j8uTwrviA38X59WYDdIeheRw2KYBJKzLZiWJOEGOF/WL7Aouf4PcT/AId2vDFQQI0d
9+CoGwgbKlgFTTsesaAOSk4qq3HLZa0FNa5tE5FupTiOW6lgFfWWO0bazpXdj7TD38Ybu2IdOW54
SjDZzkTAnYQZEP21spmEK3C61UVPnNgvLnCS4AyZdJatUDnqn/QCxtBU3J1uV+3U5eU6kCHzYzjO
gRjZKAappF+6FdpsH/8OGmvXhaUUCFQN+41XMrjicPN8QKsnHuvl4BezxpDz/8BgJ01v9pmCv+VR
Q8nXFba3c/6ehS7VEFukaym4tZV6dAl4I7W57wNkzDE45N4LtOLTDQZiBBQ1QmnsWj67/xayCktZ
7mtBRkVBGM3OLe778WkBGLZeRcBXtfuglb34iFr+BYlcr72CLuSeqxhzzw+ZMLeOQmPEQGRDZfdC
PllaKf5lQ6YGFx6gSofcUI4nb+R4bbOaffwGSXOL5imczlSc39rz7vdclt/HW27UAWkzcXg92n9k
m/gBolCnOA4+4yCwvjPZKqAw8JNwByERjI0XPdIuGcd6IhEmFJ1SfYgd9RROLNIIMTH64pwtBRGr
6nnvlHTQfyaAIUeMWbOIloqwy8GTGxyxCqSlpGclpoDGvRoh8sndE/Py/B/rKV60DEx/8YVEte+y
ne6th4YqbRQz8YsWkWJYNg0XH69EkE0sFzRP+As745V7lgeuFhDDCH1aKYvHbEfCy3Y+WcWdsXx7
oX15DvcPhPwzl0mrDWZQYmJbuCZPMWcc9Wv8KfWG/oHyd1AX5FgxAGHOBtBCxIASCB5ZWZbRf0MQ
2U4zwYewRH7+098MtRjTzoVW+YXAFzHIZkmMCUePoscc+La0Xn2WZy2d/L1cSxB97ofM4pRZPbH1
xo+Vd6WKKDxCfq/9CyZS5tq4xiHOgCZ5Y6aCBo/bePquRhwLNAIdsH7nn01P1bqrOHozVy8cqfi0
0iGAZEVtX+xClUBf1O2ieTRImtVlJtV3A3z6wpIUaXMbIE5mHqUOOLkiXNlaJKS5D/bLmhYoPpsN
9TZl3u0RTh/gH9GRftdY0BpAyY4a7mg3xY8975VsYaY/2QycVcclQiQyPpav6y2bPtUKC9BwpZXV
4bJO3qXB48UdwXasmBBOslOO54HgwKtahC0UHuuj0u0Wrn+zD3Z9jNTsjwfmW2UAEqpjiHclNaUq
1xg5BDPoUvL0lwi1+Ud8Oj3xbc9BFAChD1C8ifkUjMwpo2njMct4wxUgvoLY5FbCG0AVsBy3YBew
z+q+0sM9yVjVOgnmJQX1RPNJR5kacxUQoi4fJYA/QJgbUF4n9j2qrvNyIJbvS+TJYt4tMnVObhe2
8fH4217dR9ye+30uSxOpCMmtQ2i5sg/QAzccEjYMn7qyRhgVg4v5iEOUQoUgWcmsw33Hs5/liuGm
818RCK+yo+a8+fO5CNxAzM0oQkDzbfLXcOS2b04WG1v231BKY3svY3zLCVFW27HvqmfBboTephhT
tfoKgEVEOz5XoC7rd36fKSJBPFJm58wCKG1SKYA/PbTuOgPD+0HjVZ6nn7n4fAbSru5rxW9fbU+9
t299ZJmgQ5XEyUrMQi2QQOJUuKroOufgPNyarhX24qCkkscCZCCZdJSci0JeDT//laFy1oYIyGKo
a3qBrRTZgGFp39RCg0LtMDHUD3FIZMrRpqVzgFtLg0hhX6bYuJ8KHf7yCU2LF4DwpIcKuwwj0cxX
5Zg2379p15r8ZACs968OxSf3mgRCd+7dKSp72ugADFtzAIaev8M/2WCFvn7oBYUeE5oLKtoUG9fY
gL9USucnANS8gpyBQAe55lAe2CFyt3bK/n8Rt1vQfA16fsPPbSShp0HOBigVdEQHCXn2RhT8BV9s
ii0yXlETfKGiTJbJbLbByuQne3xjUHME+yKNxQ22K30jVUeQ97uTQ/ihd9ynwywdtF9EZVRe5ICt
yptpJbR5azUOW+q7k25BOh1m2R0Fi2F19HxSz9Y236rv5el8saxSkmZvgmeUrazJTe1JZ6ltEUpy
RlGkYl9vpUdoseKKDJlkulEq2dQ1DoPyP0EqpuUF8wIALXL6whT3sdV7A7Wi+3cHC8p+Q2OE89aA
haPoeCQsbuDVuy5EinB0692qZR0jpgUXHmOj68S5DMHf/vxIYXZEq6csP5dBklnVAQ86Ob0Yg/Xg
dLdMOrR6Y4bu2NFdtzEiALagF7YZEM/N0x2UMcqZYl0LY4yiPhK2Xq9MkE/5Ct+clHT2d09sRDxo
DotxUcE0cnsgvK4+RbpWnu55lRKwlFoHV9xD62SwKfbiPam8t4mp0TUx17jJmornSwK+mm88gkck
acBe/n1ZJ7tnbNU4AsuvYe/LGgDBDilZCOBgvwPbGAl0VVYMFeiMZzihFGt3MDEFlViZmcQ+SFzU
IHiupOrog2+6NTxWwqa5fJdad+24X6qKPZN4/GCquHUJjgAiv8+grDl1KtUYNnphKv16oMSaAWmc
R7QwssfGZSJqsVEEvX3dqE6q6nmKX7tPo8fBZOs/vEgACmKkE95+KnLksqiCEtNRIX7exEP2YmR7
YrXMysiF85qA1HLXOojY9aNYXiO4yQFWG9nT+hReaG9mf4QY5trT0gMTVvBARtXosCCYlNg3hf8Y
PUmJaR7B17eGXJrN4bxTmptw9N2rC0QKzrka1G3vmo7Fk5f4pNA6LJZ8LZvilklY22sCTe1cm1SK
vTvkpjn4C9WSpjTtbYaNe9/gxb6r0O7gXqEodX9XgYleiVTwu6r+YdsvFo0ohAjBjmgtKqFafxsE
IXB4hdbSy3CdR8O5Kp5UWEVaVoiG4Z357oYUc80rr4+WFAGF9OyE1ts/r2LNz742s1hYq6VPQKSd
orA44ghKQTYd41IH9DN+fgEyqA7saIWuRtvP1ZHzUg1mmE9GsPkmdXx055wu8IFjQr3G1/O1MtQC
O9QXeXC7aH7vUNmEVOO5q4YoBDmyqYGIRZS87LBi7uVpg4xQIdFJhVrZCcLMS5UWmAgrh5TZvFng
inszyPG9rUaaRJJJIPDkkPygaWsijGQJyhV205QKuOKnhs/ieIo2pA6rRNKW0tRidP8mWAQnypCt
M18I2pC8GEVisfiEvUX6GqZ+LxqBKz+f1uvH056FdfnZ6XJltrnlrezthNcDz7uFgcR5NLl6pam2
1vCInuW4bONKEgXbmwIcVEEJAGVUGo44V0siYCwS9xWgoziBVd3OOFezYBZ9hChEJPnRNtNjWk4L
sMz61h4v1j7kUEKh2OwiwVLldReEasHhKU2/wr5JPEtcIj/rVXmH20CVBuW1vrW3e23F4m/p/uJg
0yucYyVQYF6k/JPMKfjwCx++970KAVHPHtikuWTK7YMf3xNV6WQWQkM4LdCcHkfvbiQjjnxZ2LIP
RAt/LxaByeEvnwZkd2G9iC/yNHgY1YdcT/eyR47PN1JLfMrkipynf1D7BfOnHMyo1PsG5R2Ggco5
7BMToLIJ4JTJ/PCkNtaJik4nrwMAKwK/sjjOjmCvxSKYo+4P6TfD9S4uEED9+SPstCGGytA8ZHJL
+PNVtm5QC43KpZ5RoTUp1Xjvy+eb24doMLmsSIZ0dqWwj7txuPmKFybzwA+2jbTMjwSWDqDu3qDW
kFTSYSlwNqzPNJZfYtTnutB7Vsz/Yx9uB5nDCoEc+kP1bn0PzJb8aYCKok+KlNuPCr9+mXogAvtC
t2bsKpTQAx4HNXTkIq+FE4gISQxKFSs67nvO+OKyXstYF4Tw4H2U/8r5e4ukN5N9buyXP2p1MLWK
Gs5ZVneIec1dt7E7DOGiHS8dclnYWknHZfBnm/8l4NaC6LPXfaujhe1Vk8Qi+qRGvL1RGamtthc9
2GMLfvdhhkd2U8EPMfm1uSsosQlaDKfd1tExj5n9/Bh3OG06j8XF+43TUVGQou1zX0jIQ1A/Mutk
Ew8Do104qaZ+gi+PiR44lf0gC/emsZfC0w9yX4lpIDsUV6Z3oYJvkenOFuFKGNqLsxhS8dpaOp/c
XEmdc1j3n3iNpV6XbkUBQj7JeKoaUUPDcwDZLj0+zZ6uyi5lsSCxdgzDBTq+OCq9iBpzc5+18DUl
qCu/rHq1I0+NQfF7eshzo/xMshqf6DPErFgqc9YUQ6q4yxmD6SYklQ4SWcn9Q9RJASUiSUnhWxTO
eNXRQ1KyNxiVQI5rh3zuJwLiO+4tMq3slVS/UuvKxd7j1/OjT/HRkZToMmm4UwX3DfRvIwYnKWcc
Mg8mQA9wArufgvKVqDsOR+OW2QxWUXMeAwpV7AYUB97ojk+r6RhvwSNEbe3XzuCf7j7mnAae67Ep
3/rsE9+gBNLp4/l42JN1r8yInyGVlCyreoOKViHF58VRTfG+H7XUUpknohe9Vy9KuSaIRYIs9Gwu
beqmJXyv/yDe/EU+NoAv7qVGLI5QCHAXiw4THu6ZqR/jEQn3od/5lBm53NNS9bc01ZbeyfGJq22Y
hVlw/OKaV2/PT4u1B7HmnbgwkP2CUvpi0Rnm+Ht9cWZhz07wjrMGPViu6zYS9P+eftTjyjMPS6+6
JfIpd0EINnhV+BSF2BtYxM5kgEfUEd1r3UurIu8OKe9dqZxoB6yJT9lDTC4i/jdOj9Qm4o+BVORc
EWOIiu9eIkoWtRydEqZ3TAUQaqTE1E7QB+J+7SXXmqkizSAoqkS6EjcWjYEP8fLhKBQybdZ9V74I
skhkeuzOZes1gLI6/ez6V4dhgzVI7Rc+x3F4H7W8AaWN5uhY8AniRFE1SqdT8YlaegNh+FXqL6nk
Tg5AsBvnV29lD+L7KtSempHzRQdEfFZPG3x1riVo0V5YmJb0b/Y/hTzGr0UzUH807G8quhsRD2Va
Ho5zKTNN6KHqthOTgOQGPM0N4oAq2VbdrXMV6SUUjJ3K5CbG8rmyaJxBgzRqfGj+i96wBeTa/wG0
8EUbhvhBQQSTcBGkuIF/+GBAMzkwV/NOIkzT1KtU29NonEVsnWiRUwtLVW9uRRXlNUQ5aRJKw6qD
/wg3RRI//3s4gwZehYD0WLY6EEF5HKzyUIIvGGZc1XDZnMyw6p46IjpRgUJD1gGwJyVmwfyHO3Ul
ShTriOkpQc80GAIRGC/1Z8il7JkJ80cSsFxUVxsxDJu56hI9J1mlvsZqwvTk5z3SlzzJeL2+y7In
a9wE95vHNsRuWsufMSvAXbEebSimUncc35mKTkxMozFOXBPnyZ6HB2DeFVda6SaOaI+BQLtuFU2I
a+HBCbR91v4Gu3KGUthYDfWn/0lEOQWeArhQ+PBPbO+8KtDowt9lCKF7Ud01VHPCoVG0wu92eBrG
ryzVVep+N3EWIOj6DBioyuieT0xmInHKa7jxjI4Eib3kbemdKMakDyzeXh5xET65RyZcOtuAJcRg
lflTtfJPF8wkol4LbwgwloD6zvqZrfofZGQVXs6WeTZ8vCmZhuxjEVteadNE8Dx7CFvmQuR0ohIn
3pds5YRPTPQGzqOIvJ7CgSE6iGcxYcI1KVikSnr3z2t9PY9WDjxcR6/vbiwanFk+9eKHLWZqvhJx
jH0LKjw3wKa95a11jo8b9iRSOmy4Dmz9xcosM/hIZ1q4URj42DxuCVruxXMTV/D1QkAPnePSb5tK
Jrc34Ey87Sl/AMTcXe8JZOFHL8pSzrYFYWNxVn5UMEGLf4j8P2lSZ7cDsiJzW/XTZvYqVVKNlBQf
PMloF5Hd+UAq6u/y4RjgKK8S+Ua5Ol7Z9t+3Oq4JODLgeRwEhbTlGBc9EpoEEg9AxtTBzJsl7VpI
lUgoTmzTRC5oMrt/6O1VFWUQQbcbemV0xqhb6VY6+NSgSlNV1xtHg0DvQt29946w//myQxrMtiFO
KTJUKvOYC0b2AR08Qal6sdKeXBW8K+By7XIR1vYstwS8AwvcjPqhnLBlVh6yTD6FI2Riyj8kg1Bh
xkJgSUXaexEvx74Z5cKqxhK9uMiVIIv3cP6aQSXzGm2F/BliuZ7rnMy3+YARpwk6HxJoQNiofUDg
RBvx3GUS2Dza8RDOyt6zFoyUEb6q6P2d1+a2pvbSdp9scG1OE9120OtlfAgN9k2eiTBPGk+gtvL3
bvbYI7w/hr/J6JdtsFBpSrc6tdykU/qmIf15Ra5x17rKbbz8Qpr7uKxDW25N0jtNe8h+bpFU5TU/
Ogq7JrLn7IXy1hSlnqLDebewu8FBsHZ7JM+E9meTPDxpQVW7yZjTK0x4IpBRNEUrtb7LRkEYLjSr
LLPmvQwycZN6djDuWsrlb0N6QgjUJMNSpexUuex3xHsOuYNtbvmKG2XP0n49E/9EXnKucvUlx2le
0ONVdCOR+LjEnbc3Sl4i/Xw0b99E47OvjHRfmE/h76NGcM9v2bs/4rR2VXq4rFlSTvfvZZYM7Vbt
gagONKMUcCc1MHB0yBSX36pVhQXILzKRSf7LJcNeQHnofs9fdh+YXO0Y3lnRx1Isqv7Qv3prtWfu
ZgV2PRyOJC/rO64IAylZFZfwdF7sAisTU9r2hQvvzgwMjAPTK/mZRxkw7peDuCYFgphzlmkpysmj
ukXYwdtRGrFZHA37N0NASC6bnle6cHhMC/aq7ERNVoKQwEmRcz55Kp9kvCO+uCi+6evIoe5+PnJd
z1+LdH6Wzi6DkifIU896iZj1SSCAjy3UCNQBLeghBDLpJ3Zk7WejElIkQZ0h3rOiqnCIVEIgo0CG
MxhVcWJmKHjpcUFmeTsHau+V2InLzTJ+vayWvEF5Yv5FfLVZofxwWhDyB8ByicB2o32J+WrYbjqg
7w2lqoVPdGAD5Xy1B5l3M1kRTP6hIAdamPTPePNMtvrz2L1k+MdAlHKcFgwPwGC6+tCkrMJYS4EM
1L4SRisetxCHywY9vgit+hC6QyUjyOFOtE0/fy/u+ELqbzwt2g7N0pNjFSgd3A9A1e6GwEB/OpgM
in9DYs9KiE9Issw5Die5rhm1u2kvIOf2eHihj9+aKN53Rl+741r9VmxgYB87EjA0QuIselxq7TO+
cPj7Tl4H0VPsjD+jFv87G1yJvM3a/fRnWNG0K0cdPGIO5xM0ROgN1Na2YeoRvfaBjAIHb0XnqtVE
gFyKkQYPj7pqP6NNjtcKjX2AK1pD4E1CjvMD1tBeTgTLrAAldEy+VewMP1xrXrRo3Uj+ecSWp47h
VJhiqK0q+6lG9q8M/HeYbVgcyZOoDTmlTfF/JPnTbFtp/q3o8aYeGMGB7kfqKsv1snwl7bhb7l9D
b4KxXRROSfrdfu/qrb3FeiMmXwAeGx1Q4pRzNCKijdHmFRWoalVx+ALFFurbdwbciE2HTAYzhogO
kTg8dhaTl5OsMlO7zY9N1jpuOZcO5UY4Wibd3eMOBMMyqYgxZDtdW0U/p4o3X0ZLh6/okXuOvTrz
DXtcHs6+90wL/Kve1KI3iupd6SSRgxavm8LbSQPwHDhcS8TEChyQVvd3Qkhu5NnhMB7rDTK8749Y
xxXnMQt+wujAVqaLk4SjOvUIPWlM4O6CX+nCTmOtlZnnrHmpC3jPqeIuYPxKN5ebWoB1oGvX7My0
yNoqfSlfUcDxKOe/H8tl+3b9L1hAjqekCDYKIeh3b/oYiJetNCRe0K7xidmFgThn/OTAf+8GU5hC
2vQm2Bhx1r+jy8GbCDpd7A8ZKWcV6CWsAHfsyGWpUTBoQM7ZQIEKQqzeMUtLnKK8K488dNCuxWqF
ULUqfph9tDdNUDoj+q1/VFwq5HE4jm5m/HxInDgRny7ByElT6gopt0nVHchLFe09R1Xxq+Dsw7B7
JNOgAqy7v6FCwVSnR6GBEqotihazinQ1zQRsGd0oqyQMnW4X9YcFGCpn0dmMby2+JhPGMIJFQ04o
RLCDZrsU4JpyK2YeqpWdZnFOT6KYoA4RIvrJ7OKsPFZVj0a/ChV2uLBhJ0hCIAf2ag1CtSd7Yhs7
S/MkQLFM0TezZHNGd5/POpK5/JAZogtNlD33v3jdWr8rx4sPCq7/z8+9HNv/ovuyqYLlC/b3ctUq
+DYNgBTG0xJZPfGUtA0e/iQpEyB0MZINcVFU2aSEiG5GLGkEtvLaBtISmR4Lpfh+nwAh/Q+BHXB6
4Vspi5fyLunzjsJil+6QG8kkZBCo67hwEKYtoAff4Oyvd3lIcEJ9l8tjdaBBZDJL5DYl5AXAo9fy
8hG/OOWc26Rev7Wj26GtcgT8oecdWhU9U7iXtmWliCyrT42V9V0wGZpTsYVSlMkjTuwpzR1e9Va4
iBs2+iQlJCJnouW3eLzAgec5AbbQwFq1zTH81f4fza5D3Gn36WZPd0ke7PIZoOWmEm2U8iW2GbSG
7URi0Hy9klhV20+JuM2tnHNsEhM999ZlTOiyNGZ+nw/I8YzbTbx0aXufobGSFR8xaAIChOi5fy16
Ql4yQpQDqeUACT1ITGYgSusZF/vH/MM88iSBm8Lc7hS4nf9afuWlndtB4chMwqyBYDY7M8Ss1bHN
+DcC5j7qFNRhtbR6KIAxYYLLUFkRX91lhIG5nDdDGskfELXxLzP9jmWD3TauqW+7/2seC6lZrQlt
ZrCSKHvfNqkuj6qUcnxyPTsjhd66ZteJa65BwY/g1iulZE1ZrKc6lcIdgFh4bytZSLdfyaFexPj8
iMQc4SsfS9N5OfF7tR+Bc59RaY2oU8UtCWYWnGYyhlGV9Z7fxg32bqxDGCqZSLJR3+yboSTWNGH0
gxwLls+jNPdnrsTSSgxOkAySd2/twa/EKwDqYYWu+Vagmb9zjhYN89vKUOyknxLei3Cksacq0kpB
OQJmM2t5SZuY+9Rd00JQOfFfKOGH9FmuT4RoXqYw8knwGr/XeF/j92to6lRFemFHlhe7tu/aQ7yg
ONkvq7mZvOqXbaGT3+Urp4gtm56Mua/lwXVoEDeNT4TV2fH0rmP7nIxZ60qWwtTUila9UxvzD1rS
8rMgTCyaPEZr6to73xy5ni2vPM2XGl+UkUB9D6bSsKJX6E/pkqaiwPmnPsNbc+QAQjFzIUO+5BMH
L/3IfW7v8FZTUNcbemy0sPVu4AIkpQYA9wob/mDx8q/W0XrFb2jjfCRTPy1lyiccjKSf9lkt9BBl
RvuKfR0wOz+HMdo6oIAfoqZB92AOzAj/ncXFTmO3rjv+iCDZc3d1cb2dDmdKVGlPr5U0Z6JxBj6e
BOMhocB+lpMHqdt1y7mb/OUj1xBqBbYc9Bw8ECIvO6p3UeIr4bwDl2D2jeQ9UQksi0fnQXF8yZ91
8rpQCZ1zBhA8JrUnbzKEkwk1CXCRpqcuLUJksVMRo0UnXVcbLM6WIeiIis0dHciqeoAK5x8uPU6v
Kb/fAHbGOH2jig1tU8UDmTLSk3RwBjFX68Hress1FhcDkruW9pUhqrHK5DFyfw9+711PXioHcHPp
BzpR1NQdG0e2NBloYEPnUecVgKotQUZP+aA8syESZ8C5BPQeWmenoKPpX+9pvhp9aFgCZPq6T6OB
XCT7WcMj7ZKXDHveDhjXRGL8pPmwqG9CYydkH+DrN+EcTrz6oaQJNT5mUnlMqdMVnVxraccu+l6o
UUrkWbxwBWAiQfjNs83gW2hjqp7SKc2w0PT0hef89B5S2dmJMhbqoln+1bHSTqwIaBun3Nf2w1Jf
ozwplGtHUKW6XF60A64OCey+QxVCVYbWPNVsWN4BcYosGm75Y48/n+jmeSJDUezooCUVtznASjc4
YG9nxPGxJs827pxMMmBiRskB/XiQHOB2PtymIPAG6BExjPd4b/TtCqmKn18Ghl6gqY7+Yy5l3LXt
KzwjS62AgLizK/dE+xKYm9jVva32nG2MznjVARpM9ATyp/16fm304jSZMkITx9BNuxhnv/tvTvOo
eDssf4t48fq/kaZYRvDi8u8MGkkgDPOdiXYmIntifiloYMV333egAf7JS4twg6QEjOBrLXfXdPum
2kg0Zm1fK7TZ4KkrAho+rGMuQjuLVN7oQQcMX1QJr09jchIXYEzRFiERhV1Ih8ZHmo64bK5YGv77
9OjU7pHpg2jQgRMPejWNGeETanMIZPv3ddqoTi31SHL7e4F9Z9KzOuPFe93aHhLTAHhXeSyXgSjn
krpseeceb0XcN+bLRvVm9ebJkrrobWYIuvPXx6cGvVevTHk7G/3SKWekK5TlGX4xBGG8suIWBFUZ
S65dlDILDssN2h9PF6X3QdKEiYpKWZFVsTo6kbiMJbIG8eQIawTE/RUhhHHgcirqBqfNtPCofRaJ
RQSCPeCq5H9P3A79NzZPpmJZLMVHYPn69Uw+lZs07vbVv0rbFUTwjijMSCF+z4xjzGRB3XJ11Kq+
wP1EkxMTs8X1qOX1ScG0DbWoSL7rlk8B0tuI2gLv8M9q0gK4gMwE5P69/8Nm4x5OeCmOpEC8x8XU
/681JDWoZuxKppeCnkXtTgqmkJdpF2oyqX3mevoxAis0bxcn6JdxOK0BZuTmEelci586TrOgGd1W
T77gTNrgSF3RrFzRbWYqIUnuY681MYP/C2SrkWbSpzAKGPqz6/jpoWNpbzqGtfNRr5vaQ07BPc3R
03Q0lG5zTKEQHSiboz7BgndevnNKcvah/OOFHsazTfMvaxssJi44KoVnRX6dRaz55uV9YViQd+ao
ngESWTe2h9UQYID54iHK0NyOoD4blipmVG9eIeq7zoFBsrfwl5iCoNxpcHzDzLHn9GpZNe29rylq
hYAejzsZ4T6Aa83yXCGn97ycYN3m3OKnzgBOBMvrugRD2ecCM4vaCwG9oMqT3PisWUT/RPKkB06x
f1SKLy7KRX4KReTfvJDvg2e2pkS5lyukIk9135l4IVeYGXqgN2h40uCkl6ozYmPE905XVJPFbx83
9Oyyo6dnMNZYt/3vtkE1xrzYiLz/hGlK5zmg08RxajFltWSVpLtoGClqFDOVrjqewwmvUx/Q+GMv
712qDsOOpykio3wQXPmnkRfyuKVdPObt09s6lC0+VTvsIC+5B7wfD0Hq/SPcopu687WBVff5dBzc
dJeuSaIeeZgV3FN3d6kKuPvJkWXch/k7PjSw/SXS5Gq41krrTDjr33KhVWTsfpYi3KJlEa9RQmi6
bZACrDwZjBB29HMahNm7Dok59FcZX9QXL+kcIzr7zOKIzUXBzlEjWJAdDfDac+j1qANk1KM1whjy
xbmaDN+oyl1SL1jtPQG/3iP0Nl8O9xMudbf1iZ9jUt7oj7kXbjxX2VajrQpWUDncJ2dpT0pxjrcH
wuA3VYSgOJtmqTgTfuJuV0C0VVeIH9+4WSUIqEvQ9BK/diWFkamSjW4/92Bn9Lgf6kMxP9+nktH3
YbUbsHyStn4DPFdqFQBRhdOkc5OC/b/H0iSvK99zwlJe8nA2KDn6q+Qy6sU7jPU8siiCQ6ed1oRW
ElA3wk7wIcRz10hm465pIFhjX71N6y/huYe6VPNtXP5y2xrm25wJrPorBFhy83jP4j2GqZ6EZ1l9
sao1GGngeJaWU+S2w7ZhV6wC6wGzIwGkf1gRHcFtyIuf6b8nHm3997xCJT/kGp9iLtXUS+XI2LLm
N255gRszkpbbhccUclpXuMauefzeyM0YkxVRpXHtP9BabPaX8wtBzoS/geZUR1fpXc4/ltqmsttY
hpllgeJsA2ih5eBKV9iNJKUPkenCNnzU7KIZ9pS5txbReLEqeVnxQilnSnwt81Srk3ZKD9suLCSW
ivPr+1yRycY9w68WmLMHwvyKUh73hFLUX4q38StJWGX4HwgQks52F/9FbajMawEf5woRLUMYepMQ
VvlvDFt6yocL6OtUoDGpP5NOjIHTP5hjflJlR3b+7wtw5xbCe/mOZBqlCH5ch04kOqaMO0Z/4lbq
EzLQmUnTMuim4Nmk3PfMiilTgdB02Ow50hpEkWbtDaEF64HfUfoDu822ioAuaKb0bLGLgzpjCoIH
uGVeVFuZJ7tltFC9g5NSaCj+Wck+wD4OjsWwzXvre1XF12NiQ1r+ybzc1uMOeJeOXOWxLoznU/k6
t/YYYUt2lEn9CXzxqxCiFnSQ13fevbtVeOoA/tLZg2yIauexG75wW169FNhClxMklh1w5RZq2cnC
VImUQGa57Ih/UpELoGTfV9kodgp30MMHHU+bK9a8O4yXjuEKz3KgeLJY/BI8b3vFa0OCMpRNnwhU
PPqerj8T7X6p1roQRJYij2W79ZiT5PM0JTd66gsVkaKpqSvaneAT19a+Ta15jLB3EyEgIaQCq0ne
GmCr80kc8Fj3zfr45aR449YT2JCzuabsbJODVCP78qaFWdJaNi7caf/CUBnk0kC33uyPCPXKtuJz
OzqOiHE/IPyMBntGynNwd0jEBBcwS9XlXsIUG0x35329wZ7P93J4dg9poHVSednnKUPO67q5aJ2g
wIrgJCILfqpnskw/J4irJ02iA+BQ28+KJuKPcYLRLlIAfe3J2wWFJFg6QlyqtaA1dRN0wCxtcZnI
djZqryP6QCKtC2iXOX+RL3+wxjkkRg3lrckqY27vjdO83vhbxj/ldpc2HtNzuAPOB2cgpVnkofMz
v4lt2xaAvmX9JAgeGO5KoDrPIBGOdGOKDLejEugTdNNStZLZ0359rr7dyPZ5sTO10FG9FWOeiC9y
ROc9LwrTxKbofFyyWfQJX/EDRY+xrnKhLCvr5lTN6f+gGRdg/2n4Qvdeze5LEjhh5jz4buFntJTx
CJn7E/Nrk7/zB/oi38P3PHkGSTonIGgc93cMN8q3QVdtd2eGg3qejZqboxKuWCkHm0Vx4kAmOLmS
dwkReLIFaVn9K324clLj9R2pIBFTc3o4ODknm7un8algl1NVSdobCTjU4M7OxlLscFSzNtsYWnt8
KDCVT4k71QXnesABizTSwpr6PmXKndjl1Zeb9Y2AaAbquPuBf8ggFrSdNpBz9FHtlV7Ksh+6418U
UzJeJxytNZ5pxJoUCs2Wer5rIsk77sudhLD9KCivR1f8q2PdGuvLlb/3LWqdNb+vSrMiIAPxFOVI
Tmkk1V4QhOmgtSf2wmCl8yuoZzyHjF/B6BMk4fNVCmv85Lb7lDSKQjR1E7TMhopdONhLjTC6drWX
AHsu5X/vedblrKUG9x79eRe7xOIA5aqY2gu0elH2LskGK4jxcbB5ZMEnzq7+xuKwHE846ZW6hBIb
0NEoW31FKFjhziTW6jefrH388XEnkZzCHZnHNphQMecSSN9lOIWwT5qgHbLJ712uNiGFA708IRo8
MktjaCeE2f2alOQdHkETFTNVo4B6NT6ZLKfVJiil9xqNO82y+nNKYKcJXCQjtqFen29fEbkqAmyI
iq0vC8temlk7hg/QjmfUFL0C9IJMT+/TsKujndu9PIn/JsHhdAs5a5r53AlTGTCIE5KkFYKt7kzg
Kx+8ngRYtioAZbdZdDc7qu6jtKVHuOLZDzKp1R21cjV5pz/WIlTRW/wm1NqsWncI4zCLOfGEh+5v
TO0EBxsP7rgLvDvKBG79/QbkQ0asyVmXNd+MkceAevlyJO05uqMwwAaUr4mJJ9PEUU/fNeoPv7SA
OcnUFYdENwWWdTA5rwZyeG5G6Uew6JClFP+aj+/wpTSyaIS4b2l7Wl8zzMHJcUpsOtSNS0gLUwgj
IkyeZbU7PBxhFXvpjkpDeUf5Ncz/L6qP21H0bj6ZkIFIku1sTl6Q7Bmn3S05GJBaBHKp0+8QT4lr
EC4QbbMkqYT4p4AhT1NH4jnMn+4wS5/EgLxjlTgs22UyVSSLCh8L3ne4oM1VUfvKrXn8ToZJMgIg
GzybL274I643jSmN5Va965IEQ+iGpQzvOFcDEXBecZm5IZ6MdpY9Ya4ZYiv2l/e8z8owTJiunh3I
L9ZhqnMpUZ+mAAyL9VstXetFrqMqkyq2wIX4Zu5JmzkJlnjINMh2WmHwTdTAGn9cf1aLz/muOIp8
0nnppEtJDJG37HwPK1tLSF1So/KABKt9++bvsn3hlW6UgyQCHB1nNqd+7smyDFG6UAybj5oCVlDc
UGJYTR+D5PvWkfZx9IZ2BfWG9054DNrm0yfn3VxDKjYcXPlEIVNr0Sc643wOMyUBPymWr5ZIh93e
WODFwPb3azMf855hVWL1pd5Jw3/Qof3p6/F8F59v85wAKVikcjmF3G8UNpbQ6MYrxm8gWcK8kXWC
s5nKhpGj3EJSUeuGqfJEVQEJLZxAbkJZMQHX52Ggy9u5JBNAraZvTHIX8GIJGuDIU4F/+hojL/zk
L3+aQC1iDilImaPOPHWoRT/7EGVohllttfrEEOx3P+y1SOSvDx+5D7fe02WNIcDplGAhZzHq0GD/
MHk5XNBFgBOfCknbyKj9u5HgWqIbme43o0VL6+xO+6bscAWFyUAmTgHGwm9Tm+ClMh4Njk+NFt6V
ff+bn92ZqW+cs53zujHhbwkIXMqPXlcBXHDqlxnpMihNcpZiIeItOiQ4Gzfv3p0vUqDXR2wqKrRQ
VSZRtUzhqokMeFUEXWrYNdcP0kDnbLVDQdtcZu2rzWWPbazGjghZ3zUBAZENclKvpGB4u0GS5JJb
X1TiPDRyK9q3gKVLDcVy2VOTNKY58SYK7562Gb80qCWbJ3eFYY9iR1xkhaZoGlo4+jZQliXMh7RO
qnCl4bn++kn4S2qXKUPGWzOKptYiqDft0/IdJwQj55JVAWoK54fMGpC2THnhX+5CzIBJ0lJiOaJz
ZHMgYGl1YE7f5eQvfF+L7AxluOi4dBTQt7SO6BgycRpwK9adOpNLFxebRSWkZ9WyGLinnZh0AtOp
CMgPvOFobLVYzXGNCrKjY4/kb+Z+TGI+ku2hxKa2JW3XOoOD9RPElNYebDeobMVeS74P2fh0h0gA
KU76mVOIk2Wd46y7c8nsRXAZ4CvQnezNTAHX7tXpOtGdkTt6q5knAp+lPovK+emgwQ0v15lJvhiv
uvGzRlMPc7igCXiGSa8yn7Moy1oU9AFRjnv8/NqO5yuK+xvCSmREYE4WfRiPqS0TzV4+SHQyfelE
iey7FzyXWasdFHqpeOyAD0BVHspzeDkjLrpeYLYmhl+onL0zH/cqKkq1oAfO7tLOG76bK4JyH0Yv
8HSxnZCSc9AsXGljGIsQcdJZWS/WjmFIqBWbpohgqsoPF6ev8XysEFfxKS6irEvJ5mgV76vblPa/
SusqotUwegB7DXIeXkq2lUT0PLMpN/vR54KDxGGIVrb8FqEnCjL/RptYhmvG5EkgEibg4XipIobd
Di7PQimEvnxs1MUgLm0aU+wc0liJFWh+aWh7coyJbAdaRLZbOOPeZ0Y7TgmD2ocxqaYpeZjb+pPn
JgRdvovfym9ltCKdMzZ2jzEb2LWSDOPi6xVX7ZGb5Oyc99fwUnggrtFDW+KV5+tN/wJq0k+7qdNk
2IWrrCUqqisAXkw07vA/IvtWV3QPi6mPGbg4aFw/yEIYVgNbQrcqB99EVXAwD8VNsaSYk2VJSMSy
KFDQ+Ug29TJwEyXGUgDTaLdNfNsaW/0dIMJJ1zBM/s9DuBKs1V1VQhH4mp1f1jbDYKVolbDuFSgr
BCarKf2YqE+P479jQPBMmRCCMNn7QlXFZ/CFPZ7oar1hc3ioD+IvohoTJMibFskusnZYUdyun1GH
JJhlkJ6R1keraHkkq7QWhgYwEkjfNk74B9D6eUvh8zydr5l0evEbY8kxYPgYXaLkNyrfquz8aCE1
cuDcwlJbyWHnuoTscCOmcHyHfiJ/zfsD/VAq7vf0zFsr/0ANI6Jo54Pbaurc2IgIpq0+0x6xGGci
xT1AKAhtlVY1K6vNXOsMRHh20ZepJJu35UuA1lRE8sLHqJBYa6l8d8MjY6N26Pd5MxZpOapYmT4H
sz0eN5iTHJSqgF4ALFSaTJQXP+9EEAcECFIIDtAgXtK1iurYLRUi6BEnmOtCok1jnhj1del3VgWZ
xllrJ5jvT0XWcZXrxDDHsPKS4A712d17F5ZOtkLggEFkjR7mdguUozqc1PG3YvUdfmdkLAgGFUe0
jgdJDMFH26PUAc+jJ5eF+uyojWVb0flRV3Pe3/PyGMFZ4MJV4jVHOyq1tl8WRXc5pgFa2HtLoFJx
9+xwJ7VXC38bUJ7NAgaNcj258rfJOtVnpblz2HdwKkh6GQ0tgb+S8LiUzYgN4VWb3xV34SBcNZBq
UxN7ZaPRICZVDgDjF2OnKpl9+schbiWrjlKA+Gq8ZPpAwtPtI9V+dwGunc4GM9lQ5AwhAygUYtnF
nPRMw6a67wQOCscFe1Vtm3ywm60IpUqbD9yzitWC2TOWy+QKDIR9/H8w46ZNLsvuT6bIY9q6H4uo
zxRdXrZgsl9d4zJYNyvnGq9pgmYes2Oq9d6HDtrYww+elr15xg+8xfaQtbKjE82Lzmntb7/URwxd
VKbBU/s8nHkeamGMhkRoTrJoKqgenkjiVDbobO9qCQs61ykVxiusJ8TTTybCOm4Ow+wZb1dsdSL5
Hg4zI/cY5KC38gX0r1MXL6nm8v01YLcL5zH6fvUERFVi7xB20jH5MnxN/k2fr8T/8yDQNa4EPd3F
GtO3BplqRmu5jsqfX7k1BbeCswnwia0uFKXenQAabzs/uFFlG3uDE0Lvt3ytFj/7oqlkrtKTw/UU
oEcDNE1t8C/pPB2mI0NnyKPyx8lr/8KzvVFrP2NGA1KdMZt5480wlwLFcEZlKJ59Y6j5TSMqibp5
DjB6GGMOb4BPg0EeDuBT0lF1dfz0KueR2L/DWyVe9mzzgTSVH3UnGQYZnyvIsfEcwkjxqP79RTlN
V7+Hh/BulKuoNEXXfUcOU99pCzgObNPvLJOByH4DsK6xnJyQuDuOggCvFdf6ltKvUvZHIH/t5xsQ
fLvSuxx72XOB4+zYgtXxdvTcGmLdHpnmeJXJIPrdHUsyC+s/x0YZymCT0X8ncwRb7czjU8KzftSk
gWoHz8L0gjDYaQwRQKkJ8ly7i6/xIyVNla8NzYslq1E4fw2sA5Ig4RyCmUxJbqLHviU60roCgTpo
fPnOMGrnrqaKHEdef/BD6CfCCvHTvsV1SZj3AOhxqmDoPJmqRiCBjRH/E8e5I0V4+qjhifJk29bj
cDcV9wZ+QvY8cLTM2SBw5gQ6eLsQhb1nPgmC7kDjIpDNuqMu3HMOiBYkqFEebMSebTupgTDXK3VI
seuJAgSsHQkPh8b1LLSPgluOTXKTwMgrJMxG+RXOXYkztoD+n1uJfZQQcj6qiIYNmgohdkYlzcii
upcUuZ58rN53Jlrptox2GWuOJc58u8CHCJnmZp33dV4/4wJ3DDYeMIzxljwl27wVRkhTYjO6buBW
DIMpurqy2obOKkNJzoJL3E14c9gkrJAVQSWpWwt1tvvgfKR2n335aZYuYwvr6Y/DwQ/llTL1SPID
fpU6gwSyvRkBmn0VV4nzzlHhK1Ugm3oiHxv8jcPnhX9rk33xI4WxzuNfVdcDhPXLcqnVJsSfxkYb
/OrghIpupuOmg6iKIHrv+v8qsNIQnT/LWrBjxv+jLGdTZFu+i9vD6NQ1oOwXq6EoDL21oM+MMsB8
VseR1RGSP4nKcy2wq+nLJsdrXORjivr63DcC9qzdeawULlIYUrrhhED23REpBgX5J5O4gE+3ZJnB
irkbqIn8it5GboFnNruUPDZbDLvpymVRiQyF6RtN1BgTLmP01hx79X/n2gx4KJS/7EuYKmdOYNpZ
7R29+OJ9uLHX8mzDeLNvEm3lgrHgN/accEdO6ZW/7fPh6TUcVG9ac8rPZnPVLofDp5laVoGX82Os
KhlUW0n2Ams2FIdk5olKqIjcF6shgRytvXx+D0VzylGPmpYriv8YeDzwBpQfc2s22mRal8t4vJ/H
nZYHI5Uv0N2Y82IiuYaoAkLu81ewQUsQ7Hv7i3V6dmAj7YdJcScv7lWgJME1Iix+TMh8BmGjylBQ
8a/JNcdgVL4zgXIPB4DL7F8DRd1KWW6DAmBt/V7WXbzBG91IqF75iGSphqHBJnbcSJ1kB18w5BTj
GrsWJ2xNsXXZaGuFIZNBLQ7R8ntckpxOgqJWdjcg8fX1FRiw5fv52yAN3MbFH6+VX+5ffOKoiC1w
Nd9iC+FdUOULcdg0ijERPDNBS1e+Q1CLGt3zZMwk5Qv0kBTAeKQrAyYJdKPpQFDd/aHrRJ88kMWz
RaNL4u8RvyB7XqdwZUvtoAZEXmdDFVgh54T7EEFyxs2LZLwkQCPGiQm6sKYFdlBIs8JVgAP7Y8P+
j9ycPK9rkS5ShH2tF3rHsipGtVgCMtH/SmNCHS7B2rmLF6Yhul0KqcH5f/IcEnwkC5vsg+Hoatj2
144GghCSm49HQz52U/SP1F95zFs0r4QtJ2H48pR8kmH6A6q77Qw/k3jwp0lMD/bOYnINn0TutsrM
wODlQ1NIGJS0nSTjtLFNV2li0yxeoOgRGlycgF63di2NkbyBrjQMyRX3wea3vHtH1zPo38ZTODhR
+kl2pJy/ox5MMbAtzHQkH9IwegvSt6p9ABO+8/QQYaiyLauG/XYn8WPjf9bghyBuM4D5f2giUnZN
/bydvtxyU7UFLtsIsPBgjmeiH43PT6y0n4BGhxpPCKM3suJARJuYNOFzxIxLpijj36k9Woo25VBd
LGNQ/9OxnT+ANmGw5L1tyqjHA3Njx33RtBFWqKkV6Wm04fV9iQ5eekPs+3mlHRcqxv9mSsAgXLxu
XWSqrRSUJvq56RXSaTePOTYkYQ+j2fj1PhfkPE5EvMNjq53CuUZvzGfaV8zxGtJELad/yKQtYPrH
8rQHLizyFDxymICTqdG6MD3CeeJYMfCV738ST9ndXulSLLcpNcyZkfvvghj8McqpYN/VG57ultJm
QN5iLCjZU6gXhaXO6qEB8KA9bF9GI0/TA4H73Bt4NFUAaYiBUQTktvugb3O2a02Dq6Ou+qaC43P/
ioO6twLtjifO7MV18lW/93lbT7+Dbp9CH1V4zB0gBYlOcJi9r6uX4SKPUBYqhgYOQuLQWEn2qkm8
NpPSVHdPCZIIS+3UTfphNwqIqi5wDIrfLexxVXdJ1ZGLUWepm/6paC1mScHCvkX7ffCpD15VnBp5
oOuh81HJW+IonCA4yvuGyA7S7ltY7/NitGQNfb0jFjZjAxiPS1YeeCjBnzDEECfvrafO77AKmwy5
4OcMKO+s2sdzjlB8INsrNdwABzljRrDBDYGrbcVEYnw8Z1yzFAEpoaWItkaP+j5ly0aLEoJ6GiUg
gsIQ9C6MxCzyLfnSWiIQPvYQNsCbLggDk/z1rGb0FMAwcs9RmGcwhDVxkoZ5DafNWOiVAWRHgeDV
r9/V8pLXyH0neIX578Ax5aM5OmqAL4TqJOdCfxKlJ+pa0J9vSwjJkmoUiqfOryfvJdh2MJLvOrai
jcBDZfRBlwhUqWjHm2lEe4uRvLFd0wgCXwFemmQ/KXguU6trn3KsC3zDa8ogpEhQqdRkeqfO3O9f
tzKF4N7Qg7Td5anb6orFVfMbO6y9aVpbSY4LRXx2tiPYoQLiaOf/8KycdEksJMHMnVXxTT3H39xv
iwGRofrpja0KgWdpKP1tk3Y746Ysp89Lw0yo5Oi0vLiR+8lvrUY7szMhWE2yFCsKk6uZITiafsVz
oF/DOZg/Ax6Qh5Sijz5+V7Ke4clDeS9pb3dksh9SgWPNpO4WP1ElocdpmbyQhw2Hd/t51bUmhWHf
beztvy+nCIjtxU+Xc2NshTTnx66WilBEU1T9nsZ9I4Gg4/450j5YXemY8uF+/kw5DIFjl81WIRQo
oHsOZTKhX4P+0golmAdDIoXjK0GjUCON3RItAdSVEgMLCLNcfsVbnBR4xiHo3niTOS/EZl4Tne6G
L2V5OKj+58Kz8Gti5Q3ln69EWam4QhvcTSXZcQTrY8xK8YcwQGPY6nk6h82W9tii2dptRb9WrwyG
zD3qpXCBbQpR8g3quNJtlDRFqzjXUsN+dqaVJhrTtR9vaNu/bTWkpX6t7LR2+4LFFm5/Ox5OH9yr
s+rzSUugAa1C/9ChrvtQJ+JlUquQlgxjQ4rBDnH5jjh7W1cFj4RK/2muvC3AzIuM/G7weYvg0Mi1
E5rcit1vaoV2XwTDtGO2KeEMVSUgHrJXIZD93UDV4o01Z6HjDgnzCE/LEAuDMKfonrz4JKvDCtc3
uCYb4mX6w9fpyJTYogTncezBtsB5VzjtAyIkwVU2b7URYhHHnx1SIsnfD/kvejD0H46Tm2nQFLAq
ANg3ruCTt2ClQgN0vSX/3YzhngCyRfuADrMuOZNp2y0OVq8m7AMG1xkXAZLYfXcI0wmL42hLi8qr
oiuaghu0kC1V9zWscIre1rfADVHDKC3xILiio8oZ042nOj4uTM+ImGhvDvxjHdPvdT+6Liuzs/BN
dgGatAtN5djiyLqgJSko3gjhUtXs1os7ktgdXgMZFETeucLhdx0zdsyNkO3kyokgZGJR45S1uPfA
yhIY37OghphroxBCK6g+AVqFuijp5aeOUTbcNmuKqGCu2OHu+NOmHWZcih4QVtUS813uAEE69uyG
5c+/I3CMSolAb+Vs7fe7zYIG/381Va63lYP7P27LyEJEReN/r/icujYzVnFIjfk4Pm143ls1sTML
I6d47+4GmNv+h8uWrad53s75AkpiCk/mEvXplpdJUUqf1UloXZpENO1A7F/A28gvVlnBg0G952FV
Ce9t10pAvxFlFKu7XpFc3PeO0uEwAVER/eFKKTVU0GNKaQkrGD5Lt5KvELjGHYF6XH62YuR2ZjVm
atTOlcsAtCoL7Rh9gvI3HG9l3YUQPl3+diOoO4bl3FK9OXS/41hO9xuHzja8Vji5ssjCNB/pZja9
j2DjeUbgQd7NvnPHDq7RN2SdcTXiVDLKXslHA6kw2oTMiMq6gsJYhH0RgO0TqXk30f7vrTie3WgS
YoK1JGAuFvR4z6pEw7xyxCTd30GQ3RYjV8YvjnCA4GMdFbnhhu6h36DQb1g4wAHkG/5m7HIgGGSS
VWHtW7Hx3lAl+wMVdNC5ceRahwBV/jRYJOtqftNCu7EnfDZJjbPmH8IqBkSDtSqg/sUtOlKklRXZ
+PaUwZr3LDAZxqaWxJ7SnFXt9cCfrcdPTF2Jgfm7lt5gI0wsiLH0GGQxFqrZDiR+MvVgMudQhw1J
/b+nGqgGv6HLWbc+YF0eRNTB8RcAsYUV+d0hDb2PhPq3/pVFcmNGk29/K0zlNuqc887QQr7fnBL4
/Cp5AxyQZ60RDeKiGWMwIDHVHmebOWbKenBkPlZB6WgMbolf9N+MWZWyyvauSzeZ63nzHaQCTisd
blZv0dBTnImZJiM1kEbsUmFxOWcxScbEzo8SIkhoeo2ENzHVGb3U2kow4WdM8elahdbLOVfBuG0L
PKvxn4QC8TA67QH3/f5jIuYIzpb21Q8lctboCqFveZIjj+nFw+F/SfJJw7OEpjQ6EqG3ooSoALea
xmV4MqLZH4voK8jkqysvbWm5Fcm9M75xFsy2u3ss5SRG5eLiY8WFL3KFEo56mEP9sNFzSkFR7hGq
2LMFCC57BOAnTAO2rmep2S44QMpfdLJe3UBPQit8bttdWL9WZUy0cQgyOYh8ll2L41yZMJshSXBH
/2/SBOJWCY0OjalpiGn+74lSZ9B34GZtOnAoshS30XOUm7SrBbDZkLHw28GYDGzbjPxHM4Zc/n+C
Vaw0ZYIP1BJIZvfjM36Ft44TpoP3rfd28c9en7jtC+q5Rh18Mr7yy9MlOMiWWVaHBklFaMOEo83z
SEHHv5L9E93gGuL/B3BV+jQ8LDfCmCqrMDWx+723ofsHrWTa6sUHlg3Q5D50aHl1iN7vKB7zqgTS
gx389hxZAxzS2ZmIa4+aqrG8gPc+V2NJtdU6BPqXZBRq0b62CI4FnyhtRe2TuJ1RC6jnBMyIBBte
RFgZTeE8V1F5a5uo3UJfXNCwmXgHgViUTWDWfamikZftZbUbz7MV3skRa3Ocoaed17FT5xjSjoVK
C+aDr0tTuYVSJESiQfLgsa2vi9+hQerPtsv38nzTNECven1H0A1nC77yHmEO+tsXWEXkgqc390Jf
R6c9gfTvSf5GLxOOw4cN6Y/awnShgAgzM89M+PJfPeqDjcHTYQXjooPNNsqqt8yJSvM0Vs7pNt4Z
/ydnnATnCNh+LPMG/SgEgqSXw/NmH7izY3ZlqZyIXngEVTQD29l3FPhU4zJ7btuS4xGNasgr853q
r0O4brPumyWoMOH3HQJ4eNnHRV3/tfO+c2a4dbi+fjjw6WyvbG9ML906U5llcFgkSBXS9ne2Fknz
qNiDIIg+dt6ZOUsF5Eb18juE2PN6750hSrrCD6miEJzGt/COnP6Cpl9mjTl8VlwVwgCqXoNEYGJS
Jl111FRfZVPXbeEpkie1Voanxd+8Er4WGq9CB2UJtA68tLNHk9twh/6RNXRc/qAcdr+Y4ptZvS3b
LwwEAAThLRvs6vWIQG3WqKCjWWoSS/gCaa+EsjcWO6bZZvQOGEmnZ0oKapotOsZSvis6yi/WQ4OY
TbXPhjsw9Jt+WCmcs3W8soz1AS2cYwSnTIS6gSrZnK4kW9XfISbYbL+yU533XtGSjlMqQGZHaL1G
Q8PDRp9tlSron7+suMGX8crYHEe6p4HXLNukkzpGXIXn2U/Ma2cdrUBm52Mk1MsxcdTbGsVAMtf3
/F8cv+Z09xmqnzVgY6F739pXZiHMW6n0CTM+GyVb1VFf2Iv93aTFf1DVZaVHkcaxlY8CfYh+DEHF
H9kP2QVbBxTV/QhQP6VQd/L2L9MEFPPmkW3nc+o64ola6VZicxFeRU2V4G2+cOF2MZGM47IYYRZt
Hiz4OIaOtXquCh6kwkS1GM1egImc5E+Ma2iHLT37pT+MGD7mfXv8l6bHmOxHYmKwEx79+LEoaF/i
3YL3FE+mibuoLaHSryqVmIyd0Q5PgSsxzrpYGDFvzrqWRf+HbBVAUc8KO2YECdaf0b841zcWjOcP
X1BP5zvbg9xelPNmFgNEoJmuqUcAr5FGvptLc/quldvwvw2xtRHKCIDcWEf7wjITW7hNH62W4NRk
2IEEcpEdBioUd5kMAxfIdHqbJgjTv8MKg9yP+wyPmG4ZVsjw1ARpZNxAvVGqiVFia3103VK9+gmc
jFfqkl8+yXFlLKcJbkm3Dy92MT36PxgljLmLB2GUbEF1c7+6IpftGSfrgUsdyNpW+Civkz3Zwcih
j1XBc3MwCqSn+ytbqrdsVG5YG+cLhruhg5YJbjSwP6JVoOr8H/qLdRYvOA7npOpwlefep74a5bzx
Zi72DZW3gMjrhxFleh/AhDvMLAgArnj/n2jA7ixxdognRYcxMKLsGGEyEuj3C36IXkVe5Od+vtPo
jTmL4uSVnM93ABmOzfugcZhJTviW7SS1SjNvwVfh+W8YI0u9N+1mcEx/+Ghn5zrUg07/2bSc7Qo2
TS0yBjqA4V/UZgu/wALfO5Wxu71TqpPawasPo1vTs9f027fPKOVlKXW7BxNDLUhwJY1V6u8gwXFF
SShqRRltQPwkRumanQioWhWHYOFgarwG+vKWANaoAgs7S+p3cRZsCq3MqBz1pHI70AUF0U6oe67z
h2Mb43QwSIYwHXfuv3pfDlV+zDn0+4A5ayMJpKEcdzLifIZCTG2s7+e2SzlmZcUHzhWSzRcLEwDY
FOm+g6Zawb3Zw2inAv7ycFK8hJ9wr2PI62hpLmuLXWPS0kQTnF2VfS9C2Bntl88XFi7ccX3PdSbx
RhYYTtyWvuzLBqNtFz7F9AQndEMgsIAKN2Uth566ym+zRimMdmd1B43RjYZl331x/g58GG7lKX5v
yau1rk0GTOMx39QHdeFpQJNaR4Uwe6McLLK6dyYT2enPoJlJNzaEWRasg4d8jj83+WwIjm+6uMtP
0Z5KJLFUqW2EClp8M4A8meNjb2ruiuPTcjW10D+nTjn37g+xeZMFJn8AObNtwEpqfvcGsBuvbVk9
sLpRZ4UGAds0k+sWzeVhL7KjX7QfxnsXBpaeO4/h84akvQze9XJj3ACPOcrWksVF0e4WXX86Vbt+
Z2NxuGQ2sxaAHLbqc9VgU7Gpo2eiN3ffznq48GjeWlxxeyb1oyA/qy3t4Io1uCY7x00lN9cSYnJI
v2NVN6W9PYii8VKVRbple/1BOattyZkOmyfToF80/uHOBDirMYsG2qB4Mk1YMUyjYNUxaI/RVPJA
Cguq7d84/3EeQxu3aKvWU/kHsAKWZ3axwli2TeCQWNOGUV9M6pdRWFpukIcnU2hY+0AE0E/R1kRK
5/M4yWldAAqebU6IJgVbx/x2LGEiRGeZ8Q/W1AWsSn2pkSrpGWqLotZe42Uk21TDlWAG/sku7EKW
BR9+foOXeKTc0+Py8K0fnUkN1BgeCbFyYQMQAia8RkRmi38XRbYX1wAVK6QrYuRytzKXyW6Vkyqv
+HU/eNItqTuc+Mbj3k1iyGzl0T3+mX7ECrfiBPF8diZSYS+5w8EeSDuQWGVa8nURIXKZK87+cUSh
tqh34SE3D9jYIZsFOMx+f4azjWDI1hXfWncMHjD0Sf3H1cgCPOG2PphMY7ylAzeHPSGkh/veiW//
iqA2rNk/s9vw3SdoLAWYvYr8kFH6GS+Usq1pBcKzE5kbqbEvNe7jwItDtfO6HPCNkxnWmmnjy9Go
p9ItotXBxt4gG7zbrwF0BAkditRvDvbTf7F5fbv2Kq/+HeCouJhZShdR5f4hnfFuJeMUdwbNV9WH
ODygkSE1X+zw0t7pC6F5Fx0QN9S4vZAa3i27nqZZdeANTqcQq+e2EWNGQDaNPjkyf/JF1dfdQoyv
UmOFSAifwRTVwBJfrCOyq2iE4vW9p+8vlloZuogjt4qqgTScrhMNe1A8t5uGIa25GFJV2b7FzvwH
MUulenHJS4V8iM1M76nr/8/JCSJ0s91x2wbH9UTC0DkX1Pq+IjvEQD7EfKy2FXe94bVSSs1QN2Wy
Rz96q4phG93Jw6GLwbbup1t5woftzYgkVrCkbsbdsZF0shv1py8/ySofgA0hNazrE7m3gqvB52te
cuWSI+YaFIYu8R9s5IbBc+za6V+ftvduMLJgmWm+SI2te2cfNNR7RkiRsUSLYjIvcosAjk2p3wQ7
UoonztljLDzVimyyxQBaEJQJSE+HFNE23hSnFmieURkK0KE2yRtp9n0wJ64Hfxt2keW81U9mvsSz
LhyEdjdzE8xx5oP5hGzoTY+kQwrEWErSG0jPDTyNR54DkP5g3Nc1zU3FLvfYvCiE9crMFhHAmYwq
gkhA9pAzZ2EUuRIY1TP0i4/K7/So5FaGSSSAhMPs2wf9X1t8NyNieILs3RpshLm2ttcvhQdkIuta
3BGhnVhgC8hmJqfp/UrMMcK5DWT2/p699jv4oFVPrb4for+AQWsi79kPJZakmc91bnRF+7QL0JSj
2r4EEB0zvcYjGm9zJ/KroIz5vgAlf/Y8IxA4ct38QlHfuAQhZM0uT0nwaRwZZu3tmpji6/jn3DR/
mERowdSNgD9wth5QQ3kdNKV0CsS3F73Ty5g1EPQ5PSx9O54uw+1lS+VPrtm+jMrHDQuMCo7nPGQ1
3R9gj1mkSZj6RHJpRk4JawXfKc8e5wWDxgRYXpwM9nMy6ohheCxUZdCJYAY22A/DW87QUuU3mOji
fI2AgK6aonFnS5rLpZunN5uW6zJ7LncQP+/4TVEGEVQtbgyNyD5A7sXg1VG/1iAHYhvF+NRd/TDV
Qq0YB+l8OXvEPGq9IcAx1f56wnefMWCdw//ocI4tJPdQ08f6B2TWp8i7bMtr10NaHnxI3sBDXKVj
rpk8fv7CzX+NtTBzTtsHjl4QLI9IxhjKil2nl+tpz6+RW+bAkdEEFn/NrkrjFHkNExbrKrALAWm9
bJxB98yTR1Eul0zBq7uU3qTkJq2NtYGM/zv4OcqydiVO5yo64qGwBGrHgPbC0sGeFqnpKEAdzdyv
wb+DTepfza2LrdY7fDDCbhbl4eLLqXw2QSH/hSP41Y5Oj0tS3243SwirHR+iCv8pp5DMnI1p9WFu
yi3p0dubFMinxqlqWsrctG54UVhT/j3M20hTVmHhzOMmAS7VDjODuzAdx/btUlO5uz8mzYpS5XDt
Gf4wHmQduz+gE/1ApcxyGvjJ0oua0TZrWG7ylzswRgnAMwtEkm4B8g9YewYqdQGx9flBH/Kr9x/Z
rpnUc63DEphyMnV4NEmPrHr0CzoipXg9ypWOVvQd/6wMWDeYccg+CyyAIXzZ0WF7or38Atz9FYxG
JmmNteKsjWUQmyUE2mT1fQTbZgh4yPyDP+Kp/6Z813rSCQfq06Ez4OsZ4/2qBT+n+CA5lz8METbt
xDfmiZyQEw9aw1bMYmvz3t+CdIZtsU8zFWJERf6J+3XeBuSu73YrJlDPpdYcbW3FLcV/nzGBskCd
FwGxM67KG51cPiupuQmIJwizTisQdY7sYnU/kDbzFid4yukmxv6KFj8U2/pVCRWrD7eM32D8daks
cK3yexgcz9JZm2N2LJWjgf/Aohu7P3Wq4fq5kv8Q601E9U51+FE48TtA73SFBluOjnl4+viFMuEC
QL6EnghIlnMV90VjdvMunX5XXmxDWnzqG6YogFsnNkDLnEbPys+xBnVVojAB2lubX1Ncu7QItU2O
q/IMsxavu7DXh0fLoZ7g9c7e3llxdg+1tDQbi/UxW/559XqFbSKegew+sjjHbJREJeSJ9iQt21IQ
GeMtAmGYdtspY87vfLY5b6JL25LznPzemdJ7KYq8mDD6vbkmnXma2qm3HJ/kPAimEkBgogF6see1
EnZ2vyHYTUgvp+jeQFkLSGcaeUKdtPWduVhrKWJ1TWEJ5vT/RN8T6ys65zvebPx4L2K+nobDPcYF
026izGi67DkC7AKUHM6jCxKI6gGH0+25hfiQ003ALlsaCAuDh2ExfHr+HngtMu8sYlCN7r/sdjsr
/JtAuIdF5h8xWQXh2rHJfzEt860dEoU56FgFLwlHtUTSDKO7pQSY20xkkgHBo7lxq0aLiJ9Y+KJR
h/ei4R4j7Vx02RuoMiHQJFtJvRdEEHiWeFXlpqtZVdpbAflW2Up4FO41Ioq8lzXoJUm/0XfMASsG
hC631JFqqyqBZsJj8qceKuJrcIowXcTchWYsDgxV1thSR4qqA/2S8d1DSheZsbTEEekrOM6jZeWy
7ar6Y+u4BH492vMcx6jQ0i4kHksVbeJJ3J25Z5/JbPfq22Bl2HDo2O4d9TGLas3GJvwQuRQNfXr7
0zMs9qTCnO20U5XDCMZ1RcGzZsOhjbhZecx4JOM5Jp341vjkLGE0GQyIIpnPwXmfMZlv7RQbRk8y
1mLzLMSvHxrupuYzuAYh9NYhYC3fWZn0bvMVT2Hd+KtZvY08EC2V13MLWG4Bi62RnM9Trav6dRhm
l9aogjrA9z1dHhpXlGjZOUj44yT8hdTwStsL1ob29StpgQ/RpMHhYGOZ44OPt0Wsqh52Pnb/JMbH
WUpYs+mKSqnGNV7+8YRLabg4W3tmppKUFHUSlgFqekr5xaPp9fx6jTMLyhFd3CsAycdA8Z3Naszy
Y/JToZK9dJQWcn/K0XGy2Y7eLkQoDBGG8snRPcYLPVMD5LIDjH+fvGmNCZY/IAnlaDBdIOrWx+2w
jLhmQL9nukHvrBmUskqHh1+luhy7lxm7IlJrEAc3wO2YEFTAr9dQZCPI4Md8+VvFKwQQsGAGe5S0
pUTe++jM/tc/guSIYlBvxFxmNZuPrMjWqnnaJa5+duJjRZV0jn9ErcAHbqYPJ0GbbiW0v+WCqIpb
iKTEWxm9xnJo9OvoJzfePK4ZdQkhl0peuEtp5ba4CUgemk8nPjuzMonob2CWHFZJ+M5YWBsw7ouL
rChrRGrtXcP3gwc53U05fcm+1KfbcB5yNhFIohEiOYK7E1aOwgOsf6DuRGGh6ucsbepCc1TnXlq1
BcaamvgRV2HP15a8CrFaH9vQf3CQyiyyB5WerTn07FXCUn3JtDpE6Ga3i8l5vgfGu3of7KXgmKqJ
43P2MQQuwwp/RTx+5ozW1U0J0tLoG7aTRewXnJivRLnSbMaHqicGqQmD3AR9EWd2T5Pc86Qg6sjn
k5KHWl/VLFqbcmwzmA14S4I3tNY7z01ZgeKPGATROOUF2QbV/a5o3bCbRDRmEG2klKKqvMkdDF6Y
lIM0I/g8X8Fx8HqvU57sskGxFGxa9/lnJ0i4dvmdbz2KslAZ1njBupCFO3puvh5e6ghNMfvLyX9m
Icj3tJ3dIaTf5lv+00UVM7NV71xla9M/l2oSqqoznC1Gm7Jx1zLMVSm9KUdby2APmp0hGZj0BgNW
fgFEDCHRlJLdLm6hBF5oWlwICrUeRPLt4TRwckineA4Qq9b/dAH/nsc9wYkZ38synbQc6c5exAck
wXls36DjyVL2y3eiZ8fISZfOhbpH6Sl9a1rZ0K7V21UDYAXVFsXMY6ODajilUSqXUO5vpiZrBOQv
Qiu2mzbv7S8RKtWBs+5QsMU+A65uY8p5IzeN2loU8p0SweneWrO6oDWdqt4c6ADnJQfKZ086+Te4
0qx/dE/cG+r7yiBKNl5LHqBbiPRr6JxErML8Z6hRyusRJD7ZV99Wqz86U9XaAOpxrE/zhizcTX69
wP0GBpqbvl2U7czdq0B1obYxwygxxQcljQQWS8zCYUh5R7JnxolCAmIw+yUJ1YcnXOHZ9+Z0caq+
Pg9TGdzs2fxs3izM2ysn2mttJ5Y3y8uMnYIYnLbrDPDQCjYyk2GkS6XOo6IkYjQKwqE4cqfqLeG9
T2HqD9ZxQQOk0tBa87A9UVli9TOtdUVEzJ2uegb11gYYku2sKrs/MfdZBCqofnwWsQt/CKaZyXUQ
tRbKzROGsdzZmdgkGdXR42nbkBtjEsyxw7QTnijWhRKd3b0lcS8dI4VdVTVyAupicyByzBmDiFYr
kArs5qHRJT5bxJzfSwac/bj88FcJXuRbJg3Ht7jgpxz5qjF2HI8hfTDKK6ifOnQR5ZnEOJMpy+YJ
rMhplhLfZxCTp5XQh2FsYG1+Nd6a+96MzR3TWEB9SWqVv44qR2y1lPpdmMxPoBChvb7QQKFKAbcp
1lrl3sf37Tt92aAZKrjnGX0tfhRZ425mNeASlGYON+ZGte0GUU5As64pvt+V06P/Q+0CTdqcUdBO
MXCIY/zYDm7vNvew72yLdwS3QcVRa14ummIpRcK3tW+o5cLuOdpfPYcJ6Kf14Z7Qf/7x3VMf4gHQ
wpKOLmdTvWPea83Jm9FZrUpVooVNT0EVxDasV7iV3qRVEf1WQ8D+MAWIvIgr/DuB4jhRfSEUZL6c
2riQEvw69uZ8dVJCCsbtuNH+onwV/FCGnEPAihNTygszVJfids0bgTw95xY9vB2anxI33OcdQmLT
acUPmYd2WQITu4iEdMj6Xxe38PRtjeHrHuEHVd+Fx3zVtrOZqKsN8VUJrei1nc//Qxy1zV75V8zK
t5N4OeOs+zWvuqbmw4zwWjuNsF37gM5nI0/G0Q7t7BcNROPXbASmkXQQeCrYZO3oK5AEMm/eMajD
tidm+Psl0O71reLM1J6o7Qg/g8GXRjS76h+SoJEzMIehpFqOAquuKq5yroLfE5FmHj6R/8DVm57U
o/ZH5h+4Zkh1AAHirN0oAeRDdm6LNBp7E/WnTB34xybxvqePFwew2vLmM7JWilOpOuhZh5Fm04aX
9mGDM4XpTuI2sjPSpHkn6VDu1sfBGTgNPIJxSYXBxCHLBPecEogZdxcJIUvS0/gF4purclnko373
N776KZaNfnlFnWRs7bWoREmvBtwLI98r8EdM7YI2kJKRCtYWFGb/ATeR8M0iwo4iS2Tr9otz36I/
pakcZ3511PdwAbOc1g/2eGddh500tNK+aDK9iFg4k2HuR8yhab81aB0Zfu6XzZKIx/6DbdkmE64k
UoI1WgBuo4skq7H6E96Y/3VK6vPl1Mycj2R+vnR/8lVQOF4c4gXNQVkJQcP75VybbKrXHm4Yq1Ej
hp4/ZtR4hx6EQKWbotZTeWXA09J1JzAndi1GrCTqqNvd/iI2ooAjCbSwNTeck2/YYRr4a7WwQfye
X3wrr1mFH+G8Osu+sCJe9KHboT+YtxUtXWKFRJBrd1bgJI6vqhHv0D37YMjtzO5sOhhsHC+SQPii
NxBsUbwvSBOdYwXbrhynRxOT4jO3QBYHoeKMDUde13+Qyzb4SMG/85tC8ZrvMoqxhE8VKhk1NTIh
/g9/qM21y58nLoBF+hl7c32m2P/BTMuTW5HiFBHtGo84zxT5GC8iAIFqRDnpT6wrwXoGI4q50rDE
giKM4EqGCCUFxpbihRLBb8F1bIzRcwjIm6GMhhYGZIJiYb0otuUhBCXvgfuSkB4/eeM05qj45gtV
FWpbWyjRCt0sI4oBxn9sKcVXG1rpYclgt6ZiafcLrTIuO6ESoUjIPggsIfW9W4pGa5cHqoWm2GJ4
FAfPQ5EZHxertDcKubaMMWtsa6P3J0/ddqWPziwwhWpA/Hj0yBeKwWxrNG8+E1pDWWtLCbaAB6o8
/avxYqirW8GrFWJ8HUM0I+k8zePUgoqSwsPRbe542b+VbZV9KTg+qyoYZSpxPF3gyykpUT+htIC5
aaoUtcnP9zGkWpGKib4vvMJ9sXYhilTeMpAVo2yyN68a/qVzsD+EgFerXmQeeZTEjXkY+GbAIVVQ
I5MYwCIL96zZyph437Aa/UoMsPFbhBqtRi7IMMFaa3l1e1sZ+t4CRJiiwuzNHR+bSY653CZfNUci
Ds6zq9QyuG1hqDKQJVNrzl48EJcNvmrnhc5kcFJ0DtmXjXSo247lfq/EVhlnOXqIc7mDCZJMqQe4
0Wv3KVnEpk4brZ9dbtghlB2OoDtl4JS7IOnrSbQpGV8SaxTau+bsa+lycAyusoJOewt/3I1dDrhv
/UjnK2eQj6sxx4ULiqGSeWc5KUJSVCAXynaBLL8ZZa1iUBHlSp2kTyTgfUb2iwLQlROLYWleGh5q
iUBJC1n+X9eVkWVUJrTRjrD9dPods3EKFOK/2roilW5uE0qtNnVi62tmWUeIoC3arteZNsshh8yW
brDjT0i/4lN23ldwH/d6C2DP1lnCCB8scVobHjctaI8iEEPSlIlKQSh1IjLq0NRmOEd+FniQrEra
mR2k9b1b/C4UJ46oXm9lj9rSs97FFxJnVP2GF/xbKBsBYua9aWhjlroM42vm1ox0swrdXQpWaDlb
OYrg/f3aP0xmRHkEniOkhRX/OSsGmzuIIatk+Di1orrrmKOO8sFt2JQHOc1fgI2gOHiORm+Lra9P
Kvf48ZbAir/vnIQuovKkx7Gor7Zg36K6ni6dEiYqt6d8XODNizCXVhks7yN/MfKfMt/rzldZKYLm
Gj5aYVZ+uPUyVgv5xHK7UL+f3//QyzMRtc6z2R2avl/CfYFHWEKV+U5s4c1ox6UgH0d2JpxWFVGo
hwjWLfV21V7IkAhLyFc3e+/qyGk6LTGBJNu/1FzBnryr4Tqw6xeon5/iaz0/cPErDkYQsGGJWvDD
/xrotccp7o5eT1HL+EtAj4LrXWKvEXEjzsCNJJR+gg2Qggzj91TEXCnAl9bN3KjShFeFYHM92swT
8lUtVDX5KUvPDXyKevST8B7L0OThGOpXqhQuc6hebVH/Ej7ydhYMbRbd0RQ/WeeVe1Y0+C3CnK99
sGUYyFRjM9OXyXAkXM9At0Gk452zTS8EhGHksc2TZVw9TzcDsSNHrm3zUCO8LmYjnuCdQeKlkwZX
ApXagMFtIByzYx3xWfqZLuW17r5sFUA1IGzm959AH5NnDTxbkiXxADLKwOvn/pZo61ly8bBiyybD
i+YMs2TMg0uSeCxxTmVbZ5VPRSK72Aq7VUb/Jb3qF1YH1pFheUpLKdxhTitEvdKCDawgBRkFtHew
jRy7+MkooebuEikca/9cCUKLszD6LiAqV3a9kM4aB23Rjqo68l+M1zpOo2HRWP+CmexEr+E1zHWB
nMYrkBJJqaJ5VMs1N+cSZLixa/8r8Dp4+5ZGljo+BGFpc4aZcot84d+FC/v2ltN7YxFrfwsFkE+1
/tpXeK9dxByPI+q0rJS/eKL4161iRbqkxfikGnnelXgF66egpLvBluunXgdCQya6mBJczf3DIdv7
PWwPiIwLwDlCfG/YJW2qG8KGot2ExBJU4USCoo443cVmuqYdLHnAaKaOF2alMvB46gOJ3pYRe759
lnLMd1jXbGk+BFu8ipaF0HCMikdV+zoeTZTSJ2yk7g+5LeQawkspQbh47DkMisFGBHjxAdf7YUNn
JacProH/6N9WDP3+X+L0VQP7EocSELZEhdUDaxHZxK749G44wIpVms58UgZWiNFhrRlULhOnpZmB
f7f/AY2eVa4hXjUu8MMdRF5hbhTRX4IIxVw6qT/PSt4dFV52hpaQCMW3swGfMihkL6pZDf6wY3B9
sRQp+3oMBuKOvrR0ZtKyiCOmOKpLI+pskcztUNbd90IKy7+MUclHPxeT+hlamA8Vf3BOGOFETKNA
zTCRbbYT63aYZHnl+VCiuGneJjyHvXV8LZOq4GGNNwmxcsv5IAOpeVyBozwPe1B0cRSqyjqnIT3S
dst379bkHzIXf+ytOcf6Vd7RnaWM23wwg+LDWp6Yl6304gsuSq/rexdvXISUhUXLa0bbkTOJS0nf
ziYKwyDlhHjC/aUqpzAhwEd0+F2n++M5oQ7hcozf/zkO9Pxzo0a8P0l2i5gqFKKXCSZb9raJr2ja
lzg0h7K7+t4xYIapGbk41WszWgVA/cfw9foGvXKa2rWhXbleMYMmwW2vZ5gcNz+lz6acgD3dt202
uM99A5Qr4DiHPygv4+0JFLKU/q/5S77/cVA4x7EYYXLOUxpc6DRy2g2cqcqMTFXV9OivrfGjCw7f
aZRqBQghRdpZUBAgxnsGrJAKcpRKe0LZbgZZMeCRNhbwx4jIb5YVzoGZjNZyg7qelCXgcNKC1Vl7
Cytx+uPToGMwN+RyNyVZMT7bmEMCzdl190WiHuYttc6yZACv2n7jCnSH2nn0dI6eukS3rxNUA3WV
xWeIJW1+9dDzTp0T50ccvWRziJN00tn4MZPu7XzNuqOhHdZqpbOKEbxKIQ67VP1/uHntFK40UHCG
fEa+u7nq22OrQw68HMgeSFglpXWsm8paj00bx9H2qW+LbY5Yb/Ze4dzHUFgtmUrnf2zDR5isox/X
q9d0Aha0KxOKwzoulxsw6+7xm4Ffh/S8pPbQkjDu+WFSE5pjto6e6oIDN7mE0ZyoEkrmXxXY8vDn
Q9YLCcnDCbXCGHp85Q6xwUfurfyYCwlZGCrEnnvLIR4C/dsfC76jtTdeD2xnWrbD5B03uHQr93rT
zEYSIIAZBUU/alcNsXu3j5ZPw8R0JhIVY6Rfoxg9dG+nNbiTB7qJvMaTu5rk8Sk6NmN254RNogv2
VMYPQfPojBLn104QIlVIpbMWLf8YJz6gQfHrLYB/cZa/f1akisyM+2FWb6q/hU4+NUCJdhCHtKok
kTw6estvOL2oz6zkMmgExBo3B49Ai7hCTvQZCtfDZMfBlvL9T7/cweslpcxBITDeE9XN8sEQ8/+D
xqG3V9MMpeABfRiCU6SrRY7qsWRFWkGItKj6b/6NfUv4fHT5OkGvS0YiKNxXnItgabiuynVLHJiW
+or240F3m7ERYWEBt6k6aXjZNB7CMhE3TiZ1OY4ZHd6ZQKnmZb6Clm2BghuONx4/xjercH+4jTc6
cOGt8egEb7NCYMTO8I24ylektFFYi2VccOOgHlLyZUOv4Eza4oR1n0PorLcIn/4Lb+7q2w4kE3Cy
mjqC/JhydA3kyvnl0hfYAKEtnKrTIiF0dLdtZ7nVTsCPLFJZ8zOtULDnXr2zWljY32YBJBdrEj4H
kYY6EkTkk8LKQ6FZfp3jT/Hy0rInO3Xm9XN0/TPRIEt57cYT014CHZzaE7aXA6a0Vu/lqpipq2Je
Wpuw2CpAOQF0QA0Z6ytSnnICdh6RohgsVfnhvH46hWmG6vFsobJSgiCWmXe/GR2KUiepyCBKyEwZ
tqmAN1lR888Jy43IzTgBurbyBeUV1SyGgIza9DtjQIAwMYvVb3jqDbipWAPnNQCd5JcSHKAENMMv
d/2681N1VTPYl9QFYxijtrExmVP9d5fdqwIdk3OXA5BkMXhr/wFeigqZl08pO+P4Bf/PY5A6zSkU
KvMDN77QEbnj/4PHxvgN97iGpu27bSfWYR5Db8sP0JkRigvF4px07VFTN62Jpg0PqGazTkNtYD8h
h7VWShYeW86r4gUIlHoIk3iaD6bAni1gzkOCXlhrwiHi0HMXS0JPnTmpJMYCVJ1yha5o4hBSLj/x
zpDva7ksk8S+vcRYGbWLTIsqzP5Fm8dt/FGnon8A3b2top4Ox3RDxAUEKWWtm+T8722lk1Askbcy
OVAcW5+tp38AEtwOMJCdLtEQmsTFdeRUix/DnzCYGPUGSx/zwsQPRuZlXxdi4PumOtbUR+fbMV0a
/3CdJ0Y18Ngs/pbSSvyUZbz7w/E/MHZW+20Pyn7RxPNbd3NP0Ya8tiHCmjhkpcqZTDXWMg+FXUM4
UffMLkOCxBGaG1SYBhR/lHz4zkr3lnXQ9Vf6XX1nmxLBpg4eUy0+as2IoupikWIZ/R6Zj9cVJfoy
IZnjk5rY4iePfn5fz8ffhoPrT++feftQyqFy3P6Gh0YWah28B6oaubxGuFj76D39Q8S75IjIHMOD
mBvRyRLsLkB6lMDvrpg7HoQCXLUIAAoexrMFzcltFHZK1NKwZMZv85bLF0efb0zyPlEoPV3Mu5bm
ZEmVaZbpj2kzYd5ZeQLcURYZ6VQgT0PJP7+5v9qU9xYak0Wh1t6ugsCyx7kpdXP333D8DKTixlkQ
HSXpKLGx/T8kRF3U1/2VRnZXWkSr0lySKbx1vOccFmUAmBZgWrstAoWuuzk98GFZkHK1PedQsF86
e4DTHIrTBbq21XMABvF8hrJ+vw9ENew9dkNzTZQQAyhjM0utLJq3yS/vH14Nni5UfQaSjTbexwd1
zVhI/Vo4VFoMjlPpe614reqSwavvhPgoN3KXilRp1bKxIa9NX+7Wo3VSF6lMNRNzmLxd3LhtpVto
ZQawgA6CYJmBypbK7sFetZ+JEESzc/bLFat6r/+bzcYMC3QfZw5lsyqqqwhwcO7CkhHZjuR0fNBW
U1FuamP8+UAhugFz5ed44iJiIcX+04vNOk8icQo6CroOefjAROOVD3XlDpH+cbJlxcsd6oLjhheD
5yTfmY5vtRFZSbifTixBEF7pL7dUYBxjkHm0IBRQVXSgpRv2/J2TdNBvIMCoWNCahKsTlGM5Yr2l
LVk8a3SFun7Kd+IDyZwUkefHyffHms5KBW5DaUKv0xLzGtRO6WBUlx7lySWJXqAIzq48xiPOIh6J
fUkU/ziSZD7aN7KDJ/VZMebPSDTiZ5lPWNZ10HW84V1ydnUjA5f6vcqBBSTFPWiMHoPyHXwxZeQV
bZnvpSB15QpNOGJ4jU2TEUYOlghLyXUIxtWHxp1CsPMHMyqpQCbgy9TmUeNxSeBfetpgct+U+SpE
TVNq0xZgvdmwieBUEVN1aEqFlRHUDBOm8lwhEbdFzzXPVLDEOqIaVCbpNgHMfTlxlCPe5qeevyTV
S8k1NbVJxueA2zfPbXihoT7mBnjkKi+jyzy4kILUi8qRkdVNu3zrBJmmVs7kgiPaZhrFUBoyy/7J
d8/TxLtxtvtHQybuoS6M6eDSYEaEkfFw+GDk7DHJEzTUzgrnw+dFz/NTD8xMSLrRX8uNzUwnY+65
2Ttw517x/vC0BTxzXhv5zqdo/cWp0yHYjHL8YeOSBFqP78ICU4vTK4t9nyuLEAD08axJLklwqCaW
L3WZWGfoLmv9ZMMnD5iSSav2xlX2mCEZeZOam2h+Jzc10Wb9SacahPsOx4ZtBzemu/1lOMBzLX1j
KWMqv332slVC0u/1Qx+zN2qJH0Tf+2Nkn/6AEw8/NsWstAqlTOFWxcoS7p8CXYJ1NH5Zk5JvwkOe
rwzO6d6PXfKR2z0GYUtbVTSt4EciqFRr0NZW7lzkErOnhj3WIl0WcsiOnnDnXay65iULcfffmBjh
wN+HPRSSPvg7Ev2/qezReM5LxTk1kTYgveK9rU8p+etMGebfVdReUzt0Di+tQx2KFF4vn+j08Ql0
/qsF5n8l+SO/5Wgk0HVpSusXnLQDzPZi+rwwhD4OKYUixFXqFVcotxfogepzm5m/5iq11DObs5c+
artNLNiHB9Sqs5PETsXc5Aq82bD/Y9B2Xe1ybAWHK0DCfYa6JGrSfCH/IoDY6r1PVLfq3S3ZpKbo
cYybrpG5BcYTqyDv3pJ2LZGw5HYbFdUzjNNMxqdsgFLdT9c3nC2Xyqp0PJHqYkOb6enHg1sDlnaV
npigKBJjIhU4RkYdraGhWciYdxV8oCTOiG5GqZMXmEH5P44XQWLHJbawTJrVDIQhLg8rTAkKrxRb
e5GoXpZIbMk37r6tSljvJp2/hhUS3zG08dyDLiC5uITRQuze7Fe/TsNLdtyvn2HzUjCPF9WTYeAD
gB6uTT7XvoEI4zMALAEZOt7koIbe34AuSKRw1NvcZz6hOuj3jwPVLzABMhIAKsAzbicqaEdca2VM
Qu0P6S7XpYgluKYdODAOHUpMNOyvQvk3yUnCzIWP8yDMLK5r3/1srBJGVBodGQPn4f4oz2JrAPnj
U7VlFyWSZTGOs3rA3AVssWNtrQEnOSiqGwmueB/SsYDi/bUCSebNT4a+qFjSb4nMxt0cEbaf+gZC
FrNm0RhInEFRIjspLgL65yHhAm+wyjcnIuk/wtMDlJf3Nh+0upxQ7YUyGgCPaOD4aHa/f2+jOnl2
J8fW9vQZ1M3FhONQo8lVJjBGpiZ3dtUCnSf1inQflwsi9c77g0Ja5SIjKvBtxo3fBEk6xoewq4v9
zr8TPfi9pm06mU8CvAzqmzUZhGcTn+Tbz8pL3F3WaRlDSLaP5Zk1qKaotR3QtWHEPcHHg1dY10jW
OZ4weSKXWzcPwyezy89nQcJ+6t23z1cZCJxEeuS8vgU2WaXlgwJBIke+eDD5KHJwDxfR9XJqaqji
bl+Vc26SiUYaKGsxR9jNQnEqAahxemy2oGHBqHOVOuwU/p6l6MQDxYiLRe6L1oI2AQw7dDCVC46g
mH0yRWQ1frtl6zxpLt1MPT0x4nEfskTRqtfC2lIPFhg2sPJk3JaWM3URuRP2MoYdsi59p1n8vXFZ
vQr4Qwp6OOSfl+P3slnVOJMsisu9kvj4u50BEgYuvxkR1R4FhSesmw/udy2Jy/soXN7oL7+sNz+f
WXIkcx6SzAM8Gsz9ZMbf2CSt4XvPWUC8VFGuldYVKRoK60wTEmaI2CmbTa4CGXKc6itr78AZOK3G
W6BIPJDc7Ef/FX7ukSNeopMR9K9WaN5zNb3DWwpQRIIJxS1z4Geu81qclkO6ZJtir5atm//i0Whm
0l65VN9qQelZBqcjkC+iT4tAxzaz0sPnLXpFV8bOyq1Qp6DCuQ4XLgSISURZ6GAyBnlTB83WCeWB
2Yz6Qw0053hE2qXdCQ8hx3aaVFyoW5AJ9+YPdHBG+MN+MCz+9PaYWSjC59mNk23wH3Q5icL/dsv7
dNlX4ZKzFA2cd680G8qy7HBOTrOIddH8Ua3n8RIp3+0v+tfeWUcJvaXsejJqCqupDWx/7QMpTcr0
0QBNWfa+JvQyWy0OG7KVM7vaLI8QrMi+w4bh4Qli764qin08r68/OkcMiZAls10KdXycsExYOWMX
MA0hG2ulqufzk8Hozi/wkvPWsPgOOX/2ZmtRvIizCZkDuakQBDpbl1DaH4ewvyyPHAEobYsYbETT
bkw6+jmPxO7Ne4cgizW3ufLy3q8z+JqPuGXfS4XnzkUhOX+c2SriIx/cS5CQftDuXIkdJOt8S6ze
Gzxj+n4gGqEnMhsSnLziv4Q6uUaem3+3OL3T32LMkF6tvlZsbxubExelfUNLhZcJLMjE0voTUFv3
iPp/9ir7Ldl+5e1IEvFxOIlbzMEfi/LsIcQWmS5BZrIJPiP8k5HxmzYJ4GPrkQ0ogZW72fMlx7YA
UK7D9eX4OdMwJYK/cJgk8CpJU0lTmoolqVUmI4AH/b9+onMJ0lzmQD2dc+T0yIQ0NBZEyYPH87ZV
V6xFXeps+H/IZQ6tsj19j+gSTE/QQf1vF+660zSb6tCWyq150XpvD2ka/QO4xVdNQ6i+dHmpVHT7
9s/nFW//b9hc0C/ObXo08/ZLtDhUK0/6DX7vwNtN3PL0SlCNmQzYP9bOpDxBoAC+S52o+uwvS+f0
Rbpi0qc1OMpi3f2u2mmH0lEhhXLG7Qchsyvq1lK5Bx2ybD4QJJB3z57mscq7P7hrRlZ0BjS7plmm
fs971TKN+l5h5g4PXJXelNJEnrojB2eyzrKolUHAA/BlFwtOtlW6/UqcAFwnf6XOGSRgabHhQ/sg
UMJFdjgi7HBa1QF7ISSEqb/54RiQtnRmItT/gOuVkWR5sKAQ2r1inKlW09LB2Wl+yyokd1ycHjd1
4boFVT/xElejaqANdQ+5wwYVRyyfOZ1H8wvxlWx6t6zms1pxxWvrVdQDjvpM6L3oVQdR3Rbi+eqK
favD4ndku5Q3URILWQ5OqohMcvOYuxK3kV4yn0a5n3Cbfo/Gl8pHNyaQ1oa1O7iIibYwFpEiaAHI
b0tz/arkyK/ou3Zn6Kkqi9ecvdBdKKSb/vPYHRnzAhL7VIMTq8MCxDEg3MANiElEAMcUr8+UxIIq
y6vsWjAwh69PV7MdY9r0/CaJzDYJyXszvJcczXlRqq36lDPts7gjCy2VNx+mYTQvFpZGT1l0ftFm
ZuOYf0cCWbEOpx+VT1582TwJAmdtrFUDc7R12PP8yB79d6/zKWqxWkcJAE2iRf4O0aYs8OsHywuD
Jz/OunsIEeDL2dtuc3mXvdFymIh4uwJnbbZxRS1mLxxmRNyna6x4ASzaq+Kv1NZ8OXqlm4184ssp
EewY3YnJWrgDvdgbkvbWK5fsvOsbZfOBKrHktqxqoGkNAsrSgv2itbNGBtXwEguWaguj+NreOiSu
lu9sn4Njeq1uZpG2UUg6RXE4LnrHYDGJuaIGnlaQ27AaQ2UM31f5wIxONzaX0Q62dIA7gQZtYay2
Mam3DXEmDqIeeIIu/SQmmU/WmBDCXZ1YmMIFHNFmOeWquSZJ5Utx18eLQT+vkANqhtrjBwandjGI
ShljkTeDW32r9mr5UqDd9vxtgDRnnkLmvTBJMop63uoMhTaWfArsoHtwXerPcJ+WXIJ3AKfiL2+/
CofhVwT0A85L3ZUJn5Il9bosmGmUq84Gy5qIfIKG9xtjDDkJd3hlQLX1BDVdhL3qjMf6gedQrLuO
HL75X1iPBg2X0CqOpd4pbjPmLvfjJUcKe63e7f+ShuIz5kmSnNwQIb+33wmZaqfTNyfkHohI/ATF
bTvVoHzJW1NyjwSpETw+6IYCnTjwLCjT+HLfFCuAL7Jiah4V7k/nkPTMMATvicDDFnLHzwTxbxW+
Z51A30KRV6SLNltPgblyM6WIPLPngGJtKeq6LTp9bxSzTt1EnCsnSB9rz5be5g163wQSespfqp0T
hKNeugTxXBassy0j8DIcpHZnHJLYgo62AzA4yRdQnH9mvZXxukZphvBE9+cxOybTbAFxelj42OEI
0m7so5Yercy2BV6+FlKb17/KYZhad0GnCRzZcyaetwximyznKEywbtOjop+fCyeXZ3aK1NCZvEv+
7FKzsL2/jUr76lmf3MCe5VEH/xpCNvrhjwwl+o+fy2qFsaQuao+eU1vVY48fvxp1GzdaDHeWkon1
0Mtviw8SyjlBvyYFLLIWjyHt3GrBiLa9isUDpespbDzTvGOMLMGBnLDN191KRONEKpD44u/TbGOp
IhnEs2uNSK9pngaZ7xKM4tZv2dHYPm3ueqXuQ8dgOiIXZEJyEw2qNNTXse2ZGWVwlBmo3j6Z1Pn5
C8gLNk2iRvqr8LLiUx7muXgmOT3vh7pyhEBwUcwJ4cYS9ra0+LqTELMrjahVwBdLEY6T9j3VgJnt
NXvaSmu57bEfQKpkVuhGmRvinHNjdvMqnsUfeI82asQlauYj8Ri+HXITxmUfumIxwc+iqgepMktT
sIlWQBgHxwzVJ8AUVaJAUW8OcVOhRnN7l9CkZ2p2TNZnP5/TdPgSunJDwtYejP4QFjaNbQS7p3NK
B0qrnXuREOoS2qrnU90w84Vn6K/AZtQAbUlQC0rSYIxVvKcMzm2KDlmeye/O6EGchKee6aTePNUD
+C4KDSWpI+wIVnqYLpY3v6Kj1sBoH5d/ckt4LshB2OHM37MHjWb/qJwV3qPcdB0lp1owHrbSW8rm
+NqnOMGmNdkUUXYLtiygYZDWhchbSgs/RIazb6O3jPpxe3xe/1EcrTlcfWkrhOp+Fb017xGC28hE
qTZBnbrGBqVaOxEThywQIqdGoQRcP087O5a3AYRrYvaFcFtpBIAymZFCxbQ7c8e3fi6/TljlkjMi
3sOGsHtokMCdDER8A2L3RxYDd6mkefEEJAmlsrjT0PA1ARewpDgCIP2E7FvDQxZwKfvflfycZ3G8
v6XkHpjS/GYUC+W6quccN1gk4wFPb7bnXQS8qFKoDhyEj4neJHvjtYYoW9Jj1d1BJK8icD9rs7nA
EUogJYqm3CQDPiNN2AMHkZxIIGc6d/Y3Zf+hxCekZNHNdRD+RDdpMJytrSuOq7QtldRtr6gvG7eA
byQgUcLC8uvmUAfaUdlD95/yNePij476LiKdktO+RVGPlEXH3RBi/ViV66lLMOOZyUevqPRc1mIh
9wBvdKJM+GyYIfoEa29qwrwQijej4RSXFSgkUZfnDvPISnadITnbEkcVuqrDmFLn6IUr8HkTCbYe
kjvXXbd6QV7vVS+tTNlAtv1sMXVQt39v5Ou5TSBerETvxSPdTEDQqR2LMW2Cb6SkkspTHOhPc3N6
Kmjc2RUrMpLEClqEED/zbD5GVGCBD1ZPaFbHlbptwLnPGky+rTbrpcG3jTnE00lvdFLZ6Wx5gnKr
d8F9w0iPb0i66NIAPiXXMzb9aiwTvZxqhjTJ74caMYIbxefnABDvlGEQZlATKHzX/4pMgRbpIMI2
M/SvWxCUzNoPl2+mUxFmg9CbNa7stFd0lNJ9e0FEPV+w/NFAzmqkGJSYJyq59bA2zEbnEHn9nJR5
6VXStjQA3eW+w83rzdXAQs5McAvyx+rQKU3hoqulo9ThaV3n9Uh2OzhOmAeLxGfY95EUF1wBtqya
dD871OCTt1n7mdDcxNMXI0pLe65bkyClIQEijBfqQd+iqJ4eRGcmyI4yDjGe75pVujF7m3deUiah
39UsTgO785PI+6mT7UifyCxBcnwG+d9ug/lT0xFDvzcmYnhstphTNZqxMjIDBRdWfAEADwr7Qz9f
z+8Sv6q9N1keQbD3VbDjFEkuwuWc4UTkPLyUR5KzW/gmUGXWVApglQxaR9B7nZcVLGGvZifDAPRs
UpjgUSf8Sdq+vML3e4DI84WXYQiKIv6I504pSeumlcEm6KWIajGamtCVtZVPlhZaUBDllHY5AGES
hTtD90QOV78GBWoAlI2D6phlqXHT53NK4b0EOy0uzIFZ3/URc2JgJinoZZdmyoCngofGdpe1ora1
i9reF78QSRU4k0umpUvkpBfz7eQRW46I1pv+hJxZ7CG34Zh1gNrDQQdSls/egurG6Jp1eqKv6QWu
Zcor8crKuIDlJNVXUdeBrM8Wd24HxeDnuV2tSuMLUR4tDdUEjaiq2fhmeQwM3/PA8J0423xYtMEI
ior6spFPc48tSh7ZJVvv7wzShrOMImxmFlgALP0xXORi8fPxKhlG9xO2H1Bg0WJSSCCbdy7MzIJc
hTNraZMsb3HEw2BAlmBZyousrAHxscfKJE3TxksBmXjvMArIfqeAk86E2Kwl37r8v1mf5ibY/iC7
Ih8xLiSDBupaMnzy81a/vYGcm8sMLNgHwFYoVxxOfsMfuf6vEyq6Hm2gUIlfr7AUtcb9lCduTtpf
Aj35TOd/hTZsauePrTHK55EF8OnwIjRvw0b7f8GFdwF5mzIr3/x6vf/x/JCtHEmGUTvyr4U/gZBk
6aHTGkyoqo3XtoNYt5G3GlecWnQ5jr1jkSX9Q+bDimbZUBwr8hQV85DsT03/IMPmINc8cO2PVCmN
6RypYNCUbC9cKQ9ICbuwZZMs8gORWmvzIGIwHBQMSGWjQbCzR2ooAKu8HC/wlhHCZLsd2YfRHkqr
XYVyCRDCAeai/4FN1UbSh5Rfbn2+t6c9QW+OBLYPbMEVuwaDwfa8+yzeeatnQWZUnDiGrUvf9izt
hHBIMgP19haFx1ZM7C+IKkd/0188gbOekP9zHBIXdQQihnJVpWmNoH8z3qaGPDiMKPf+nznGgXG0
EtQ8jkwEqKmPFYVJ/2ClCEzHPTdmE6mm3SDZUIER6Ig0eD0vgRncIEvqz4HV84BsyjbkdhKSvplt
V2eJgCjbyYeGu/V6XPujMPW5PsqPwz7Y1LoLy6DPH+Y44desIWQRiduCPGL4hbbb8DuRip1zwgmB
zDvAdWcln09LRtSgEpuG8mVsrRolnp2RHKgMNL8sL8KDpBM4dcBeMReNccdq/odl2IsPTHC7YkAW
Ixwc7gR0ItOQ766w9dDZZggGaDL8tGaMQTw5F9n9wg1FnYmys8ZwjFaAPNmQ1XIjP+S7xLz5oxjE
ld5N685tPLWB4T3WmOaNft4ciQNx01PNs3c0FCMeuZUmkZc3m0MN+FLPRwgQJONHy+vkbLoS6WGB
iVNZHXangWSgeh9hCNinAvf5TzUQZ3IeG+GcYMGqwBey31nCNdVo94loAG9ZfrCzec2zPB1J+ZC3
wFUfGGEz65zuXXIeZc97yqhvlMaBKSKDxQxBZJo9qAeqMONWumnUBpMl1IvflO6P7YWnvhA5pFjJ
WjgQ8hFHk9EmqQi5vG3US+Vlhx3vWvLtB2siU9fcimWWTyu3zKJEoUpq18qYBHdxhXDUYrSAuyaR
P1ll78+hBLjVqr7L6UcGC7pW0EZl55ldSTMOggbgqzbMwTVJRqya4wRUVXDen8WBeM2Z64m4wclV
x/TLQ9VZeyrpDzK61TNiH+KmwKovuW2UbqvG+qYWWpHWcp+cXtDdGUTL+UUcozJjgNdm9gabJPUl
H8xRucj8TXxpeAz+K1Olu8JGjR5ZSFDrbh4bz33PA7X2Sz+dMxCmSksBs5B3K6JNC15DOGj0wfS0
kTU2ZIbHSA3ofyvFYJAs1cfo78l82q9DSG+22TnXrfbP1xMkCaGqhqaLsNdAD/zEMte2n+W8YlSs
iAzpdqX2T/i1cYnsRZ+R/Ut8VwNDTzHQMv2yRzJ+6jAPvo5+obNny9oMNry+yh37Eg/pBQwiEuc5
umNybNMKVjJWSxrHgAa6VhQ1PzzFXix+ziNTTQcQktrvxKNotLBRenpYmTwREbie12pnupJvsHZ1
zsBU0D552MJ9LQCbLsPLAl1c7NbORgd4Wefsej6/B7gS2k0+AHJDJSC3k+9q8ZisJnJfGqkXjLF9
4whCbts3d8URJ8Xr8UcKGPjGXZtlNy2bC7mkkj42UqQFeHNFCLE7ariNXkPzDCc8mb5lbRFJcXVi
OeiB2bxzrQzjDmtLIxaVuONgesTTjfmJ/RG6pJ9018L2U6/R/L01G0OqVyxsFonRqhv0N2+7CbUz
8yCSP3l3/thfkS8o20MIRgpp0fi6lqTcU3DdMvKLjECV1Q8y8tRS+aZPfvI9pneErTLczjsQSiED
kwO/RYoKHyh8pUuNw4DPF7JaoDxh7epb084Slnh4zo0jTOmED6qjjcWuJ99I3USDWY+A9+peImeN
YqhmVpBs/F7vTN8I/FBXGi+ArkMts6Wr9x33EVh3WqDj9DkPSi8sVFAb3yqRKuNyUbEU/bax1zMi
4gMQIBG6h2TCCrdK7ByBv0A/12ac0XiYudjzplDApsKxHpdBl17BSM8hbipeOdG6rZuLbOk4tKAM
lwFCbRaIiqff1XNHa88JXt5VpQZEL4ypW+auyzofhNN7QIhyXgpXxS1yjVdCklIlChgWzrHtizqk
E7fQ6tC3JZsA1AhiJpJuYQh2qAvLCTcFX2z5NsfRcTLZ0UPEukmlR1w6jAGzA6cfga1XbGt8EERP
bEgC6u3Dm/vY7m4vEb1qaBIeIWrN99FgOvgl5AU3GYCYX5pgdWN10TAxHX5olUIyr2sIZSgb33Vy
zkJ4Z2ATXAZjD6FybKr9X5+l5WOsfwe49vKrUVyJtEunRiLjbsqJuytRdWtWv3HNAzQ8/kykqXw7
v/2a7hpZhLdXD0a9MV3LDloMIhzdonwlHz85qnKveR2oPmqLDqxV99ni+QagjjUqrIlO58oQTo+m
ae/7snqo7f+WUplmbu1MEOmsbRjCkLHCj1XT6wjks5qpMDFFAfqWk/skOUD8k3ZlEiP6v6Yjv6zV
kLIKos9nwCuLG1QnXipazG505snYcxZ3IffraHQ2n8O5YyGc1Yn/iGumTU8kSImBQ+GGlzye1are
Xo5TPOXzfMi1nrMWuAlRAmRAExCKhVYubrt5osRhkixqRWXAS/PcKW1c1GYfpQFoujNTwwh2tpUY
PSLWULsYHe6Nd8O4sVLUKFj58Yz9kZw0WqZbd3PY3l/NXp1ZHUJZysMhQ529fOO8MEgRIbqJHhTz
e3O3J/5eWCiy9WNHYQ4jNeZl/aJhhO+N4KCywtj/ND6sfr3CE8qYwID0Vf2GpUYAWn2KxIMJ1XPX
GkR3JH36phWOYo490UUUWr0CNhwLpcHoZBnCtrs8LhPvjmfuUl88b0KMnTy3zRx2f536jFeW2Xfn
u/WrUoYa+yNFBds3+m6SpyQXmFiD9jWdYXGz6usvnDo73nfi66P/7abH1NN/0OmUjDOJ/TBNo4gn
dNelgsWJTXvOZnzmyqn4sZF6zOQhkn9l2OGD2ylRnn64W2kRS6bxwQmRmQWz/hMK2NwFMipGHYIF
XAulpIt0NjIHdfigYdjuH/vOk6Xzdk0aMB+0vXU7QsaD+Iyr3sJmE08hR5Opyv61mDOnW8QcyZYf
2IPKYJ21CnzEZwk5uM1sPJy7SBjCJUBPnMd3VDdodjF/0jV3V5ZScR6fMEZZ+EUWPSV65XDpLwei
Rj3DZnszMMKpgoqQGCiRwrhgppBWpHjll4tr6pz4umMLRM85wHYtG6g8JyALsqhzkBWAzDf8s6Zv
dQuxWeMrqfPlD831GpcTMNac7+Rhyf7/LMN113K3ZY0gVKKH7vQFkXbKBK/HwNx8N8b6gjzdw+ak
eNUiacSsIHweAqKQ86ll38vY1fQdstXGKPc4sxmnGATMWN61b5k5EyY1eEqW5sAIspfFxJ3kTS/X
ksEb+jlSQQuLesn6hc0TSHbdl5b5fhnO7vQ8A4O8Tix4mv9XF5MC7JATfJEz4rzhoyP4sEC3diLa
ELqEjhKsqeXsmUoKov/bYoFa6gWzoCW879CokKxno+jNToCUZVZDTx0gR8DUivBUWn9Xl+k27HT5
+h35C+fdrECwIRNslD0v07YefZ0CtMuUkJeimM/3CJItPsPgODXDwNDcjvniWsSt4kiZUJxgbV+s
FWo8O1i/ZVqCOVSdj/4TtC1XTRbEFbxENBkir1W6w0qJj+Qkxma8sPb4E5XGlmUCmmfupvsbE/S7
3WsVp5XtX0S8VqCNtuGW4IFNXPm68ehpidxaauO1m+YxMKDJ1Pa2uQRWVpZDEYrleZj4MwSAoGZ5
+PZi78gbN8B1KqCSwPijBdaE1z+KAIhoymJgHcoAHmUzfKE103Le1sR/EDk/lYmBotIsApVIprq4
VOgPO+BWkyallPRUwWgiFIQ8NZhqQKu7qjerPLhzgBd54UYico3bU9WGxFnvD8hKmk6VzELakApv
E10scdYkIj6ueaBSdSiu4yPpufAsNvoamdccOlk6iQrLBv9aCYupq/kuxazF6YBWEeunX8KG2E3i
PqP4WEv7Zyg92kCXMaDS5GIEEtNDJuEhnWJnzbwLpcBSKc8X5CSLWntYz0KZmVc9AgaJkmUs01tm
G+1XB0gx9kJotNCoQAZ9m02eEaTxydQ6lIsOYzyVVIKocr9F7OPf1CVmFU7Fr0YibP+H8vlVlysz
SzfDFVpjBfQvlaa/gGXEVx0ImtMPLKhoxQJ5/Mb14vm1g1KEyQcowg2rkqEFYaDVPVCO5YbTAM4v
OyK0eI582jpjP1We7erbGbvdkgbUhKrHEtNnwX5JnGGBSh/9na4sh0y8fuvqPtU6oSFIHsFyu8Gb
e/Z0yXkVjWTby6aFDJ3Rpa5OZvYcMBDypsu1kGao3AGqxahYd3I+tYEq1Ftwb1ERZRgeyYatyIE+
6XCpNatWczI1x+DwREkJIjgCQqH1e3h4Hum4Fsq35JY+TkOymoVVPdknfTrK3T0Oxrm1AHo0rZmG
Thj29Dh0Oh41sLc3MMFW1bLy4i7bvbXMUpZqbaWq5XwAFPlxIWQDqwVhlQUJj2K3mbZpQWEAIKuU
lhz6Pho64Zgr9Smq5R17QorxK5NJEZn88xeSG6uLrpK1kV4fDQjgLBpI/RnDLVNT98DCh0+o6RdS
mQs1wgRoZpehrA6p0+NcRjtX3KT3htNxU+BweMGAWU0KEKvWEO8xbezrmw/NKARVQMEkLgs7fqCv
KLfMEu6UcAtJbkPfwCI8q7Z6M6Uhend60U/umMqCp1mr7XXTY6hXmcuceaCgyCASVKq6j0Wrb3cU
FiMomigXTp1iTvk+bX30TDcGO9Ycm+joNAGBtwhxnbWJofKj3OLqsEI+8DicPdBfb1mSkueS4Fr/
MJaMdvYyIRHkr7U8/Grv7od8w/ZL9rxCsrB7kGl4a7t/sU6cKn8uL5n9jVSnjUsMLCFpH8QjuCBI
28HXbvKhWQd4yBTpns7Iks3J71lPl6sCR5RM+zA7hn6tU/QubOSoiHhXWwiT5ZY2utMl2RfiOgta
XA/2/rQQjfH1kKPdFdp77cHgPw1McV/fYQRcdF2r24bnmzfEffJY3nIeMQr/edzOJrWNZVr+CWak
U//F1E5fBvoWQsaA5hbQHEE0DaAJ8LFbk2Ltyw1/GKOtIo7PXSisWQGRExoQCo6Xb6z0N3bBs4yp
iYEYgrVoYMErfPoOGnGfjTfuvYXLK7molnTQBa2+mGvTNMBpdaBkzvfNBOfp7CDQEbWOpFHOejjm
9XfSXaU+ZjzlSO+cR9aM3HNpisuaIuM7n0iG9p5YSlTSJah6IhIFIDC9cChQrxqT1s/9UUoupnXM
+0jZqLR7lZKIspylDgLvJ5ZzGA/jLbjpOcKxhhaqgnDHk5nP+w19XqnctvzOtFJxO2qTS5a4tBG7
BVtoCzQP8GGeACRGOO9ut0NKId1GyA8bp6azr9AN8imJ8sMKEOeAd1THtN6SRMZEoQq+k9a3iU3v
yEHuyO6/TUJ5Pva3/Y3MgOMbMSO6nEXT3zZCh1MFHCTcRwPVwFwF0ML3CgpkrIFyb54ztiloJWRt
3M5KoORUBNhHm2l9v7zx7baS7T/D9cp7NtdVqNMOTnSTbBQaIS+37by8pkQaJNzs2RIwI8QcGlsC
k/Vk0tyjI4pwv0gy+h1VDMVwovSbLuKRCavd9WdbggVIiFK1ub1f1oTmfnGIXBbf9Pnjpbk4cXio
AX/TRAOfXB4vekerxtW0z5/SO5MmEJzE5Nz8K4zGTP6XF3pilDMsVvlxCZ7KGrge4Rvp+2mg5Zna
EEzV1qL69F8/ZE/+h3acXkr8Jt9fn9cb9/ruRHS+2tbgVV+w3VBngj0qu+Gh+HoOfXb7/VqMuZWU
wF7a1VzBOusK8asH0rw/9qgzU9nQ65hWAZVWaKtrKpQD+pyXY8CFkK2NWq2VTDYGUYFjyGJiVGjn
OsgyhU0k+3vrjptaczO1e82v66o6WtrleL/jYJItEGiSlWTCTBtA1LbirXz2VrmcEX2/fx2PPWMI
rgoujOXo1RgukaOg+7u9c1nhRr3XUb6Q3YiWrSzeljcLCHOCrnsMEUiWZCps7PBw0CqvY1sJImSC
F801KzAu5uf84i5F+LWQXbwiwxcMzvfEXQeSnAvS5j3rC0cNk8+onInk05wYqV7PFbpep1t/cLYM
Y/jwTBXOA4Xy3tQPY1g1hBDUBwub4FOSLGYZofJqi4lt9qDX04FQs7tfutUmix+7AG8AU43Jn+bw
kRSONnWvOz9aHkDWChHPd8h3FR5eghLUCde/MAATjLV3+DLurvbKQke7iqBUG1gYa2kguPfDsNd8
2fvMIuM3TXwNproj5smbK9zK/fKpIUK/oX6/TSfjFDk44fJyuYT/geqe0TlP6C8vWaxcCusuD91T
OXvYklv9Th6HaQT0nGGBvzAG6Iv5gyRAYh7NDU7bWGJ33NfUOerM2euzUtt/DaihvA8Zt1RDtU6n
l+ACgtohRjF1dxXrccBKSpNtqBisbVl2vEtsYnlfvIc/Xubd5zNXVt+d5wI/bCMCXPh6ziovf5tN
UiS4tIW9u7AftmfBv2sRIk8QZySj+GvlRxotMqcZYTppYZrDC0AC7etm6FiGvZuQWa4VjlGcYwnA
HNEO4xCm2OakLYFyG2t7fC9UMF/U1L71Jnun5EX6A2+gIqRs46ZM2ku3xZJ6y73KpzKOayRZ3HOq
ZvO+9wf6aERSZiRClDDdsz8WxKqthgQbT9Wj8bHjVNnTsRHC4CiIftOtw/kwEHOS8kzxnoXLB1AO
7weEnakHCV8SRk7MfZmfdG+Nc6wZ5DXgAL9dKrnhsJdcolFUEWhFhi2gcgXDMe6o71edC9AfwoiZ
AMCvXz75+VHcE2I56TUXPdR3WeO509RVj0CBThgvAGQZYviZKQZcnN4MGjxcDUbMVEg87/Y3QQvI
dJ1A4NCqZTbGFj204GSDjx50biOp906ICQg3nzDFA0MbogPDnYRQ1+uWUdNGzDO3YTDn3ZqEi226
C/+q69QJi2zFMlamJZKeDtUup5ZwUKNy2gmx6Z9QP+C8KciFhbT6nEccAqTZvglunbgyHsDuNjnH
z6hfqy1Ct6rzSa4p7/Z+eisfsFYR+7IH8I/xy8i3CqgWF+awOkqaMmCnXEvd9GAdWHuLopE95690
SFK5Zl659pd2bxBIHJwrj+jH9No/3S4PcrfB2hwTfYGN4YWjrvnEUsuz0pYZQcYSuPNYZbRjmMmC
wnpA2MXwYIkSz5FO/guJD1WM9wgZI1XLIRzNB7QB56Rtn7msaPABfXPvaAFwWcGFa7ZtxjLDYfmO
sJhwOg+lAcFux1v9NjDQxu31P1F9q/uzbCle7WE9s1puDR23Ysi1YA1YJSr5tucb00gwS5chRZFd
GCAR5hHwqZZDsxvoq/2vhd1gDfT7p252PtLUIt9H8LY9OIZrj+S27ZHl2wDd95FskCBScR+eqH+r
ufo7qCHDzxTIFaTeYD4laZcRJOx6I/Hsx5JU7PvBTqsbgzd8QORqCPflW/hemG+jnHZDxRld6bhH
H5hRN7X9uP4XLOOkoeLaBHA27T0b5h8FIPGz4Hzqy9ZPsI/s99I8CkUbRQ4Khcp2sMvJw3cHFmJv
+FhdanE2OdZyxm7nsUbdmS00DxME4X+IVTYFcsPwm4hMd6tqInuflfztG4zC1dvpfnLLhg9Fq7NI
Ik71YIZxOH4aWqjUP4Rfgb+MG32tY8Jw0dekm7Z0kgXNO5Izqdx0UHXgEi9a6WyIqnd02fwWpGgW
ijnZG4Bmj59KGIO/Gii3NrzB42G2LmoMteBy+74mXwqGsajAGnwRdQQnNZYqCEM+TrPXG8Ao+lRf
69iiZCAaKFdrOTVQS1B3sTjxk4fZU4ZKuJktq6b28kU3la5h5Ra+u9KzpI3TK1yRFC13m3BbL0PN
pCm+TFQ20mkF1syhPHiwZ+Utkhhw8kBSt7W74KhR7BO5ZU4YP1OAPyiHY4IW93Ot6o8ItnEAmNdH
NkDMDx1+TnMyAdlnsUOqq1+6U+XijjR6f3c/10Umn9PsNsYK/zgvHbbdFop8Ynyo/EUFeaCk1mcc
gQoDrRQIQyh5FM3b3tmdcfAMNOYk5vrsrQUVGzNvpzIaUR5rTzWaRLh3lGPqaPBzaHEH331vQHyx
Oak6LB+XQ1CCvntZB4KXB4U7E64gR2PkBBtHV0/mCIWGWEThZ8AzmNdhNwFSa7hTrVEau4Hlfnrm
8XtdGlwHKLNJuNITvAxUp0az4KdvrkO3hvQslWqPN7oakXB9HitQZNQQajwXx0CiyI0czCA9eVRx
3Rn6tZNXy/ssV2CytfPZjn1Id3YuCGz3+iCJf0YiJhIHPDROGUKdT1CaXaiUguhd8+DaP/g2NO+4
qgoGgwKH6GDfgkdz0OQROi1t38L+Za28hI4AkFILGZM/qbAW4HLS+4zH1+ZCGeUOLl9wPb8EKEJj
i7PQxEVeUReWLg7Jr4kvOkXTZ22Fn++PVU9NDCaNTx7En6f/y36A7M5a0UoiIR5NvN5PS+YCdqf7
GYPm1fya/s9R3Z31ACpwIayGykbL0m+F3czZBIc+PGD08xarsPHZRQdE28XwuA3ducxjq0r16LR7
SQYiklxfFZ6THhW1cBvetR3RSErHzyHG7aNT6Nyk4z2vEjn2qLrAIsSdfNsZIf9ZalNjI0gOXbkq
TyCrUA02JabIxW71EDHoIDEyV8tt7OY3p8BQLiCgZHsQ1QBOzgb+AgPggYK8h3Sf4ARooVVD5yfz
dax70ZMew0q0Qeu7taTmoHowuCfvgZlTSodcIuuuHzjiPOeG4f+8OycJ9cgTPx8upCqEKsY56yYx
Ta0H9B81Ve9PXZ8yU/kwo4XjHSmIYFYpLLvdpm77YVYBk8aTvKhfVvv84NgWwMCyxZvWjHcZz9HD
417SadSARBBy5N+RQssd0B4+OxYRL+fkeLaNPe9Y95qJohvsX8JT5I2a6Y/oH/rdjvCZAsi+QAXa
ytRVMIagR0rTsOTfyWCJjy9VtGcrANKgXh2yIRbaWFtftdiUknKiFy+Dv5yq8YKaslqrepKsLR9g
PhRAXJzPHfoFX1V0ZUt++u/lGEzyLtnLV7mdEXt+T9GNc4wZZnV9Rj/f9iZZJqpEfsTQP0lzgmYn
wsFgbsiVpD6TPV2pN+jNyzhDuuS5pcxxaVjNuTimOYgaLDwYMEnI6iWIHFpj8Pc+k5FEC5WHbqPw
dYz3XJw4CSLBaMyoHUtacPbwdFNNUWipfqUgJMOPfGGSXiWs8iHWppm19WWKPIcaRrMQx0SA4kQy
0MFf+c0GTVQpQAfntgrKQun7GceDTm6Kv/8ndNlb6lJmB9dmb/EOwVjGqZfJbwVdTfI59wp+hjgb
ASmrBamIBpv4xHRscztL3CXSf0oiDSk0qf4FqwswzMA0hb4NCBZd+L0tDBk6u9lU0ukkQNy63iHv
dsafl3LFmcBHuPmLbyZDmPqOPmwT92OacmEJIQzDf+elbYH3vzmai/lcMnJfVrIa5OVQXM32Ib77
zO1DD7dj3GynV/NEknGr/Et5nTt24opZOUNyESNVtBhQ07+KnR0wALMh6ueIY4HpcO9rE3aIO8BJ
9toJ92h8prw9QOBCEqp3gqFeXuzkjvcTpAlptTcqtprSw96k3MD9HBK8Nupv0DWzIr7JOMtxaBMN
kFMoXlF60iXBsrBdzAg73gdlCe1jPK+2KWyy1HENcG2AdsQNUq05I8Gsw65uLwSjS/xGHh7Umk3j
QcMXpnYTfxzElTCPv482mj3J5KuCz0pkZVLzY6XvmPlpm2owowKS0Zegz2FxrC9dRcPBMpzSUOpi
El1vEexBMmAlbrh2HJOPQnBOvyuA5H3peV2uc7EzZX1oCIoFi/UZGL0PIrwhEVYM/OOfYGQ94x6T
BE6X/ZrUObfJV+3E5yC/9Dt71QCXZCL9klUSIU2wwuA5JlkMLJgz9qiNdIR5ADsJ015zPu2nl/XY
5SB/LYtcxiN6EOFMxYPR4Tfq+mKLlqiikbk/lHJC1U+BTonyRvQLZ/9c0T+dGG0IWEvApMbGvzEw
V8K/0tYUbB9pJJCBsCylhOaO6oZpujcq5k/yHzWqjIgwlZmn8koFgAI9R9EgbgUBcZZCkcqHTy3g
sl5/+JQgfkoh58UYoGjp+ckCzIhwoAm9WqaJUxwV5ylROhwiEmLvC9KP8W6NUpj8uAzJ7bu6mMoA
h1Qb6b4utPk134/5Fz2JrFE8Fnqbigsk5HQpood+2iilEpq0EZujsepbR0iULrzzNyWJdA4rebwz
q/AUr0jhnbod9J1xQL3OjrRKXMadvCsu46Fc/WOMPgZsTbGYiGYP80WsOuRY3tfyhhkFDIpdr8Rr
K+9piUnG4luCcGRfOdLEQdkO85lcc9PYK4pjsILABTUw/TfD6TTKxOlX+W8zjpj7hhLDwT0cIKux
jec4gs01HP+JsDOaj/LcvQJnuY48dXTLpLlTBxsMCdq3qb9lsyLc1pO4Dt52aPZ3Q5sO5rSrLELK
6zKYlsws3sQqITzk1PcVWuOQYMqesl3c3yHgGpv/azAPMbxpeFCxzfn4JeVi42f8a1Gg5uBCIsgO
CH/scKDUeFDV2m8guC0n+bkHwV5FNkBEJJCJAhTTK8RR5O6eXqdWcSiZWK4b+1QxjHLYEDjZOHNb
lgUPE1ERw9PmdF9jgUdQD2tQo/uRJFnlvFJufknSmxT5rcqHZ+xGONl8zrvi1xRaOj98hyf/YF7b
KNZnIg+2fzDYZKEmaZwmecvQdH4S23l31mpV5j6epBh7+lWfRzRVKj2Mpo6j9i36pvsSfTeoog2u
IISB5c5PiIN9GxjXIdjUSvpmGYCqolU1IiDzaxQR6xWPGVOrXRCTp6B7bdpRKcNG5g0P0qcktk+5
4Mtmvge60AgyiN6mSMpxgVv3NwDxliBeUv6vk1Ll/H2UPnPKnlSUAch7lAJaRNE3z3Xc95CqThac
DpPlJ5C9fDiWAZPPMLYSv3cH5vAPGtu3CRPMJedfWjxpQyuiQ2YgcxZuBWFefQ+tTnEwo7f4RfK/
o0HYcfofZ1hLI0D90ml5J9tqIcwsfoB0td5iW7l4zbL0kbuzUquyZnJgNXJqJaCuinr7kzTTKsIS
/YFIaQ9QQ15RAy/KkLepoibzYTXqUmeA44PQtPEliftM+HD9oFSlv9W0rnClrurbKAr0/ra/XMmU
+dIG5mXTJMqUQIsbaajdeaYYL4o2QiqjYWEdV42zh1rOoCGxE/sdOq89N3FwZdw9QCsRfjhuDX7x
aBwUNn5mery9z30OU2RHsQHdUuVmy4w896cisXgMMDXA9JVPNZoBwWxqsSDF9nslxMMQriG95DSI
tHRbWP79CfLLfmPvZUZynHxt09WLjj6/av35AvjQlOQ6//zLjpjQp2CfBK1uhnXppDPbmXdvDNMY
uQsiCWq4w/mKXRMUXar6kR9HVuFOA5/Si/zj+PG9/RMnSjjX3ILPS+s0kQHY0nXF9Vt4vRsSeTgb
01owGfJNkqoApBXVmCBGvURzQlYJfeKV5SmAl5tWYSpulwn7PYSRWOU1hhmCZ88CVkfwXmWF+eD8
VCV+JI+hYOlvwZ2YUEhOMdzYzJTiIKdTD56ILvFe2oZQchSiNy372X1Jg4xACQI6t2ZcA+6ZMV/s
s5ww7jk0VmTfDBp6ZULTHrit5DSnNUpxT1Jiapyh9/2G+OnmNvFGByLnoHr5/PGNIsAS2+2px27i
nv+zmdFAirfqSD73GEKLtq6e+aDsARW+kzGdJ2euqcjwzXRR6VH2yZfNUTlRNciZ8X7dPj3Xc7Yi
+5UzwRysagZmrZQM+Z4igEbF6yy10WVk/ZD1QiLTS2AlX0f/o1PM8yu/ZBaP5bkMjwmXJAmuGRru
2GEcQzt1y+YiMKPbVZhw+Pxoma7ay9L0FYpBK6DXgXOJs3Tq7cRz3yoZWBsBiG+V975aMwlG4eKg
lfxRSQnwcLtELpyMCDTButrSRlh9HjEUuDioznNZVI6TgPnTsLa8DKf8TJdRdj6Om1Mrdjaw7JDg
tIi/Mi1twrcePAZXuSUee2arP2QI4peVLvYx2Du2LkKq5c7pPXgTEEag7odV8R4ezZoGA0OERBak
/nV6kDg3Izwtt/bVBsu4dRAotBSzgj2IplHhyxq3BV5m98b+hcM17r2uLr19ryveM6i1e0rp6WWy
Mt0I6Orjy8jms+E5flYlwagkf/leyZ9vxn/+b6GWcp185I3nlk7lj6Vg8JGWP7JkGf+222KFdyGA
LDT3msJiX5mA3xqtSVWoM5+nC0KtGenvGXf8kaHi6d5wLjiv81vKrAg9ZyCIuwK+QNs02A2iMLiG
/Klx+iMzaXgK0B9OCphMtfgepep3agD0CEProtcWjT3Y+crgPtX6YBHfrl8apjW90s6G9pNNALw9
38rZW7R2Ta84kOf1QmuOWDHdnYTes0IsW2afFqEH/4ZolxexTEF0UGLYIwz3knbs0wWwTR3EosIJ
zHOehNTFfSNKYDG9jWtEtsXLByGAjUkGZLi3cv9NB3Z9qXZjLWPJWKkaR464YKIK97N9n8CRGUr/
BCGFEb+no8ISne0e8rMKzOlYnAC630UwvAC0ElVYhMf+dZqDjNVXnJV8NFg9XBpoDH9JE+D554nH
ffg4Ly+2S4viulGgxtN9f+5qGjGgdoZVsIUzBEaJF7rGc/8okVJtpnDpFynHfPpezb/Y9wv75903
ugbKEY6EE4CXSmOtpxIrrEQdcJtW3TOGSC55Lk0uyQTlEmAIH8+CkM5kyDJ3A7w97vbq/BSYFol5
4j1MTBRA2lobXatmh7wpjiCfXTyP/YGEYAaq3KGxXGQTvr3uZYE57ccJz0z/Gcxw4zaJarKo5Pvk
WN3iQO9KmveyPOnB0sgCS1gktA3cYcVHRBXvHJoc7XGmmdr6qadjCu0oiIIhh/MjgnmG14JlM2/W
6naIgtejFABe+A47gphQb1aY6Bnpxo2kysXNupwFTGN/DnCX9B0AlBig9uf4kanNZBHSClJlVpM2
lfq7J5I6PcxnNua7jMq8pBQ2jE5Abn4ORZ5Stt5L1/lfE5MEfWLbRQN0hGUtz2cwPe7o/SU6pFHR
xKhSdLk5ZH+mK1IvWjYUG/B7nt/B/8smSVYkzaYctofO4Hdkfsi8iiadp9qVzn9MYBSrQMfYP2SJ
T/1kYzWTRL/tS9LfNuwtmgA8k94AfvXHtleDCPq+aYRxWt5LmYYk6sSe3JaOstsv4Z1WrSqZCWpZ
pjR1PeIk9m7lYvqaQScVrX3gTlfyz9VwRa8uUla8JCgO8c/XZtv0XxMfJklj8zfgQc7r2Q4CBWmM
MD1bRHnFyQNqqwRn6yv+o3b306hg4jEBxhVSSTim2BFVFCFvu/ng8WRF2eXpXyUZftX7VNK0aptR
CqnegcJk8QT/spLUDAo2qA6p+NXpWcB/wZbj56YBRtKWs8YyeVTrqPEuEDbamMIOpwMABYTevfIW
lNAxXR69b15vdzruzw7lTD42rXUcWooqpovgxp8e1P4UGgG4H2m+bQEUrRGkeW1bXRB/+RvgMeCJ
6frckynFuM5gIaaOKBq3b72L+ZLiN5Xj4s5pAKdsOu2q0Q0eRYgR5JaPA0WwhW8IAyXYr72FBmEU
8DS4RORQlUDc9y0P4+yT6QxNhRfwRDG6hAUsppFZi0X/ZY2zZYINwRfrm+OY8FBugU1UZ4gI9jwd
Qbxd/DE7i5lwM6sEXwjA+9ch1wCf+2b3/sEX8NP5YVSDFknqguGnebERNzh9qbTiEHhAbdcp1udh
jV8Pl6m3eyiDot+xfrrs1TiWJFzHhHMEOyg3Ekwuc79+juGQy/TR8Yj5Z/zpnY9DncrlQNbbyi59
HJzjgmwmHd0Br29G2zgtlGWdJwcoPax9pHFX+uyIPbdCR46gZj4pUbTcHWYvbydNSiL6saKnmJoz
Hvk7Ja3nZ4BkjJiLnowqSm/Nud70JIqVtZL8WX0+2VZ8d4Oe93HQGZMYqCNbYg15mVfPakAkUCes
frqnWXMibv0iOEoWmi+lmHnWs5ld/lyUrrKVeQ9bT23Z3inTvyCW7C7ILOVkxH/xS3NGJUKm9uYg
V3OjrXS3zjtfjqTELE4b56mgfpUmWgSIrj3+1z7HkwyhB6iAWvmAeJcFI5FM+l+hVZ77rEFI5Rj3
04+mrQBnyH8gzyv5pO4oUgehYCM3O8Ra8U+r9qrAJ2nuLFzGX61t+k3GVJS4IRVJQpEQq091u66p
HHrvG6RTVKVfSo5aOm2CHjx5cMSnM0JX3Mdu95oz3OZNAqC2HZNBMlThHfyNv1HRQhRLZEekf5XX
vc9WIxcEielt7qmXZm5im7AjaTVZ6Egd/tPnT58LPsHceCvizpJ87unrGXUEf3Gb7rWi6LXqIhlU
zq5PxR/oDKmRRU/my/r29LkcXQuZpiB5+nz8q1teO8ww70vFMKoWlkUnkDtFj0R0Hhc+PNaMYqta
AvMr/NEojLC+QNPubSD8GtKootLIZHpdSNBwrLlaq6sooqVohK05swyhDLhZ5MvY9vp58AKSVrkB
4Y3ntO0QG8pgXwnnFacarqWjK2tn4Xa4Yl6O4xFPLdV5v26rFq//SZMeAfLEOxbXmOaBwB1EUgXh
54uN9qm1E5t5jxiHQs/zvG5rvSXofWk2Ju3zFfzvT/tjqkOeSg4LmjE5C2PqzOTjdWgk41fNkkj3
76bkuUMqHmz847MCDgpT7zJmUVLT80cZaH8nM7HKhquTouMP09AdWtphwjNZdLtZA3vVpkn5r0QC
KsgK7atJ1zZXUUPT5LmSl/laPsN4V80wfuAvHQ8KdlgmEv85+eVwn6AP/hwme9J0pYBwAye0/UIH
dIYxZaKfqp45RcyRRGGPt0Ru2nECPbSed7FQkdX6wSQehBnDloc/Gb/Ml/wazP5SBU+XQ14YGLKz
yl4PxyxYNrLFy/B1azaeMgSSxS2o8N6y0C8kxocJqOL0hpkAyTZIMmgbf4ti/HxYUhL5SwZ7iSNH
AMkgyeHDsi6LeL3WK1llhvQ0RJGqcCLC+nepxYN+rcCxjLYfhv0U7rPB7h1HNA3r3QbyyOrvivJF
uEj4hB0WdcunRx8VpBkS2qzszlSup0Pkg6H4z1NTk0lAUmkD99pkr27t9rHtF7a2g3Puk2r2Yxqf
ZurGZYCUjeEXQso5c9ON30/htwOfGwCBfIErF6r15nJ1rw68/9hwVWSfYy+36sjUc0laM644Bu8R
x+0thJv2+P6BmbzA+nhMiDOx/HISXZj13j503ulRv8ykzjCCLjbWWPbE/eupqIMaNNJojEZOVM4R
RUp8WVhAS9zNyol1tmWeLxCxpzKWcOjG5GSC7uTvHwxH5vN1Z1lgnQXzMvJpXUcZKFip4I6euEYd
/xsI3wyCAfiXRQ0ppdXKow5EqkyomaAkpDY6K4//I86kD5I+5JrjgIRO6mz5f2GMqP04UlQybSlw
9iaDfBNygdLkYkudCrFMhB5Og4AL75HPRM5ABwIIfPnWlFGeTQwvF1q6pZQ98Q6ZEjtldm+cPL8v
8cwzpnChnRb0asCo8No39Y3G52+owFZiff2qI7MG7Gt37GLtFYhGsPKG23QoDr7lzXl4IlVHuCDA
Z6bMxXLfi4/UqA6s+tyXCFKk7hxPGWbwH4uQK2XitcdwiFjyZnd8+C1gR3LoUmn/GBeNcB3/M1Gf
YOOKWA0bM0xhj67Gprz4+ksvkQvfI6zfe+teR4y4KmrelQUF/NzrUOeoKc1ChRG6sHiEZBm0z8hc
hRjGrWliiHrlwAM4qRi9R3q29kKo/qolb4oDYe+7RzyN443/XFPjwz09Wz31UiLoREwajs/mAMNm
O+qAAa2ErJod7jmRrJLDq9MKgfIctr4qRFtDpIBBUb6leTpYpbRwxrOeU0Ov6YPTGAp83ilPu9Ls
qSq/G62emLypt9KpsRhVR7tDymTQ7t1lHr94bKQfbE1SFelYEiiRJMnQ8oNr2wx7VmGT5q+Y0V1H
vYMDo6I2LbSJKdCHqDjihMP8V6HDIzUcREQvzAsoHwrcoob8DAJXDuuhNBbceSsZ/+pZ2rMfRf/L
WG2mjr+QG4gkWHLx1oR8tksD7v06vSyXJ2mAgLQKKI7zD/nJB9zsNRecB0uLW2bJMOlfAhp3tYKZ
2keWPdp1FlLJPJ/Qu+Y1ft115USrNUI7FlFUjIlYlwiCQGqx8zA7DI/d2rs/q4SjrD8Vcxz6qPuG
neRLV7kPRx1i0kc0JJ2GaeiKkjT4UGC7jAyA08wDNPD1HjlN3Q+Gv/WhtN5ypHN2qMGu0UjrqknB
1NZEZ9YJKJ5aoZqzlAxvxxDUYVOeTbj8bUmZ2hW34h2v1oA1/Yc3SVDBnktqan5tytBwbBbTWUbk
UFsxtVFAw2dVoKNvzZJXWNb3RQsSgRPPHHm+0bfKfkHx8l38E8fZkHu8AiNrul2lUMH3iscBdNsH
q8P32lqUYxaqva/dKgZnGqvrGTtoNL27dUfqZX9TKDGtZKSRU0GyVDFSoXA//I/gqwAUJYojsNdF
36oFzF78US0V2I0as+PQKzU3KV8x5wFoYleU19Z+2IfQHSZJYND4Fv8M5aNwkes0UUctiTXW5WBG
PYKJ07neT2LU0R2zCQk+voYTUcHskwynU77pRiNd36mIC0X60j0hQGPx/LgJMpCJSmhZoNSl59kO
E/vtYH05q8LJaSwxHKHFVv22LUSTkTLGx5HyqqXc25Pol70v0gQeP1nr2DYXJodafLeT+j4W1/AZ
UptWEcAIf+THowlKGY/yrcxMfYHC1u7s4vgt5o5ax+46YWWLuky6wKoY3+mlh0DbLdOxrglMmhdy
HDkpTOguZ+DZejq+RzDsTrsHvfq8jBSq6gEZsK6ydmOOKcQhdAGF2YGA+RAEekDclxX6+3N3VfSc
+Ycttr8SNCgtWUBcOntaw2kg594+1GAgOfUVGcUPf4Fy58tpZA0tyItQCQUVnh6jyze0tBSTYc4h
ybY/KZxq1R1gZpaaDA0Ik6MK5Vt2KmF3wg+crXPnW54p5xrdObx8Y7XbP8M618cRfQP8XSzIbhIJ
KUjo5hneiyfbntIRGgC6AhfHhAWeLfCGABjdtEwFq2eLMgs/nfjhndfwqhnlKSGGFqkwsVdALD8+
WokS/FDo8k71E8xk9BsE4ItQPnWNnwZh3ufKxGQoEHZ4o4GMGuLGPV9txdqcFOri1ii5fhsZfEJb
mNpbVmnsOKglHtuiGJdM5aryCG5kLES239xnRmM0+DZZAeTd5dhJn6Hss45TKv/ax3qEgmg6nLcR
N0D3LiArM68lfjzcKHX9OVLzW1QRsah8gGmjpsmz4MOexTzUbeaHwo7CVDmzUan+Nt6e8VhxBWQr
775dqP9i4+Cl3DSbkmCZeoRvn5nhVCEOsRC0XYfzHm1S+4AaTfqHlsKrfAfN6lnZCCpJwPOsEj65
5JfFLxHb14vSro3vF2cE9JLpp4dAXAD0vsggR6ARHhdRSd1WDjHJUGfH/iZd5/m2Ib2vKQ25tHNT
EBCBZ90LtM0LDwkNlFX/s1mS/tgYx0G4NvvQXrAJvMAeAsSsyRCjfCxTrA9zjGvCUmWXMq0mgDjk
i41RazvB2TfypDLtr1Br8Cijo40xWMz/KhGOJIQfxzYVXBIkciDAJoA+xeTVJ2b4vtCw1befapfC
iVAzSxGRKBkNUKNggmd09pxtQ4jdzsUmq1jFRIG1V28MS1CBz3zAKY+x1+yDLajcZAdWqyURCB6M
I9z/WAPcEkdS/2J5CbCnZPrPnpOWnEMAnwKS6jfyEuqLyvkUNPsaHuJN49CN7qGQ6xMFrUW/Q7gK
gtAln2jG9gtWZGt5Fqqj4Rk7uttqIZI63kNL57ctXKa/erbzKgR2hEYw3DFcsJRvFkOTMUCJdD7d
jj3uILO0ETisqYYt3ulTBOKjJgFpFXYnmX9Alc72/KRWDt41BFb/trEY2UhSo7LlPloCBfrFMpj6
zHyiJerbhpA5w9VrkcknFtaWRKhtw9mBWqophz7Q2AGTfQeokA9HocDiz37Hx6Wdc/Q33DXBOaDq
gpd/u7HTrCdkOqZi9HLd2Ji2a2UxsPYe0I4fyhh7/X+sXLHi6+EfNDk7NhyEaA3A3sKaPJLHEaNq
d1F26anltdiPLGOZv5mVqTtOsZa5WOzZzfKZCBOcT4dfCu+eEQxFCP/+fdRoI0KMAGLCc+LEoSHM
BLsRl85DwPacyCWVscYIMsTDCoEN0nEVcLitsFyKapUw4d4cMUqVhqgMHlk+O4C8Hk6AJfJVoQni
xxLxc1VXfCQbiELuxkprwp72ytcCyQyfCdrFmCng9g82UXu/prE5IOVjkh3JVs9wO/39XYn+eDMO
xfoeHz3A6K6YsGp1UBPNwwLK/K3AwDtq3xWWc1Y7/QZtHcJuU9oylAkJ/4j1jiv58KUQA/j/A6Xh
k+kiBSZz10F8JaKMYgPZnxrkIGjJMiQCF6Iyx0AvwHfX8Tj6Uiy5DW+vntY2r9KDYm1GGGUTW/p3
dM2Cp92xJWhD0LqzccG6CArt3cfI9tDcM3q2SRSbPNEx6qw6ikMPf9G1Hs7jdobNn7LDXUty5tps
+OqFX1NHkZETR8gjHOy5R2WHAZbi7zyHCmUn3CGcWi7fXuv9ABrVIR3ZTZGPdzBEuxaDVek5xKe1
JNftonPZ8KQSXfRnwbVZo+noGa7n6+mP9FoZW6vpsc1ivC0JBmhoR3ANGsqWBBqf2Y3hkzE644OR
dd16pFVNrXhWD5W8NCnHsunb1M2CurUt6TDreDF5XcaYLVjcbnB+D4lVWvBAkktTYXZMKbTbpk+/
EdY3QK0YfMIjFLxWsn0igEEBjyHvK5SkN0h2vd5lgLVqj1f5JxI5BKwWy4X7DXmFbelu0LzfWQ6V
kLbB21vOqw4NuDUgYreUs8hLKN62VpZcW0yIG4kZk3ESnXAIC8DHXjW4tvWKym4v/w4zGlqAG3y3
A2tKixbZ1XX1IulZH7d81OGFgGp5uC9p2Goh2lDdi6vTI75VGmrfTXSnZKqv06oyRRrTlSUZPN+B
sqzWHeTILq4tQng+O9mhk41S2VnODYS/yY7PsVZAMx6b+aQKxGASjFulu1PNL3F3SLE71ZnIszuv
xiMOGOYbQX53/ZTxTl+oeZcaHFKZyzJJADEECK2h1wFmX2oeMcOKMo/hADyKdJbmTWBVW8xzOpp1
qizG/qkRuVAv3a+jYtmjQJa3PFxdUGdXfuUzqVqNC7xNI/s02x7bupenZ7fO/olk8XD0urF//xXm
r5OWw8O8muQhhqIgsoMkv026mtPYxbhCMSWuyIx/sQO20iHjdevnWePEVfaFq6Ll6zWHsbX0iltm
pBSP2uAuMHSyX8O7NCN7nLBD0XwtI1Mdz96I2395Hysdhb36CkOlZRxk2vBpKYMx1uVPFNrhzGvt
oONDI2SIi3NjjoVzhqsr+LF3mTIVfFiNFQ/P/M3WZpeoMRyUEzAWICz+WDluH/47MKEYQQo/dsMt
ZvoKujTY8QwV39ObrK4/+i2W7CefWxXytSkDm3QqpLD92mBDmZgg2OjmfLZwhnBBIlPLq08zDJPV
lDrl9AfgeGN5B4EIbFSSg8pH84L8h5Dp3W8QEdbIZ2oykgzMZETOMuYSr4FyTR/RWLlyeAoxPVtA
I5UXG80YfZGv79rYp9odw+eCQxrY1TKVcI6HfLHS9LpZuDAwx49g2zt7p69a+Vp2mcAW+dXkEe5H
G5WSOIjKOKFrAh+igkBlTWkofbl1/D5lySd8SsREGSpig3dYNjDwQNsg64MsYOw1ZeiTMdElH92k
oV/m5sdHwOAoDSQTQFztzySPqmB3zzrs6+8GmLaMwpuVtP2WjOjD8ERye59A+idEKVCNClPfvSaS
L59QKnXD0ZSWYSh2buf5kxgBUV+5agakLBLm0dvD/h2OpHJFREMtcpHKyxOcAc09KmLaKtWavpOv
TkqK6LOXn3p8MR6nOsAYneTrytRPkXEaLS1MM3I3kQiscEUrntxqzHWLyELPvqxyTCX8bV7tyIvK
oNQgw9JlAC55w2lllbAcTWD/3ZNIVTAcWrued+OAd8TBq9m5tFG3Ens0f2Rn2Oz45xwYgC39vE4j
VtvZ6Ihq1x4sz70b73JD8MGItMEzbN7rbHs0AhFXPvGc3iXdtrA5mx5vNJ2nZJEBPjid7Iqxm9Gw
U8qHZiyKP6IO9huIjbjB6pYg3WVrx9Gg/GBkMNoVLx/eXfwsdP8HiFZswHWFuMaq/ksYPI885HTM
irCNSy2PopLHuIMN8zB6UWwd4XLJzPyVeaLCj5Je6HGWZSV6q+RzvGQdUVh9pIMSKYIAF/acuPKj
Pxh92fTRLcLUBU2LUneuqDHlzxAS3ZfOQ0YoqmWpBNnAIQ8KyraElZdbUAqp0De30dK8dmHI7+tr
rZY3uZkhTd2U6KhNvS1wOKE1TL+Fe/FyU4Vfj5LGDDBp8GzR7NtRrzeIr48qcweSsN0IlZvRHS5K
YuP6EidbQqcSG2xxmVWixqhHK/3mIVn5uEj7IrPnvfJQGszdgAMrzCeWCgGon9/BZQKa0jkojx8o
6iKS9e7IC6oIskvX+BEiGW5pva+tyDcW8OQvmY1cvLE/fsX2y49KDx/mkWHc7v9RC4uHoH5YSA+R
reWDRki+8PIVI+PTC+CTlgZVhxuYYKpjbMWgu+R0GSuTWj6C7eRYSD9eKgchE3kp/1AXdzii1AHp
xMx9OqpgWubD3RZIaE9xEts3eRwPTZ2huqJjRQHpytPmhBt3SU9DMfewoheCSY9RNJd2kLWAL8+v
m/+TnhQcLIHymP50UYtNPiUw/lnYht/OchY1GvOYerc9ovAQbCnnJBv3qW5XXqU2OZxcKUie5eSs
WTf7mZpdknb9Ok6L58xmkXO1edeLtiyX+omCSPCrRwn6UkeXbUPbVz1orSMe8Qu3cMc0w5PhxCcI
zYXHZ+Mn4SPl0yFF4f277MkqwB/FYiqVMDqYXFK2EgBMD4EesFvi2IJLhJqw+Ar4q36t5yYXmIRr
g9A+hO40t2tQ6v3Gzj+I8SEFQc62b+mjbN7zExtuYhsf/0RtnJ5WnfFCA9m40HbI3DFX91Ns7Tlu
Hodhz9fIs7VXPoPTsdYrgk/KLXXF1jFIjeU3wbbMkzEMg2vBv1Csx/086oKBLcKm3cdJW8Xl9s2o
P4KO6sRPNm0p8/YF4cxqVixDni9b1YdznkDfuZlVl6Dv1x2vEPkP1JEcPFVd1HKe8TiV+8NcMsAB
v+i5xQGImx59Ajkvswwb2uH1TNn1DWClG1jhcSMuPMfql6p+drxE5wTWVvqDN6OKili6/PZGGAbl
reOCjPjfiq8XHwnGeJXh29WaLgs6hFV+lEzhec1vqoC0SimSPFwloJHJftQ9SprOvjvyiHug79jx
fzIxIFtIuIu3GBW9uoDtfuQ87kXxhZGRDbrxjEh+o++LbSV9P4v+UsFFvmvoKjO/stFvWcfBYhPL
cQnCgy74gf91hxQD3yXoAfq8evYVJkehVq3SJYV4FG02ajSYcgmV9ckxGNt/BuVF1iUEk6/uqQRj
/1YWPR6VEFrWNNb8MElEF59WYZ12ft0VMWC0ihI/b7gg7NtAGHei6aA1g5WnK1Quq8sI3UVEfGng
0eTWnt9+YdA6ntaRcxH8OIG1+hQRzLyYsfymvXEctSU3q2kqxgcWtQvKdKD6lFI4XhP3p3V3diBJ
oruEhhMTNmCyLbyEOyOvBbhfCVFI/qe+WzSHxK7aaZIEYaMwuLrKGKgNCQqPwtW+nNUbNigxn1R1
DthsLHKAXaYr6zo0CBtrBjDYm7AG3dx1qiUtbQec8Ezf76NDP2tBHdsZMY0lfD0Geu7N9Kgaie9B
xqDmf1c20L1/NzI8zR1+kuOilcufpN6lQxfUlMNJmmIzlST/y9J6naNTBIOqNJ9dYMRzH3+KT3vu
f12HAS3TJy9FYFZiAUE1F0lnVJsUaUa0+cZ5qJ7bg3JmgFoFerv4nZymYqY67KetxJc7XN6putR9
LLSZ8cQ9iYCiULbsA+0nT60REQYJF8qMXAMU9CDaYIoFFGwiW6w/c5A+3UaoThkrpHbVJSs/nfYD
3J6F0laXZQHnIy1UG5pXzuXKsJqkKP33uWGzwiQcSv3CDUGGkb0Zytod9LPgLJfEPqalGYB/D2Zu
r3MiXp2YzMr7CusqdMZpe8Ezx3YgLtMiR71+FFKAYZohBElJwlj90s5z+fvZpiVnyTtke1O0PON0
M7NJPnKP5Ofae54Mc1acOreuQeJl/36XJbkFFk4cID4d+pCn3SokF5ddN9iq76YYYAKP+lkowhsC
JLRziHfd70xeagMqspJik6cZljGAy0jwPi2dj2m8Sefe2a/G/FaynVXNPNzGoPUdCGHe+kkBpauS
HtcOInCRN2grw3t2TEYe/yw4xTxQ8eh/3WBzJKSDuuhE6RvZRd8lEgIZjLQhooITLpAraUuC7qys
gsT6VotGd6jw5qovZ7tZPEl4uakLDjSil3eknlK3ablrRcqdfQkZFpTxTZwg/pw250201rtMeIZ5
XwiX7m8tzccmOq3KQc9WWw5I3WCWJyG/rW4PSgrt3yz5UT+1BqkuKcsiBonhhrgfnJ6g+ZdCLtnv
iLgs/MyEEterNcrtswjRcJLmyxLdb4bVXTdcCXsjeNIa+uX1FsBYYrA6hRDGemTiQaivrc4SYrYA
0fDymMvRJkJmffQfsnS6dbaCDWKnLUfp29vhVJoxi03BM4qg6Xfs4pw3Ugx/mq/pURqTBXDcfa9K
qlbF6Btbbbo6m1zLoUpqq1nfSvutC8WCAf3bbYLQBjnziu0VMGsz8rwdVfgaSmWRu7xB/ucarRRo
5kg9CdoXbdKSy3gtIRaKI8qSGK8gCuDAp9mFnnoKDQZGjWiCmcH9g7n7qL5Ld6tpAOHFwoD6BRTN
we/kzppa+2V6cFramn4vtpK0UBK3W0HHbJVIfMFAoMxc/MA4823nvvkuMZYrPR3wNeW2zkcdIUal
nVAnu/VZU71V2H/W76Ohdecs5RQSWKWRx9tSFLtqQoCOWR29JBz6GUFrZnBsAs0wRjsYmAxCy756
sxjBK5H+e8HKKxiGqkWxQIonbt4BvoZ3ejrTwbJ4jS/1i0wleFUk1R/uTqHiaywDB5LL1wnQS5c5
jDls22pBFU8INNkKcPI0RrYYVIEV/pByUyAr9zRQ91CnzAVE6knCsC+avQA+VN7H+bTMqIKOVgKN
rcsZGMpZentjPX4L7cebDjWWgzsnSTo8UxZrGOwyjcEy7bIv7461pgZPIDfxaPBZBzdAImmXFHKK
b6EJh9/6BZpZFGmC3tpMpBe8azs3LLZSK4Z8n9m7HU+Z2c9/Unf0u/0tAKhaQkHUz/gY6qhpKA/R
oDTgO9anNjEgUBvpe9o/VatmM1P8nyJPP5qYdz9pm78hku6SpKdLE+MGd5lnPS42Xt16KVd0hm6a
zL0ZSIAgTxZcSs7lTLwreebkMkSdfeH8Vj9UDBchtT9SVK4Gt/81oh1QzeSkG6+st1n1YDUGDtcI
kvLWFYE9ha2CUpp1yWv5ywVE8A1bN51j3duzhBPZU03VrP8Dq59cKs3QAlDhl/yK0s7Oh6frj1Th
MCRRkj2bvG7tfP/ytHX5GkKEuhjDQMwQD5I4ckxFwzCxFtjLPSdcSC7L2mp3oFUI6pKIZJ8MpRcp
/GtvYQ44QfZAZmL3bRZ9EriHj42XRu1pP9xt8JpAhPUX/6JTr33T6/no0QlXGFX0OaOUDENroTTm
t17lzktcb/JcGH2h5sKlkH/ERC7jlbYqcr9ath8B1T/JpLPrxoFpgpTJ1ohPVJ+MMUQKXxvykMGq
oxDR1iDn+sgeNpkyzXG5rcYJKIQb9HBaPELtAJJhM2bcEx5Mdhum+F/fysyTaMp/ObXf6Um9gc7K
KhqNsMGqSRdB2REDaAAQfLaaQNnxVSlkYWRALkmEQ1O1cV3Kl6SAMRbyjCIJEA3GFUTIGJkJ3haL
0srzTYkRPkTNmY5lUIKA5pEWbq/UbnJYvViqwTDySeiFhTRhMdS8Zee0lkQvKYJ8Pc4yY3S+G72U
ZOIPVrtfDaI5fXraQvr9SLELDd61lLgUJmIwwykAWerXeDusoDxkNlAMxx5cG1OwYD+ZrHQJdICB
Nb5iELX2Gg5pmrCb7/X8UXFxKYZkSk5ivoiIdP1E2RXpp0BnhEKihVWAgR2NBYKjj+Dix/stTc6r
40yBBqgcBGkITZ89w3F7clcRqeolHRFZLKvmkEzATnFr3rKggOELIEMJxyurQj6t8YQKpaUYiO6d
+brm/+3F2sIkUD7Y2eTiqwxYMQ2XcVydBBkdYfpvFFg8HrAqZ+8nqin3BMQdREeCttcyhrNat6Kr
VoRoNtqXXHtihx8JAUCkoFRa/R8qZ5VmcUfRcyjIq+VaDt11V5WYNSqiIXHMvAmUDQtedGQV0nib
MobLnJfe85yonRJ8D1bdmkoN/KwHqogOBCaUMJbjOxheD8z0mKEwoyICdmJVREfUOrnMKRZaBieP
QbweLxrVsElCGvXrvBzi4Z5Bg6xBuGuOlj94FaF/cQzPa5bJsgB9xRaQaazWF/o/nduXwug7nbL7
P5PfasqztHZhFdMiTSeW/nyNJ2btKCCYXwzKG68vwwbq5IHaz1BV+V1mLJA/qqNfbsKMDGjlvKFI
vby2TaMB1Ds0S37lRokPFRUygvGn42zS86uOl4WCM5fCFJZEgk1hQu44/nzWEJukzndj8jJ+eWob
XoKRBa8+xeEDW9YJrwyRJU8wMhUlx+Jke4E9gZLTZD31rxnQTNn/ilBYzLa/B5WfcipDFHgqBkUP
8d63U7Xm9xxdjIaMbz6lF58g5sbcw+XAOYarhsWbXGuLOF+uCAbLAD3It76+ukIGAe+tswYphu9r
EN188I7kKRNoRiCSZJ8rt16KFwSelQe3gpabV8GLTblE03Zyne6DcSYr1cS3biTMam4udr31lE3f
jPvR84SG83qO2V4gygfrMCVspGTlub280v7bG5MCW6gSPe8rIZ9QpSLyCUK62yXWg9AB1oUgIoca
3enLLu9pcOTS0jW7fNjBDW9E4wMHsaSs+cUGrvoUQKO61k54+Ty10eA/Smv043znVbiQovMadBE4
WKOFgBKr4skGDqXreMidsKn76p0vz3GttEyss3GqYuG1qCK38muus7LKcEtuEcH3DJwaCxdcxTfa
l+ZCw0X+4K0D1VwIYL1APQCIywa6BkDNObH0Fo0Hg67EtHTYbrqsG3WxtEwwTwuCxtPiR/sdHdNq
zmPDE5PP+cR3lJR/6o2tKVW4DI1GPDZKms7LLjyxLjFasepvbIPt4+87k0rkoScIJzDTzTAhzAg8
wCmO33WAVPb3dwVOKxbFV0vQycBs3aEleriCP//Lg7HONj5paBZjnUQ3BG7edncZC/F6hSkLxkkA
Avj5gjeL8BSjDxEnmCThRX6Rl60TmW9ToddmRqq2z1e/nvcxGINC8hF6GdnIR5Hx2lR82x3aSZG3
sPv0THsjDNikZjWey9a0yQdAUVoERuWL8e/Ftke6IGr37kgid3HHprxZA+YjMoETOOW9JanG0Bzs
YdRVXK3Sd5qFc2b4QSAeiz8TBvSHNsv+tLV2UR3gGiXsnU4WFKWFIuGFHrzi5Ac1woNo2UtT+8oE
QnQrAVIrTOAk/N/7Y6Spv78yuLksaiksOud6MbDYrL+ixZIlwP4Tl/XTxR2gNqLTDF0H1ppDSzV5
iY9jwoL3++x5UAjiyrwRqJXIsIv8sKQdwagwVfr1PC/ytaJEW+Fywom3AXBOgg8fARTHASgugXL/
cQMU9YjER2SqFGtUsPBW6O3e7alHHONePgLAIKF0BcFx6pmBZvO/5Kbsw7cCNh6P9hTklm4BnR2X
lC0cf8x6ysTArNFhpBnkccrAXzzbrUHxv26QcBpH0yVj33boV4cv2+dZ91imtAcOaX5hWow5F1KA
AlejkVbcNfmoURejZB4tKrkOomEVMzWpDRkkkOT8KMTE5yxLCskaJn2y+1olMThc4WBh9jrufJFG
LTbbLMW8aTFkbKToKDnMVWJ1ed8M6L+8QSXTUW1JHN7SLwXn+w2gXhuvKRzJJVo5U4blHf/zoMbe
HbApEk6r54GoRGEx4DXFzN7wr7/M+ztvuy28pDhziWJXST1hSyvlGO21rUKfstp8/+zcll9L8Qq/
BuHY3EKNITkL3Uhtvm7dM7sBZKMLD0bRXgVkzvEzW/JkRtEc5rs7qP7HUmVoFlrD6jpJUm0C/jPj
G2QQGRH5M3h8EatHz67Rnqq+sZ8/YG4vbsd3g8XIX3dXhfTftlWUpeIyp+9TetGQwuIvEJFlPlCq
n48RTQWqWnlCMZTr+44+ZSspoWB5UVtFPsddz9tCAy0w+8A//e5Ujdg0X1vYtROopxtAsXkOA+b6
tUAgphWH4NQ1o1Rj5I+wowpRXCUUqOX6nKgr7ESvUNuCrSgo62mA9qmZdDXD3Hv/etkswuICB/aV
NP6neI1XqbEr/KErE3clp92dOx4QMHr3mauIjwGl7h0qqYQ2rr6ylRS+gmLpkQZM+2GhgTr95Rgv
q2F0xZnyZOwr3hL5wvanvJm+cenAW2Nbhk+GEPbibFSxPfL1Jnr4d3NXpj5ZqFn9O4dMlLTzwCFE
8VAqM8zypamDmtz/c47azFiuPcPDBQbSzJGEENjP7bwvqIJxAQijdgjfms/3dS1oGerXrnhNSLng
qT1UlHJm1aQ+neb4g3W+ENv2djM87DmpBLKU0CIoaNSF6Vbgx7ytCUSFKl/cS8pIRK11VcF+6kxF
7ZYSxy5YjLjKAxuTXl1nd6Ygem/U5s/N397RjsSxDrI7A3flVvq+1MU/5tEXr0DgDzIzwGH8wf3+
GRzFU8oE2gtBaIEJ69HA4/tqWXHOiSqz/iTuLbVtis6gHf7U4Sngl8+CG3GaQjkB/69hXWGS8lyF
aJgWxxeCJqpIQHd39JNG8ANhf+8iyoc4wHZXo9O1b0AGv7pyS60JtQMTZrpFR1zAabhtyEAwKpxI
0/i75g7d0eWqHmrMB/7rvbBOuE+n9pLr85N0ahHUkAZEl9KV3LXRpj9V3NomhpZhjNnG9zKC28kg
dGYwqISuenN93zHPMf9LqB+KFSAIHsi6VRXjRT9195qjsGmP+3pMDcTULQkP1bf5u2qqkfu1GgVs
fnKaFhyCrQdYBos3r4gaIRqpJSPI5a8xCLCMDRgn+szSDlj0BaDGUTwLue5lCTqqwxqc3pEeqNps
FtUaEa1oIv3h6SYrwyOw9kGlxWEezkRnRQtjSnMQgB4PldIt/8C69MbOt9GQfUhlmNBBPoVj3qz3
z2RF069yMUGWovus/l1pmfSS0dXTuQhVN8KBfFxjwcvR4mitZOgf02um5cEQb4kUXHo6EK3eagCb
DBHYszl3wOavIuX2lDv6EFu5IY6oHQ3RqUmajhhAUZUIzAOoyT9d61BVHJGDxyPeQt9nBwF+ZkbQ
76aG0fZBPVICXZc354oR19nxlZ2ZIUE1iiJdIjG7EXSZMGoLNTeBnWQvotXMVlOdsunem0vOQ8MI
YGKtTWUXBktJb0Y3KPFBEaxKAAIeQO8XVso7PPeQjxVCtN5ldLSZ+E66dgLkV1TXfgNW1kWJrVyl
4rryzWJihZwghKAP5YFj3OogjOVIqIA0ftg7yyQQ5ZnRGUg+l5qQsbRbuu7y5ONcn+m845HU6vLL
6Vr6KyaJIzrahEo7WhBX1QXu32eQi9W8JJ2VQSnvPNuOZbTqleoNWi1uP4ij6Jm8I1d6or9x1W94
/W8ZExdfT6cBsR07uvO/meBa64NVNwXw1c/Pfay/Eu3p6rkyNgz9Uy6gljH9F+vI+m6g9rfUQTx2
LKmgAv6hyn7ijor4gOB5+ykdmWi4+Sy7vSkJXORj6+JdyLQ3X8nAdNfgo6LDnKAWBQj98aOPPAlG
tWqScCgtWoDqvAhLyWYdfRB1aE2En1BNH1f9T7uen7YPnsjNYz2geUVLncAS331suBcaDX8FbIOi
PStxsR8PIlxx7ThqBtULbxPRHP6kyiV/ilFEEK0FGFGIM7xCF1C7UiCtRYyxssqy53+F5FdHsJ5C
ijutN8b/1HHFBKJZXhOF50lyflMVCFbMO3/dwboeEQ3yJfv9UrBOJ7bXw/mndK/BY4WDk2e10K8C
gUS3SmgpS/sHjCrHtn3Bd6WMTKillJQmnfuaQCAdIwIwwkjZXaFiUdPpFvffQsbprY0qZsq8QYLJ
fVqK0iefMGokWf7K/tiYG+wcC24z9j2+r/hiUdJiZw6o06/IURgGhImPBFbBV5OKfO70E1KjR3NZ
gkJrExjO3T1H6Q4814Tl+91nQTqh1lYC+Pq/WXnjgXGCsaqOgrrzAE3Mf8qmHVjtyygivkgqE3Y1
Dh3678U9x12b4w15OlmyOPqY4EzjKnD2WgnvO3zAkfE4ex/I1oBmujqCAUYOCG8CvjZIq1KxWAv2
ANs/0MoLcp338Wklrt/jqVdJfNrzYQDAR1nBwMg0Se85Tg72km2eI67cBP+pnEh4x0fuIP6Ov+9d
sLvbue2rlFr0mHAKLiKjz0tREWsjHVVSusBMqLwiHJtiIVjwK621F1JQZ5WDBOHcXeLZ6IHbsJBv
pbLYcDCyx5eCJulsxDbPAvWIBIqmEpvecrQ+/uyeNy8JC7Koqtj+azqpl0smOw9k/A1nkXPXvCO1
2+q0lXZeFy4oJOHBQly3YDkjDp0OoUDMKpL2WtBTWzB9YYBHm1BFLNSdxEbieMha6iTeVMxGiH2A
so7F0tAMrlIYgJIN7h0AV2yftJOuwiuD0Y3Zdh1/DrC3n30wzgUy0ogMLmT+umT4Tybd8A25z+Au
fz7uUAcOU1XH4USaUNMtuZ0AWm4Wj068DNQhsQk0tL/Q3QaNuQTc2Dut5cNc7JcSYU6VYJG6QtvN
2xRqCasdkfwIxAqbf1DXv1xjm/tvqFl2YJwrCc6MviEy7bGTdkcS4pRwouMOrI6fSKaw/sPZN5mL
uIJH7UVDLfSuQBqy+Ew+YJo1NHhFagWwwZ262SlchDEj3ZwP9/s9LomMBryNADKsj+kMjAiR0+0a
cKKkQwi3E3duDPWBMruAw6dZ6StKZr0PtWBwt/bLwO/0JLMh9+kmd5hwep0BmcJP8YvAsynK8pS+
4G53XuD0egsKAC9IjPtj6F6P2gq2/vcSf5/jQXxDoAttfec1de3oLzvzXnBA/ochWl5cLquiP+mU
UPKSRD0X/1awJ13D6glNy6PuOTk8KoCRYyNYZuwCorKsg7kOXFOfF1xGgDmmPhbFHjm5hC+ooJwt
VsPXzAv7UnM8Pg4CUdq/ECTTnm8yLlc9dbF52bfBXKKBti47abM5nMR/z49mMe1tF4EuV7kWCSlo
xELzF4xXCWut4BL2U/uKRdyuaUJlf7RIs2m9ht/INa8GDa2pVFK4Yzf7Z/5WXyuTjU2AV9vFSU/X
a4Dss1SUKTz0umodYs1gFZnxduY6Sa5SQwccxR5/80tRxn75MbDQN540Ft6mrNY5dMOPWMvPBG5m
Dw4yuyT0r3DuFfLMq1fL3eAZy7mO+iMWjH+Fc2AlXFq9H8X7N253pgSjsvC9AY8OZQ6Fvqrf25vD
t94DSeijO5quXSX7dOlyZmtZoEFbULTF5FwxL35/sy9XTx+vD7VrmCiTfiuz/XhIFGXX6nXIF5ln
CeEqtBhP+eerQvROjBrHCZ5udQwIKTQrQtV+4BPwtomgqVQnbkZhh4WIBiE6acnLqVU447Bault7
QVwWZ4st3mNqT5SdhaCSvBKk0BjO6pz7CqKvvyPq2ZS7E2Q+AKUgUe1vfxKBh4Y2Vu7gTS+LoN0f
AH4C0dTLfwh3Lkt9EBMmxbyiNRjI1Q6ANF5xl0y5GCunMCbB2ek/Z88ZTgB7Xxa9Y4bOu4ccOT7v
qFQeIm/lolzSb9rzOEZOHc+RrUQX5N/kkgFgXRCbN/Eh0WilBN4qhW49hRyJdSAZSmEdtjXCKeYT
26ARn6gFg802a7XtxR8Kpz3vG23Ujd/Vyw7E4CSwoRLToTNpEM1uF/F0NHw5Phh8noLrFTUrdFw4
ztahFnV9TVyXu/Opp6Dmwk4nbC39jHdn8rcgaX40K7ldr2MYBOs+sQag/EOB1TLUqxxYJVd1WCsR
Ligb0OHjx+LTJ4zeHp0FD29W6uDOLtuoszaG/Ky1P7OCSgCZTgnwpCd7jgxoa984alAu9k3a5MWG
eEWYqwXovJLFSsByLQK4lYPUgz647lkPXRRIGV1Qym/Y9bT4DYCNEq8gWzeTFnUrs7gCRNRhgFzw
YtTPt4pzl574mVwK3zi8gX01OhQqSv0uMQyzB2pzMNQU76f/ql1UYz4iK7r69rbRSpuvdYIGLNXX
19wZsK3eyiyNFXcJjgAdX5Xq+/ydQ7OQ0OM8K3VV+4yNsQlOz73gl3Nuvwcrgx8bnSmf8+31mKeG
MpOISQ52+BvjSZKyj2LZfA/unEadXG+b6RSRK39vQZ7WgreQQW/4ex7dRizmhTvFcaSFoe0jMzUz
fsF4Alhm3za+GtXc0iFBvkoMoIFwGBuQR0nlqVMoRsUjkEH1mY0klSt4x/P8RpuzEHZBiWz8EhyJ
+PtNsPTLYif7IMrAtqAlBHw2Zu8unrwcgvngbEn8lK5SpHVcC/r39itpDmclvS46BM4pqeSgoAhD
02zuYRdco6t/O8hfUptvprBoKmvE0GLUdxnguhU6lQb7iZYnoQQUmbgGnWOIhZfntx8U8MK7uVNK
Fpd4nXJxMeI2b0zil1dPFUJC5GRi4HUVxrh0ivPj/ttDvHUY3vwcURTSsCLFeW33eoc0yKoUGuk9
zGI8twy286YHvRwsLKsJgJqZ7PlZiTbzVUROAdGTofxliaYTU4CayNBbLkQP/jKXIZMeDqY4ckDP
L51CwiHYB7W2V4slSh7XTEyvfWC6CCIHKb92rNZ83bbpvg7dZGs6wly9YkPALGiYo9OdA0zfXBQC
8xGSMCc1tgb/bMZ4YcrlBN28Jtcqg0n2eCz8PJgU7PF4siunwgSzXNp5P/cjs4f2OqP2EqNkIHZF
njYtTCzlnyyymhidpqBALICji6+g9bLQhODwZDqnXzptVj0Xcmtj/kQ9c3dFo2PDm8Up03xNtqWC
GK+T2UnXXfy/JLRY18xcZnyrPuqhy+Ln1VqdkY/1bwjQfu0Kh7IJKLsWSkkJlar9xCMZQsiryGiP
WPXluXpOXFBmCUxEFAff1SwM/z01EmM/oolQtAtL43QGE3+j6QZi/DgmO1VPgCckPSSSk4GyfiWk
kHRe3ClSdWFqjjxwUtmZRd6p1cgyJtAmpuEZLb/EsIpdhS9VO6i1Fst/p/Ye+0awlkpCbqym+I5R
bCp3rolQYQ/dGyH35pDf2x9SqXdcW/0w9VBJvclDHsqFN7zNxPj/9s3vePIjvDxpUGXxZBcUWDA6
njhgsB3X3OchRfU4K2N3Kj5aW0ZmmZa0CVikigafDrbJIiz8G3gCcdTTQDnvz3zUA9pDdSHJ3I2X
1I9IyqeTD2vTqZ0qDKZZDy8F9cZWN1OIm88NckA8fe7n70tJaQCM5msjQSfQ8b8jTIwMtCRureNU
1loNfiis92g4mLM9+b6mgPTd0Rx1p9tXC2x+F0c07e/urlR/N8x7TwlyqqjS24LkhhmoSWehaLSI
N+fIXDITqkEu7JT65lKMB7MbcM1NqbrOFlUvCNMitanVxTBAb4mLQbSJ/3CM9gMLVymJzPwSPJ2R
EDlBa6sTWUBjhVhDHPN4pvkdC7ecOf/CR4DAkyTGFZN/dVWsN/B7cGTvjmc0aJLzJogAbYjvV08Z
C/jKKSZt0bAdZzttc8alOZ0E1wfAEimaGC2ZzaadxnqY+XwEpTPivz+T59Dgejn++o21VO8ZLwPx
g65UndF/92I/bdNEzmItnbYs4usMynR6gQGgdRa6bPj4LpDbeI+Ky6lA7P0InUJa3tSIbhLyVESo
tv5rUXnPUFjsVsr4iwkdy0jvOQE43gO89UjGCHb4xQuWW8iYKKtF3+88Ld1PnKdZdhbGp8IgMR8k
doH0ZNnYqe9nAbzVFn6n46DjJP3TMB8sgoRi1vPFSQnSfSJ4X8odGAdLFmO447w9NAxHZI4omFX8
5X60TWLkTcNuiCrkXZtoeF/r4dfOOH3Wbje4QNvucE5cW8gvlYGY/W3DIlHEn6UMsg38GWEqH+w5
0sXS+u1selqs5E5U2MHj/zeIUwl7KhRO0N6zf9LlfpUe71Eu8ECXlKuZ810fHHbw5celhb8ZIHFG
o69YbgDuJsenadXBmZLZxtjYP3tGPhDICi38yd1rBNTNIgIbb1FKDLBbLUhUQqjmLbE7lTq9JyFl
uXvsoSHeQ0MxMNEBwnigRvxVANJduF54Zyp3iwq2VDwA1kMbW/na7sRPw2InE+0ArClZEF1nEsP/
sy6/RoSlxJ1pBOyAvfEGrp3ByVhvmtdBSn87+Pxll/418infthVwbQ+8IVFcYz3wMbJsFHGatJ8x
NDNL3c//0K8rTCnerwiXZ7Fmrxc2pT5y38Gr98WQt0hXg+7qPYJL6VyTgxaHwJYAjP/T/okS8zQm
MmRyVabpmfTDN+/Nc0wjt1QwhprWzbshRVUzN4MjHeYsMW7WwBEvJccRt1CgFivvRgVUBQThO790
uIErfq6eoEZruxEM2Bbaioami740gkf4/EbE/tgSzxRbyUuPgxyG/j+M87IWPbGP3iZPB3S0Qv0u
OX8x1U4WRKDe9FdBwg5NSFjFtcpdCDki7+xuaOrVC23QJ9HTMM1CJ3hmxNA9O1iDx80l1uTMtQve
cpNubHiVAUzXgtzxlDx6J3JhU74THEni8815rgA5ZiRkHEB2HzcBMa0mbUO3NYqHTBipYakQbajX
auj2/Y2sbl2TZaJBNVqoYQMRjkUH478OERMzYcSKSRnGoLZgzTNpFDauVL7Xze7NI2T8IEZME0g1
sPC/FYoJvebuHVyi3Jo77Fx5YnXnpyEcX9GRqzXp+OgpCWzbmW45vAqOkZ1Zfe2UW9DjuHEAHPot
mi/6BEUN4tC5rOMipN7X9J6XtqJ4l0MLgUNuWMoAiFh4zVfeM56jNj61DPX0pH9gvTdKCxN1Uyrf
i63TFuKgcGAimEA1ZiPAyBHmQYGGMx2hJ7cY1P6jVJt1m/UV9+h/ld9hsy/r78E2W0ILEIts8jrT
T8Rf+verL7UlEb8Y7EL+AKeo7FpBkLe/xlNRB7694i0CSnjdyHY6hWdty5gPCZ0JYK3ogJTau7Mp
UCgFB7O162sKqYaHUjGM+RNPOYgeBEpNtN3nlux9h7Zlej4h+HiDtyGPBbM4iHQ1E6V3YnNf0IIK
i+X2klllZKpicYA3o9aURewy+ZIWyEsMwyhTrOaxshxlwLncnAxDal5RX+RzOKu6Htf53AtlA5Wm
/aQ+URd0iPZKd8b1xR1gJwo92/QGVnpD0RxHN23jxvAmRWkR6GjlDQ+6vYujqyzi+dKZ0kQhZivd
0ZtK3HW1s+Tb1b0P4oYR80Jpsw7vH+HRBFRAbuLg/YzxBkF/wsH9F9YbyPM3/xys7RCNr6okURB/
KOne2gGDlvY+Hy3NMXxmNTdmlluw45CCdVn0RgIWImkbtMvW2AkYWAdHNHSa0sZNkmauKl7NduLw
vlfb0/CuwPVZd4FGdRkN1jeVVJWkV1Z4SLsFE/9sGlTQe075qO444eCUMN9EyNVrcsxN+gX6PWAZ
1GPYNQbI3aSUpV4cpimzG4KrvrJTRs6o4c1JYaw0y0ayvFcOb9DQqDywbCn7coSdcwZRslJCXeH1
ydaXTvrseM+ir4WVRA1g/LlA78otx7bQMOtuPBLVpLgjjip+EnJuosncg8v1qtYDvVNoQaccjsc9
o/IwM9vfn8M0nzbHig0TwvIQpTz122uro2oY3aa7yUu9P3+BL1WozTnLDgKVyifyrzuv2JcHqDK6
KvAhGzGQzN1aXEHMEg+6WBF3Tdohi+WUX0H97scWKvCb+JZ8UP8H9ArzUh9j+jhoRqDOmfj5UBox
tv/whiFm/+uskPY3WNev+eFI6uHPz8qyC3OnERjGB+zJWFNx6O9IQfws9iyE3u7C7esZpbTwwD0L
pPPboMTcrnsXPu1DjdwgYLKnkp06T+3td0reVeiqSXQFrAf3QzncBieA+R9x7bWLGRv3RZwOyPBl
vurjGX7F9cnRxDWaQ9hLleP+17yIjpGrTdSzgmfCBRZ/50vpvJq4yjoc7Y8fc+PcfISif07wtEmo
txxgkOahCMf6OKtY+v9awofgfsEq84yvD7pG3V6BP4p4IpA2wBk2HhagUq/hxpBVR0ZyQnLVub2J
397m+AkqYKGAgqOENn4iJzb0QmE3JfKm/yEhknYziRrdm+1pRTtK9qnYXDopqEd2fS55njaVNgEV
ZN6VU9IvSDpbn9e1zB7w4QgnW0P5VGx0ggIXOuytqyuQgBMFujKcoUV2pWe5duRMKYAs+t1rIjsE
e4bL7hu4OLCBKCRLgm9elL+3qsYObBjrlPWtISVC7A62emCBqok2lqfAChlv3QAUf9ID9U1f/mAm
hIlSnCiEV4oqpGE8iKUodIUEMT6OI4aC56fhBehidnfB4hP3UD6tJ5WRfRzk9dgaaijFOWAgnp3A
1DnSUp1LSonIS+ehULtXMgNQ3+XJVdsfInl4lxjDt8lUe/Pe/Eo83JQYfy38sqitBS1oPruyEVHq
DqfUCqK1jqY1iqfhis0tmd/4DVorQnFUV68w6GPu9VJ0W/r28/e8pCzblKuj0K0uCH1F7NKqeSev
eZlxQwdPYEnmKVysCjMNnyxzppfZaEOBIrd94r7Xc+8zi8IgGgUNsVatc5YuIkLx3kCmtiUqxHR+
4ExGK1+mMChblq0f/qw5WySfXXGrq+ta59MkwxAa8cEK8NkH0jSAwT+ydkrqRad4gbEwaaAizgHJ
3u2YcIy69gbmYLWQSTwEr/M5MbLGq/4LnAOEDij+rg9I/KmM5zO0fEF5w/JNhCBbmldlAs/kodt0
mexjDjXnszjzMs/Envmyo/G51fuJUsKN6r3kOiOx0/C5eCIP6M91+S/8uqNiBIUdK1BuXVPixajZ
bYEl+OrqzrHgWtdLFlUuAMuuLlY0JKWhDgPxFBG4jW4pp01kSp9z1mhnSKHvQIsraWg1fkPcDSG/
qDJR07rA8oRy/LK974nPIIdwihkvjwwwH1WUru9CXPT/6rVdcKRp38JYLmmHUWxE5euitSETygo0
FkY9PqEw8EmWq10NwrLlok0lsy5zQTwB9KcNmFdNwCnDSY2QNQry9IB9CjVy1vRrqQGx6gCz1yPK
N/TuZW4iDEVNOSuxe6hae+Waq/Ntur2myFQw+479IX/D9qeG2GtxPWbvzjc3e7Hr6bJVU5gYW33g
DLDfLI0mEnqN/IYK4HVjijmgbwF5J4Tvm6LddSRoUIX0R3zk25skEvJ55lKg5kpWjNED/+inkZjn
ihKKffkMLqBFZTwZRC2UBrRNY2tzwLMaDENZ+QOFOZFl1kkuful1GzFM9o3dBaUrKEOD1il/0mGT
qYB7kFFxto7hTtM+VzxFRJZpvxhMGEwshhNiJubyGIEEoUCLvtBFc63+wCY3N/QgzxtAqt2oIWFb
wN7208Wkujr3GpOtBIjfadTXwwYqwR26+wJMarFRd7LRPt58ObWKL/ypzQR0Msaktq7jNqib5MGf
nB21Zq+z0+B8Anbm3dKgoRDfSeImECcXKxR4nop/hUQguv7jAZuec9Onu3fw70AyIalu3cmhEIUz
v1sGZzvF2pcqtz8uHZm01pJhnhqk68OBt32tg0AjF96gvUdmLvLWIA6SJNdxSN8nM8K+8JwSWtdc
wBYdE6inSBQou8wu/7D3PXWkICGkwHHPYdtWAFoqwkz/pCtsRKtHz29sZUGT7onawQ0HF4o99n5C
lx0GlbutNAi6+Gzl6fct2S7fxlW4ijB6GXFXzUGUYbK89dZfEqbmnYHIABK4bti2p82Ixs/0NRUH
1v7ZsU60aFrv6a8m+eMHEN8QeJaE+G2OoX6qD90cq1mVK8bRYqtjQvKE1sKqTw4a+unZf1fnoRbp
vL3sRMrbdxSf1wb1fH2z30/e7VPz89KhPsIV1NEZmmoXTpcHn04EfAVsjagCaDQMcILqY0vOgvHk
ZYQbtRisbWTcDkVpAUFGJmwdh1emGGo/CuCQLxtjMEQlP2yLHPQ9+DRkMr52HwcOLTVrVy035WV2
owiNmltGgyoJQxXgwTzjiTp1TwSCeg4e9FFde48R1ge4DEv/ThItC+4kCH2ywpHuCG/qAXMPIv1l
kBkDLMXYWlJcJRZUN2UugWSgJezW7jVjKuJw6pLse0LwxI1OAxaCIGyz5LXeTsIhLo1kF4EQZl2C
YaHrY8/AMx8FnCBNC6bZPypchLk/8kAAx+lfn6SCIB8eoIRgA8gds29NhAILzDDJeLpPA6mvLiSJ
Ue3SA6wgVJDCTDAs/S8dPsmO0v0SCUfQ29oxJNgR1rXGJ8GwUldtgJIqAZQWjTpg2RgcmbITfJwu
sV1A4wVPuTPCFPItqbcFn0xwIa60Ge42oCt0iwutxQ4V56H3I/K/bn3YR7FvLPqwK/T4OSI5m4C4
gARObnnLEQOspMEPNVKImQ0WmF6uYIYcxo62VFWqB77B1+MdVikD4Pgrw8+vYpUD98PN0xvvbq+H
OXxfItLNVDlEW/hSkYJBQDMqsZCqSw34WX/UciNHkSKpsi/1o+VIEifGdTRpDNmtUszky4e8zSH8
dTyg6WIg3Yw6nMXUEVYQ0dIUe6lT87xhfzm+rf4wtPT8xuxQpEhKKT/6t/5OnUGjJTrZPUnmvzZG
+InI6ZU88/a4vj7rqY4IxyHvqUmd0J8FfYR23c6/YvHvMkzKlryo6oPIF1FREKZo2g/a2q3eCx1r
hpa+KdsIzCY+DMWo24oaGOe2vzTIzZdQpp2BeeLBAIr4EWMKc600arFGeKmf7XA0tb9g64BEX3GY
wkECFauBOg9B6kexEicYDiwIqmvAL4c1lZohGWPh6zxw2dAT5rmbyF6eI4zULs7flm/NndHNWDUG
bBXt80rjvmLm+0M1vTk6M659HspYVnN/6JqyEfyRE1FkAVfLwliO/qkox+Y61y8lcm6zH+c88FBu
XfSpRSgCPgcB9jVqlOBIrattJh4c/ucgzO0MRZE2VmW4tzEbg+O3tbU6KebUClT/v067VnkHr5aC
ZgEc4LirJc+zv7/wTAsGpsEEfv0GZNZ9pL8cLCPBqZOH91Ueo+6T0I1aAB6Do7qklpbyWiMsMBFc
fs70LX+ha8t+2U1JaPInxBQ1cqlV/BpMZO4/c8K9g0mg+7++YUOlAGFyW5R9yH3YilIJtsZ/bLSp
tbGVJ1+O8qSBDbsJKqkRHZJ4QNUNRfiWUyyL9cp5DugGKICM8j52QaB+eJSnMlsOemj478xiNbjE
7367Di7pxFno2gY7FIH+WFzPcemTn5QcBw45JTkpq+WJPteRfoqUfIY4aYL0Fxrn2AEhpL6ttH9u
KrqKcPIhF6R1oIs79CS3nyw+K79gJ84UJ2zGxh42bP5Vad0EMf1wDPTDjp9K0ygmDqgTEWA8JKPx
TZBiuCfQQy5JDQymM/aQUJQoDQQOI17eJQMnxFPukECbGHqO61ncC2XZmlUq9g6UC7uA9R9/oHF+
CJEdS0nqjv4stjqFfg+BwaHGxDQLHQDW6wM9oH/FUEHr0tUkWQ9eD9XeGNh2a234M9husfFEIsLV
Pa3uG+lOx403Ds3GtUduzZfj0KoMG7NJ76gi/z9Caeh8ctr6H/d/jG0nQL8D/GcFDtDzZBFka85R
NsofGrEi0LBe8aSoImdW3o7B2oNmdA1+iJetZwKg8z1b3Fdt/VWZnNJhjHImRGWhptUBWz5OFWIo
MTPg26DWTtwlFEUxG5Qef5wEctI3vue+UZvMHNB6zi1fdNm2CFSvNs0TD3rAgued8XtkmVpuPiXe
hn+CLRpNsW6Qqr7Dg5re1CQHoAB7icob1RsnVmCNOruxSNXFZZVS9hb8lMZaRV29UUeqBI2SRpwj
aTgCDua/4Bcxa2eKhnVcESHbWXcJ2Lnsz6g14C9pi2EE/CSGCthplfUADSvgYf4BDZYna2f9g8w2
fIlIc+TEzfky5b3jyZfl/SrRvI4bhm+XsXtPk68VhmlcgtPxmEp3EbivB3FfTg4Pw8cpUbYi/7MJ
mBp8QO2YI3AC2bkXCoyHhaE0Y3h/IGsAJ8X2uewzIM6RoO9z/GOok9FXyG842Y3XZPsqGXni+pud
gwuFlDjtJrd7Fsc0C8dYfbJmh4hnQOgPBFY8Mllp4HS7f1Jrrq2jIYg/9hZg7EByp07BcBdnZAhZ
lE/Y/afgStBFjXkJgkMCRjHyX4b6dBbBXj8LLF+/Y/wrr3DBd++yOEFu3uC5XdwbvDRK+kgnB6hb
lC4U+1Fvc6RwZw7PU/RMMmWDdQRCREnHA2+jq7DG2TJT7PDyAO+j+aeSYlzquPVWLZbnlNWOraQe
hrfUtazzN1dvayDLVePH579NHm3lscA4BrqR1SiVURuDHuOqNC+Ql2J1AufSRH966PpXkjuTmOT1
SQFKPi4yKyDCYk3wamnaPtW5+bWf4MGIGkY1+iFS/RXXChLX3MfucaiwndusbT4oJ+Cj8EtcDEbk
VXR+Mhy4Hcpdj4CaEnNagCAbzESWEhMANLSEs/Tk+9DryxIDIV7/mWd+gEuNzC6F4MM0xrYaWVuk
QawRVMdjZwdnx73hurmA78QdXRBECI5FvYmEOfxr35hhnjaIBOj52AUMnKLktiBgKmkfYo2YcUJ0
fCnJw8B5nciOz0N9X5CzVsgXchgD1d+wJ6FWbrtvPjlCRRRkuSjrfJjkckI1y4M0XmyG6oFubw9U
TpifxVRHsv6q3bOwVmoYYkZvQRrRdvFCruGcsVnWiYAUWWbUxpTjiuQpSsT8dAS/mPusJQywOLoq
uluQ+wmTqUOCK/Ufxph2vnitClDDa9cl3EYUCGIlJR4aAhzRPoBc6CRrQ6W+pRqsR0YcZzcK0cNj
pGyUec6gAxWgX4bHWOhI+NQVy55NVdDmBCpUaYmt9J+gOR07DWVtiqzkVhfUJgGc2vIQ2MLgy5RE
dLHU5aDOTstd0yGM9lzDT4rk2xc5U7+q5/32obYaG9DhaMgR1hVrfLaphI8wHJVoWkcRTvHIFgTa
CR0QuQU4rbM0OkkeOejU+RnKFEBbi+qvurjfkSVQKI8Kh7UpoLM8ccMePm6fH0O2mx2JCgmIFbmh
X7DHl6+di1ifHeHqdyngA4C91b1+XA96OzI2Jtz6l2o/jfu7HpZ/rcX6CBWSM7I7np4ODNTGZPl4
Txle94nUcITSnYOhVOITbbajCqMu/n2fbL2S9BIYyrZoU/O5Jx9z3ilDq2jvkyGPhx6deXPQqL6C
Si6AFukkKnm1jRonY2o4cjgbT5q5CkMlLLoMR6Is9VW30F69FIDQYKIs53qdFUVjVTTb1cnvmKeh
VjnRHOC6IsCfHD6eiBc24FSny63psp3JdkW647RLKcjnDbtaC3txbld0P69KbJYyPP+UO4SpUTAt
Jw55tprwPxo9aBh5CM0QnLV3K+PpXIJQpSBri2vYHuFvqD3zDKnQeDZSX3lKngryYDMSQtW9anRW
F5MQQGOryjB8hemq3VC3GehQFttbQilqclUhxQCkmrvu8BUISfa64h2+xaY+PV5+jcJlVsTr5Ld0
Qma2pjYt0oG9eS7X0caYdZycv7PSXFdjwpiu7AFLgARf7wQ9JEQfWKwFdaqMOjre4wPBN2t1AkCZ
AK4jDhYw4N0mpynBgjXe/SEj/3g7WhQdUl4mLiYTOnMUqiaSeHdUMatcBEmLNd2YutRNgxnXLv8h
5KwWcsNyuQM+uiE4hFFVrDMdwrVrRMIyUqEZYCQeW1jGca8sZoDRFCcTxxMdg9ommaJ6VN1cR+tX
YRUFyKuiXaaZWFLuawrJQMhgmPEjKeVx9/7Nvkl1LQ4OXjR9nIc92enM8jYsv9787tqfwjfJ+BW1
h8Z+XZPwS/lrY6vy6mO1+I9zSfVYoLQ9KbOBhtDHH1K7ro1uX+3G3NrV6G7INot+AKkJsDP6xNO+
T1KllRNLMdsd5VxyMpkL3HY3HINa0+Zh4YurINKImILVKdtIuYZQ9vKJhk1qngV2FCy1NojQniD4
l5LpvoK8bTqvIDy4Gtw1vV/nm5Y1IabhQ+1T/3Zs5DbNi0CQfLxVg9Mi9zaqXP9Zlj0Ljih87gMz
Svny1Mg+Hfqacs75jUjOoDusUJ+3JuRidmwhQwVDw9A0neCzIKyXBKT6yNXCM2q6Twa2SNz1xRK+
GkNV5LDxaziKTujdyo2p/sKbSzLZQlEI9jotJ0VljLo0AzMd+5xAdXm9oWdYUnvhVCqJLp5ETBHy
eSJsftiFDCv/HUhYyssgu7lEdH8tVtryVFiy76HuUojlV0YaS0x58uUD7m+6yLevp8IEZ171/imi
mPh+CAlEX/K813t5OmqIzQFWx2sBPmF1KCE2I9piAaNiKcdX+4pSs2AkNn3O3CfNSw/u/E5Rgqb4
oIN329631MXvjpJBb+o0qwsNUbXtvSNARwSxQFDMTUHuXYf8lkLGWNl66t5vFVzscc8jerD4zIRb
6ben/oXYsC6D2mP2CD4+ywxvRYM1Y+fRkVhjsu8EykXX18ldmBZmvLybCGX4+XZ65u2d7pSacY6r
9Evi0zK9tzzdhJ6+KDOWyvug3grSarh4JM8nLVwbcA/PDlxxxsjALDrghW1fZV0XAsghRf0SlrBc
WyfWO2P205eYzLlrfuLnpg+J/AAfmJNjkJJfRelyXpHvAxEVAMkqqcz7c3R1T9OmgoHFGxcr6c6o
zbrurkdxe93pgp8fmtrdrY4schDn/8ZXMI7fwbfyJYX7EDxaiFnJWc6tTFA7gO1qOIN+tgcV+aYF
nOE7pDIR/WmkH9jaI4yLvWoTAExMAwtgEUn6Lc6JfpD8D/gsd7cXzRYdQaxkhthTNeBl8Zq2Bq7c
xOPjjL4XimAAHA26UoVh73SlFSxlW6w//XmjMoYwBllzbyste0vRiEA8GgEmfYg23VPPxzRGHbW2
hV8wxYJguY50jXSWtO202fjzyXwUzyHz7hwh6yymXKUL09TUCoAALg1mRyUxUangUwrBXNlFqJHN
SdZgWpsTVhp5VTxh1qIw4WaIrQMDG5TqLzakNKbK+paGn2lys3MVu5IszHclldO0RTD5Z3W999AV
E4RDRtxUbzbfH2fQIHlRPT6JsZI+PXWxeMzaQ6nRx66ZrA/xN/6g2js4dZZadWiupm4uBXOj9wZR
HHoJCMMuaZS2O+BlPt/xf5I3cwFHkhj6UAEJ1ziRF5OyMeteodVsxv5tRXp5alQzDUax60e4RVgN
wPn2LRWKwOCzD40RbFOcc16EbZXY8gyO2Myy7y7BiMjhq0cfSwgYW/v/kZUja1aj1kDLcueuTi3p
9Or5QpGtpO0C5QpAlXCJnTWgnzI70jaAvMJQfm/8sQKIugD1+KUI/q2jt40onjeuTGLSd9ZuuYiL
qqvh8mT03T98A/Q7enSjMTCaUy4aoYbAbpUga6hBF9AQVb3A+0UEPLT1Qsd/u2YZD/iC7QkBGEVW
C9X/gWQxcqMDJ3ajKnQUqga+MevFcylMQ6tuK9YKWutprppHFggfMR4Pm4brLEz/mHb183GFs+Lu
91H7TPu5LRY+lgnymWM1roNRJOztc9P5vLFpEBh6OJ09Jx1nS2qR5oxbc+DUh8GmNmAufntdm7lV
rL6jSo66B5A9m5UpruqEXpmJCAMFtqxgAJqFRjmU2zWheK0yQ1vPgyWJkQSVZPLpZ0KrO/La7hoE
86DehrC1eDbHNWxTTU6f7l2tnz5jDa8iMulz3leocPqYP+zZ2aNoHkzUY2dycKmKCDQilnXM1X6N
zpSg3bWF/OeCH8aVn0F0RiIKg8UqdeRs5y+ap0UH5WyessvCAtUQy0ftPPmuUK5o8InJXWiJD2W9
LeglnJw1fWt2DNGiHmHLF3H1OgwNcPemTeqjVj/aKB1zEZ3LPRLa5CWSbfe5PuQ1BVxhmj9ax7Cm
BCLJbRASt7VaO04zwufTmrW1jDl28TIXSOmssSrdED6gio3/NwB2mh8sTKnfY/i3PqrTTVyWj77/
yDkNzxL8mvQtSPcf87/4C8TeWBA8em7Q9gYO6MQfWLh9UKqv4PpzAnmwqywnL2iqE6YrV0PuOv38
TRsRN4+X7gaE/OJ8iHDGK/TTOgIDtH0th+YJnnFeFG0mACzNH25UsgrK/IzDeYXXt6f+KYc383kv
Neeo+AGRn3XLDg3gAZ9aByPzrpERs/jVRJWwTdMxCdgDbMRQ6X34tpl/2S7cTlD1eAM8lA7BxZXz
OURPQxeNnqyDLgVAxkRcnmWoUAZs+19DqApSkTqQgK/O/Z3MleFIvfo17WOgAsr7ef1tCYa5243w
8u1GoRK4aE6Rz5k0TB+4oCeXh2q2EsxPGjh9RAtxVHNhiH5X9+SKFAhmEctJgOZyz28shm2SCdSC
o5XPH2eKkbR/uCgBGI+aisF/fthOvbrq+jkIzrZiFNCn6if6jj9WT+4QicGc7OU1etF7dMIa3iKm
u26Wwu0HPfcZLsvNEdRoLnkoH2pnpHch49BhplQfjrw+KODQE0lrI4WutM33HUWjC/d5qKE7XyMS
W4uqWFQGWLBjVeaJ8L3fVsm75kp8x6aAgLPmZqRSeSzBrd7tvBYon1QCO0T+qBdUqwXxSZJ57iWf
1GKQp5wmVaFujFj13t/5ENPTPqHkD1jcvU6N8SrrSVJbjiEWOMDKo4G2Updhl/lvBXJMw3ftBvcE
IW6uo2wDbCvDxNQLXBzi0KCRcL7ZrxRObroY9GAUzuG7/ihIBsRO2KL50p+ZC0dD2d3tH9bFnZE0
QeKV/tNM+ufRvDHrhWiWB4XTlP34iWmQa0TKbR0Jk7rWQ9id+tB4hTuMh+4y65A/hahaZmWp3Qlo
JWUVRtwdvWLikZqVAlP7Vj1QWhEf/khnmFdvRbAargYW7NKuKeGtLCGUBz45BVecZqjd4q0sytom
NOdvfVVFtLU9cH3Mduv/eZEySXiqYs5zIha/ul5DwWDvm86s9G6ikXm5U+RK5PYgqkkIEyLIrNKn
DB8dHztNQMnufVw2OmaJJTOagrhppzNJ3ck0/0ea72rQwSNR6+SPk4nSPd+jiJfz7aJYKYnQZppC
tpBMKCqNsNz5bALPVVdBohSt6bl0xpKVR6lKJg7bqFXHoD9+Sk8AiiWASfFWyivbqdvAr7S/5xIG
rq8jjBnDCwfbfo54q4Hdwpk+/vFhIwsMzrSxmxKcviSnYra5hLCpZFMwD5gMKU4QTywwSzPh9DI4
zdUnH+abPECf1iBofh2inY0mImddgkxQegQPt5m7850zwrU9En7eZ/uUZqHnae9gdCPnL9luHQ0P
1xLAZk1JLLT0sSNPQs2+KuVdBAkf4VAKvXoB8eVDkbQh1ZMwUANdPgVc8Iw3ep9i8muST5dUFDto
iEWyQFmsIhYHIYqtOg2+pBPjdsVjBvuVk5RA3dgMVCzHOpH0QlDsOyLKPQ9dco2ylG6K1y/4M4G+
1+b5uQfN2o3B3rS0IVONZtPiICp7MXX6fkgsVTiWLw9D0hWnrDB92EQSUXKuiQ6e3M3GDo1yparq
09oMxX56grdD1Wfhp+XQdILgrAIXgnzs7+kEOuSQJlxa3OhSLgMer6B9QuwGJ33djgcRTcNVQXvV
JH/i89d8IHhdJ+ZzCnBY4nYEJZnBmxc/ttr3OcimsDPsx7y9rwnXPr+EeBVLzk4NpTzpwO9T1Jhc
xtpXh/tWf1twpuffW+d/x86FgZmimzqtD6RQ9YgwZ/pbxOknTAU8b9X6xvngdG//qPWuR3MRxMm3
MUS5jOcjtSSnBU9Y09KfKBjkfCaeTHX1yv3wyGoVc6guEYmsy/uZyjsvBogE2iqZMHHavhWNKSat
hQVcv7GGJiDvoJngaD2L6zn4QqJnAYQlinbBMWa1qUTzUm6THexGiltINpUgVg3+AKoCmhPmyfMV
zPOHawltwj7O9tzFYBfVf0BAcxT7K41ZJlwVibYhfj7Qp0GyOSoMmoTFofxGZmcWnAqKKqGa8gfX
oaO8WOetftDf9Fe5CRAsxJIqDgmL14uwknPyM5lyAhq1W7sfMEbGj5YsSjwDdQvvVhkxapDG/wLw
l92OhJHx+HgcMwOjBHf/pOMqCoCO4OasS2lw4r4TYEDwOMXxBltCRnGxXHknIrq4rboDTnDvjEWp
wwEJAWP9ee1RjiEWJkMNFFEf2vp/8x7juBMkDmPqh+1AIwKKPeoGrHp+/KSTtbfZj+VbTUqGfIG2
br/TwoRtm6RbJepYAFHp2SPJMZPUF3Z4+yvOAupI3vXgz4+zzcMpc83uoDgii1yv3eoWB17y9EjU
j4zhNmID34MToxYhhgrx2FcdqYO1zkamP1ibUtFO1sCRPZ8dZUXzh7KLNxdKdU6bp672JMWHG/n4
gCgQq98rJNMnRSCmNOjWGYK5uH7em6EVPppMDXai3Zz1CrTB2jCy3QCAXwi33AKtdFEz6dLU6/w6
4ZVBjj8ncq8dUyh8uK2GMPSUMct05mpOrQIjohXfJyC/+HxIyicWfKvA7qQ8seriwQNtuBvKjIdn
9cN8UY6PiqU3ITucrEQTnXmj9cKMDIT5ZroyoBby7n6pI1udMn+wrVn6EQS2tlsm8JSp2yslYrJA
atsFrpSAoA78Pi7qW8o/3+U0TM9WYrlK6ALOmrfzhysW5G+6eFMULaWGWg9lYw/iSZDlx6hYU8mr
cFsJji8qkzv5M++L+x7Vrb+0sBPdoRAcUPLHHZ+LrkIlXnVCu2q/dpxxDhbYiMx8baDrZHmWG6R5
fW/Nl+LR6jaJ6hXj0c0ugRb+A5k2imEL8VX7TxPc/7RtWgoeaN+RN3fxmblBD/X59O4ZXuKof9O0
09E3Zgm1c/fott8r4U2fv+C4tKNL8fycOuBcqZ0wXe1VX730gBkxVlthprOfQj+6Br2WM8DhdRq0
4pv/dB4oedUZFjSWbNx0EVZMzjglkbwNUN/sTMw9X9tV9xLsbXP1t8MQ3zmhSh8Ynb2PCUUwJk6p
wNgmevikn9kOw1oYpKUeL2QG6TsyQfPARZiH7QBzNvNuWbFqATQiq0aSue9JWWq+S5UYuZp6mvkE
p0FU/mPBL5k+aBJXxU2XfIucZoJpIrnc8gepRMgUDzkKIGSp+xnLXrWdG3lNiMsoJWUa9IFOoID4
IaPN4B3YA01SHAgZialS1rsTGbDPmJ9ZSlOnnvvdBtBOw0onkp9f04VU0z5khiRFh91qDal8a24s
QrWU832h/e/5StPXv5vHJLVVz0AhHpPzvMFnBi1ncbbjh1ioE/Cm0N64ep9zZLIM4b9OGSx0JA6F
2pMMq3xc1vtEJKMemVeliJ8Q54npoz1B+BCY0RCOJ/BwtQSobvfhX3whBptLxohiVKpzYcyTWaMN
IwZyPoMt9DVdSpdkRlLvQHrfPA56+rTCdif3GQV9VYliRNLY17BS9h13bLpRA5ZE2ifte28hGf4M
eqUcf0CspV8V+I3sKg4gtf3FJYmzqtHQOtriTGpHkrKXQ9fGxqMHxCJFYCOk8hrZvNt7y7ZAsI+C
d9niEWrnHHVMUwLWcS0UdtsnjnkIbfttL6gjz/uNDP7raveTlGa60o0sDdcYvgq21UF8PWw2PyCO
GJHnDCieU+lkNU0mUnLfYQ685YzWBVFsd6H3d70zc/7upuBMZBfXb20wH4D1ebDmpR3sm+9FP7Lh
98+O6JYLRrXHCGz9pp3E2SAXl9PRj3nLhDC9Ji5qnqzZyCXEhGseZ9+SO9xHZPrzbEveKTfN/YXV
PmZFwcmkZSx+5wBRneq7BL1Tm9GyCx1x1+IYzTgzvP5VYO7o2qRyPQfFJ0azDzdBi6l/p4G3iHxT
sVprowy6rsWRHHtA+6K1lEYMkKoXDdHaHXugRIw2ksM14XNO9BFzAwVG6glkxlDuJthRf6eZR8J8
V8mi2gHeUICxfGnSx3X/QzbZMd6iR4kyYwNH2BWNyZ9F+oINu8oRIJiMlceLhr9kIlOBHG++qaVb
zX7qnC3dIH+Hy/R2BHGePBaEJ7j1E0XK+b7RRagZAv7tWZhrQMEjPYiV4bRQTpsCmP4nZ885mWVk
lOX1gsPUzPWgT1iNtw98xpoPi2mDH4qqkS43lrB1tyjQgOol03sI2uJ2Ma0Rp9u42VTqLIb1CNjm
Rp/ZGJPr0GHg72+D8v3KcTBMLACVRkfSVQI2/Ey/PYCBQQZF24MMLsEIWZKvm9ao813Px6QSh73w
H3qnHACmVYouVohTwU8YIHx1ROlTe+45NwgWCE9OGfRDeQmzXfuUp9R6odVK4LmwBtDJzIGyy9P1
zLWsrlQXxeaVRCI6a7PDWuqgmz9UN6nNlZjp7BdiYDiVISY0s0ywQ1t9NMYS3ni90BUB9kS6nCqA
hEFwjzplavNm+beQ6Xbh78E1PqjgDv2pj+ov6+THAnLqt1DVPGx3E8XdoVXlDQp8KoeJGugcsNOQ
m5B1w6Kkgk+cfdjijASnVM7WQTTODHZ+HDkb0JYk+NwXO9/Un/qZhHXX30c+NMJFjEQfRGVwuRai
teqUGOuUKMig4o8AHeqCdLTraQO3Dwm/XRl5iPbslDbM1CvsA6zOZSQTbeH1RnEyHpe+tFLXyG+F
rj9JiuKkThUSt6en6Lbdcy0jueF6UPkUBcLIkWKdwxVJD/h1KIYjAHp6riLW035zudVelROYxuS7
abA1zk61vmDmm8tWCpXyC9a24ukND9aFqkqvJxyTSMEHak+KQdA1PaLTCICs9+cukYmnNB683MEh
28/4jwlyLvl9h2DbghOgHOsqr3s81sED/x5nzAR2tyvUDxCmJqxs0I3ywCF9RBz5ElU2z1RPN0ON
uQO0kG3YzxUH9sye5LEvvZThk+/w6fu8JxikCGa2GKzR79YPbvo0wV/fGuEmn7RSFJS3a2xG4RWT
h6l5UuZRk2tZCLgwiRzCF8DCOe0GKq7EaH7Q+ynRhf5Wfvm6FcQ8utJkWswlLSHdttoiyQpf0rtF
RUukV+IROkh3or0faeB/pylkqwfn542iLuB3ZgEYOyvPzxXojlA+i1a+wK68qg7t0psGsSzTiICz
WXe1V2Oyo4MFAdD1McEk0GCLYHgrKzFc8Mz4Dzl8Hf0uSqK9JT1/ivYkJTEGU3ldyY2jF0JQtJTr
XF/zfzeTQAMeh7AvtyQfUr8Qukes53uRpmEXObH91bCfrK9iSOl4b2q4AJyfKz6aZz3HJEBYqwY4
gjjNgKlV947tVO1YNwHdW3dmP9LieIuYi3v6I+6uAxinyemDA4+TrfIDoFCllNM5DQRnnbLlJk1C
ura7MHwQlTmx0714GERmw0/tV+0TVSdywAovAGe0eheTqgnGORdhDEKoS89GXF1XCFMtKUrrB41L
xJarLA8VZzldh8/iIIdoz3wJy9CtBn3L+h5jYIDQTM9ReAB6zMZZm1dRteWagERo0zyu2ev2a0Ht
Mz9YhG/nIBrY2EnFuEWI3s+QGJ0Zy82ZuzJcwbt2yUDUtas+f+gaSeZ2gJQmgLWvWa6IEJlxJoJP
+8yk1ldoy9uAaD1S+BInKdWtIiMyQrzaWtErcNEhk9/dhNZ2fkjUzeMMVp7JqB4yiZnxuhX7BJWS
uxuRI4YMYITQhRrcowVAWDR1sQGM0gM8DLFFmKlus7hvdV6DbkjW+HSleq3SeEN/TEHo5eo6pMGD
y3FrbyI7W1Tqri4xVOTdn7GZQReWsWWLAPsb2dxiwJI8LbMFVHGb6Y+BCh01BoHjcBDrIbAZFH8X
SyDxnqRwJlCEeJ2Acv3Q7Wr8Cq7JR9lbSGpswZmAQEDKVxb3O0yxH36Da3enk5YWAhMywPqx3Oc5
LJMvIU6RDzJLu2neQ+lgAAODnr3a5L357It/UO95QNMEDlRuETvP9n27NpwTxRpim6aWNv/3zflH
Il9VrHFScew39q7AVjYA1DkyrmNiGq2p6NFagKHD/yTKr1z1fPv/KHl3SsJ4mgbiHv6dLDhAfNY5
8QQLs/OOC+lROBhhzjbAUwRKRWYIdkfe6nMI2utwiJzfrujHhGaXNiys1VO0cwO5vDeY+N7YaNa2
YwSBc8EYQMYVuUYp37kogLYvKyHCFYs0XRoF1jzSTOTTL6Ct0ow7R28Ipt1jHR3e0Dn3Nnx5+J39
X3LUQoh+4a6lECMQrW1xO9iudgoZs9nBQxHLbFuNydEJmdeROFIm9RFkoLSNO5d6lef9pCNU0Vfo
n2W/XNPeZYZqKgwpH7qBCrgScrIscI7qL3zxnpDrHaGNUqhyvtkr4Zq42wQUs/bBPGeTi7sKs/2S
0uGz9jElqaWkzmj7xMB3dTqjPYnzcR9G0ZY38RSm3W6SabFNsSpta1OAE4rCVFnmE4CBRmK27A5T
/WWaiEJRQ2k0eS0SQzH5mQOo+Vgg/gQ/jxcwD/AivEumPYZp32Ubijc4dl6feGiWMbWsUyJ/CNL6
+4JJTDiBItciJm+M81NHLYPcQmPiVZgAjGwwcLWtHmrnuMOK+fILSESVY4tkvVu09GRzwCy3hP3U
p2SJhLtTGEoOXkNlclcvSyRbGk8AtQWjcK16EoJCLdFDq3PNPBj9LME82/vnxJB+wi/qqA2Ehs7X
T632TeTCmKQNVye+Q2i0bQUPRZ5mMiv2hIdveYa7JMQbF/j2MKWIn0D3eQ4TIBpkVbBnCTlDK/HW
QphnesthnkbPJ4wilIG3iOaLHHGzvw9LzEs+QVrz0pmHuZfnPS/vP+tml4DzZTGCSac5gVtRG/iH
zzJvxayA5ZADgKY22kfLSPSpyQkSc1YFpXm7eh3HaQFB91kPf0iZ4TppK/XHXXw1tUpIYiOsqtiX
7I8mhsOy/+vZPYdagkjxm8Yh+DjP1GTe6Cb/yQSHMftyio5RCa2dGRFPlmKEPK1urPgHNDDNK9nj
Qy5JJYMw47IS5TLfeZTwcFwL4hy4Tv1/QVETrdNH3nbeQ+Dd3ceEEXareAjLRzTMN3t4I3Tw3JJH
VU9WjVsY7XzITf9UZTQfRWRtpabT1UDiwGvodzFyYCnNGHebFWmECxRrFCAE5Ce7JqhwFcfDyg0a
7a1h2Kdl8xYg9/2JX9ooKa7zJ98Ynwlr7+C69Msru4fzFMbB4pAFyHzRZ25x5q3rB7iCPJlcR4NJ
Gi5UuUJ3iZ8k7+NuWBNUbkQiV/PTUCH38ztV3q32s28UuD0xxzDoDF+n4tQ0GQ1iskVH6Dk+bI81
iK/+vSiFaRdIDgHiqFY8YYR/IdTUcNuRFl17xWMzRP1RZRlkpqplJvmKiwmGrJ8YPNkNyR2obOiX
NjcA5pMAfVWxNkFSYDwSKR0UbuliRmP+1t+RALjUiXwpCtQFLsQ3W3ZzTnAiVLgUg+tza8rAImF3
fxq5oEht4PuRD1R9aRkzlmbPd3K1wL+YBl45f5R5cwXuTHay6blHJoReKlNBlzBjISWWUAJMRdgN
HGP/+v4SeSa3Vy4H5APTM6hEWNLbs6SvJ7vqCrQ94GtS1kOUIvC7KyK1A1msi2EzberqBk2XFg8Q
p4SV0CR868E2DlbgPFJ1AQyTqw8ZEFeSqcMe5n7MjCPmLtVFFiAOzEajt0ESKBx29LLQIxYMR6OR
aqLndWKX4hsLs4g0TqLaP1DSCIQgCedP/NizCC8pX3QptEsgJD3TTf1AaBz+Ea3E7KUPS/qZNbYt
f7Ld6nSSnGA/oWEkDzOoppx8x+5F/J6w7YJ4loiAiz8GsTeF9iHGnz+DvETxIezRTck0Gs+yUmon
CV7E8a+txxKhq24RGhFxT/V2OovfSHoiG+kuOJRlesxTCGifQrvq8tkqUSgnqILhKzRzcI0B1ELk
oxLYL9/3zM9kUF5YZOQszXHMe8CaxDXbYb+nAYT7DQfX4pJQRrRAaT8RGBSHONIgwhUwLpXE/6fH
NLNYgVATs+6U8mPu6QZx+K4dZ63/pR8b7rFkPYeABY296nvAMPu5GA2m2if1T7XrG4H0yjGGfYU2
4+vWdun5GMC1uQ3ezYT/A6AGSlJJrz94rPu0kjGoad64VO57RukDEtHrZW/+k8y42fQIHGelr46p
nVz3Cn+tPf9lc/ylnBLq7zXmsXn86lHmPwdsDNDMPDY0n8aFJe9vZW2cVrbE4fc6awO7kZPL6m+o
36g/eBrHidvRcU9l9CkyzxMW7aQFc31IaUCNyeRnetcKOcLWgTfDqpdA+Cs9m+zbBSwDADkLGzp4
2qMCPT2e9+Vhp99suq1Ie2Fxyml4L4lTxtCD1Dx3ozV+2H9M15HTE4/3L1RucdbydX5gohlWvnzk
ZsjwXuEiv23+smQxVj4S87oXETEH/uOCFNv9KzxuJUMd/edq3zCa/tVMu+NwAWxca1zz7O8xrssM
tyevL00qv0mfUC1twWHOdzRVbAMM/rMvUJzwB+lNjcGM680eQmPie3fITVrtlJqfBLzKArE+YGQ2
lGtU0FSb7LUR2ha/+fJfg2//ctchk72MBIwVYLP8vUz3Rxu8poWY93IDTxKqqSpI3Ru6WEv5YCoc
/xhRaWstS2FCXveWdMVz2klhA7N9zOCb36TxY0ksNFM6YYwQqBj6yRUFFprGyve1+O1x/clEr7ku
kQJAQMk2WzcVIwZwa/NIs6MxXfDFtXO7fQzbeOVV5MdaiMYQHC+AdbZvMPgRzJFWJvLq7xJ74cRm
PdXaC9x2qcwSsE0Mv/1IQoMMzgiiujc3tbPae14hlVx1xfGsRxJDdQKAbUl94IJ5W84fnuTNmKMY
G5nqJkOQzkRVzB+gnhLPgLYzbTGNl4+1/dTtTbY/YPf62kbsFxpIMf6V3uGTh8yuzzXY4zl9eOcx
kKPkPuWduc3Fi53w7jJtkjtwZqlUXBJNIqCKOSBQE6QBWL7I5NHj5EEsWKCHMHeEDRf26MCHEw3r
fIWMmeCSVV1i5l5/eSxisOGjw5JJQ6i0A5L1BJxHgP/43sMEL11hnUFwNuzevO1ZoqbR5i+IlIvg
R1YQA7P8LVgGlgRWFcQxRQVjkF4f8SY32lfg4fLca2/LpghioyHN+Mmwi0JwwsNxgxwzguuJq9HO
LV3WEUCoAwnAiPpA2ZeJjWeFtqRQP97w5+Csl7K1vp6+sEonuIUU+AAZnQZ+6EPwyh9xGoVte0Vm
3bkN1DCUBF3D7tzpjwg7dwN7ctUR2AqAAMhNIWvJfCvLQBj0Sz9ErekWVbEIMUlLK69iExakhHso
b3X5Tq96sfPk2TnS4nUTqMRXoCBlSvVkEJl/YRxGiYCTpKna1NVicapFdxXZ/bj6lUVqMckMCtMg
WOrr9C3FOoQpohkjB+lz5ejzcv/xXlwA3PRLPy9TOPROPqOhl3/xaOzX2wAW6CmkiCuhdi/V2dpf
I8eopKdr2O0qVnKDEAN1gkf3VvDUKpLkhSOoPaXKQdr3zfyMFLJliySI103iogf/TcgcKUFyc2xx
ROI6uakw2pE6QEg/uj9Yg234Ki9a0GZUonSh823y/LtXGegeLRwBFQnPWPuudUOhJq0p85Lt+6Ct
+aUW0Hf4tvP5w3NZl2aC+p/AT7YdHAhdshnnmz125qHTqOjtLPJSxGc6SqP5OC/D/ybW0HoPD5NH
TayZUnoLDtOq9Kov39JjT4lDzF6RcnCo2egLUlp3vBBFl+ehtbaCSqgjTeRiLlyT4CobqhPikcph
EYbhD0neVAu3dky+Y2Bg+b7sD4sMW7T8jtycvxzYT6LuYy8RJjx8nD/BwgrH7PjuZpahIYhGRFe3
cOGpXI0fcbeMbNyzKp8yK6niJ3B0VX5ldWSNGWLPL9BrlsqpNr41O+0VR2BoktgzvgJIr5tphRjR
vMxixYmozHpuaVSinYR3oc1z+tRQaM/ztH2L2K394JIry1nS3ISCNxcvXw+fqw5WAP1mcGjIIRC1
mjwjm/9GxR9Cf4Nk1fxWWVo8u8yEYs9uBEUDEh4IODxh1d1Xvq3267kjzHKg2SRTSmlqeWrWhJgc
agBPrY9tYbCXvx9jAjdd4ZGJmtbd3rbCDP2LpPGQdwiY6Y+beHkD6n6MhXCNuv/x1C83mkp+9+pE
+zWMroPCH8D5isHS5Rr4x6AIPe3grsJkFdiESgtRfbl94vaufrRMuunNR1VIenVtvaRndBoxzpQm
DjmkV48Wn8oMSmGCV9wbtnIBWfLe6yBwkxmQqaNmfirkV3ywGMBepNgg0wqGi938MqTvdMyzBsI/
FdYOBRu9Wzz8g+lts8YLtm/D3fQLhCujNkWjMUSIFKY09Dowu9+oi+J70Ji6s6JcWBCV7UbkDYzm
WtB4iaTvIwMNwU851xjpf1XRxiMPnXQXpDaeipmMeWO0t7G1IFjXG+XOVzWj2hzZv5KbLpu4R9sh
GaCqp8AFM4HAYH6gdP2HNWLoaMU8AzLsxrcPY0HyuFxlLjOWG3fdwd4XDQ2mMnkU2PafOqNKGuEb
uSKtbyBjgGPhv8otHiNVU8y+EwM1cRGaXSBsnnQ0RlO8g8Mx+vqa0/ErNtC/THqHUSUoIPNLfRQY
78LmtyoL90pxKpLOxbVA86m2rDqxI0Hhe60o/nq379sNMUz/d8vaQ9HoclgDxRKPYiRWA+ekriuF
MnP36pFRLFnwv7DAe6piMLGNuR8/qVPgb+45cghbmT37vj0O50f1Rk5Myc7Kptq0fmGC9pc2fGK1
k3S1gl84HYC2rXmrP6Oqx+TlcyEWMg/ppLFxwA1qZy2AKODhZTCFYBVOZ0cNgYbdJ714KHk4yzLo
E69yL48DYigQOsXfzWshgiHwWq6tKf8w8CUdQJwqyhLswPOlGJIrj/LA4L0pm4BOxj1G5UU26CtM
UraReT+CUMYDe8filQM6ZxhaorlLYLB+Cl4UcxaIG5xrJAAzBKV0h5HRUaUEjs6IlUN1ejc/306n
QRF1eTfNtOpKTUfBuwDaxSfMAG2/aL0Mm/MKl41oFWxwzJ42V8l/VGeGC5/CqiTu9NGRYug6qTS7
9nC5oSg7Vstl2EaGmpKUuYYzqmc0XN7Uey5zYcxaUf4neG4oK6HPFQVM5oSW1/LTTFho2Uu9cB4L
Lrw1CewOJ42DN9gCqLJDBmZgISu4SAKEJCcQrAyV2Pzc0xuqyJOufXP519w0vHNGU9oziCI4PBa4
1W2JeWqk8lSySZ6DCpWRyPUXTtolijbfd841tkZWFQrWOJi+hWQHo8otJLUAeItgVBvPYpN2dhNH
pcTFIJgoCMP9/aUiMy5Ip/aGyRGAp4NJdNbOg68lhm894dzLJK/N24HfUQTQdSRxXKhv2LeoEuQb
rQYVrAoHV60rxO6/cS0pJWQYqdN9elJA1cViI7COKa+AkELA0lmrl7d67XyRKHfN7X3LBtNJcr9V
jeD5h6J/uMps9EiKzsNyHPhATP+E7uf9Zuo1r43eht80LyW23MB0JOAcxVCrEKPUB1EjTZt14QEl
Zs9BAuxMkqT9x3LFFvf0eXVDB5SYiVjzwIiTaKBXSM+RDhQpaS/e4mL5kKC4c8p+NyImNgMQ9X1z
LbiqX2vO0IpMVIzR/C91HMnrqU2NxUam5zNPP4YZeFNZmslcHAD1QDWUMmfyUN0h9OrNplxc9Fqf
COWXjN6yRxa0Y+xVyhEVhVYhWhlB7wwWrm5BezvRd+oO+W7w57lf7m6iHlqVWkq2OgeN9SvmTqA6
25TtAv7Q8BLZ9ff5JbS0erNMm+GuUX54lJ1RTQn0/4FiBd7fM1i2ffEbSRWbYjdyUG3w3pjPqjve
Fx/LrqZYHyNzHndL3WIwv6kXCMMzaOTtSszuGxS9uLB2E1iH8KGLx4+HAqwWWtMaQMV4yCvwD+zx
TJTft2YdLpldod1egAOrjc/3I1vuOkTFuwpNfoiyHlxxpad7WyrVxhc/m8KnPmLNsQldQZcAtAfo
8HHZ0FB7CPH1mjv70tqt2nzf0VfVaghT4BbZXRlutijq+9x87cpsheHZHUlzGD1wY3JVky72EVRu
ydSwA88g/O+IPjQUr6K0n5lss3Qnul7vaHq5vQhyIbONOKO5x/Mehm0gnNmMBUexZdedIqwnk/oU
owdfp8EjR09qFqPRLIBFC5XmL3JaGZCKeu4vo5tg15pxGMxRQJNPfsqPfpqZyysHibKjjnm8V1ca
05uHjRxVo10lRVWTnQkp3sl2kJxdcLWrRmLJX4zIDJAyKI4pjOwZpUZGgrSfpndEM4s9zxvx3mLa
og98cAjgeajJCi7x9TyFSxf5G7f9214ol2uPfddOXLIfIPqPdzs1PCROyaK3ChGFoknE/m6n+e9c
FtjqVGOvMmroMMpZm2fmXrytENQGbbDt6xryTEo6ieDCZIep1QLNu9ymv7WOjV5BFp3HRaS8kvnC
pdGTzWjx1yOtU1BciKC0BWKzDn8eKbZmVa4Dpc+gxC3F39NYhnr1LnmKfuKuhGQ1NfE49No87/Nx
p6Ek1PDaXQEGZHQr9N7QgEh5BQwThpttpyvpfNE5d19UsvdPZeGd1y+gHPNivBm6l50JXCW9OsOX
w8uBCa1kPBu4gIyqrvMmzL5r7SC8dHSxGHpCaKulEP2mgzuWoqyMo/+iDWZfPZnPHzNNUAd5Wg6C
jjsu1Bp1+wARlTSKj/96dUYiqJjnAam7HieBFYkzwGDsQXGI8SGkbb3Go19XTROWw85Y/QQwB1SD
FpH/BvlpPaybCiRCDb1cSN2IhGEKlrJkFVmkVgfVtbWJiPAw/wElTrJc9EHws2fvTawINEgsq2Rj
DXMfFrNvFRIzd4k5SX7uqDh6FX0MpzSbzFLgIrge1rpEDkWE33E03RBEcIQJujPLWwOjn3ny3DKl
pj99xPEbkh3ia03uWhrTT9YpgQy9FThUJH7GicuK5LHoqF8FKvg77bxg38kfAYzTvd+eVKhtOWso
EOtllIqMg8MOKf+XtdR5WRoLOny1ktqYpjIpxcN1mwX0eiCq8FN3i+TnMUpk/+/KEqNs7MuwYI+v
N3m2bOiBbmUZDaI4F5kU/hkc6eSQyiCcO9J6McAKKZdinETFP4my8fdHBm9rHax29ZodSPUWadIz
o+UU/V6OLSPqWjGVe91oQUCfX0tgU1yd1L5LIcLxHN7WjWgSuy//xQjbXFItOmRFW/Ss9XqTL7Us
UR9fGAWKMuudiDkK7J7Q4EYZzw76dC1Jx4ykZEYA9CIU5VAhInxM84iFWw6Nmi6EDT6zebd1fIhc
pfqwFFNKiX+81u5EiUXOCmIy4aXlIzbqR9zg0rSEpTpNPfcDpPJO6J8vMDQo1dPcUsO3Cnwfd4R+
gefQ1RkD9PHFL67lYguUDr06XXvcu10WaQ83JlFzHiMeSwl1yomxllyuJLAEDg3nT19ftyfqbvAf
oO9Yo6N9AGsoHPx8B9OU/vnBhtFXyVTIMLtSCPcKcQ2XmrofNn2wu8fLcDHyowQrPDUlSrcna4sw
mxp2NpGkJ4AX8wJ4eRi2b16Qx9lwyVHAW4NZnaYKGovpHXOfmv1hDH0UrzABV25Q1XmEoPe9YVEX
NcXQ8wVQ4TTGmFeiaJnrzGVBjnBEmf4sG77Qyn1iWFGlvwD8+zOhV0YzXY17OVZCoeXNIg0BGUwG
cwdsiFF6lh2BzpcYgvlhMzUWoYwnio0ha0x9ggrXBA8T+NYHsQrsnzOINHWP251nRFtgzjQTFWCb
dykV2vQANEQx27cx67+6dypVcrgXB/eqYSGNlb7LEdiKMOPh5QLQ6JVwlD3rDV+1/HMtOFginwux
k+pn/2r/tBmKieT2v3xjao+qr6q9qzNIMLr9/akWS1kvmNDEqYSq/RlqmBVnI7YQKb0JcK1uhdGe
JJptid1qLE4pQF68IDn+uocXYDBBVVroI73U7hmpgVuxhZbYwPaOIagPvtqW6hqQrGDZd3TFWDyG
Cl7+5xhBC+ssW4lbzdV8LkBJ40neX4wEndmL8aMFUyCajSTKetmIIZSo0pHEkjjgrZExQ7sn7JmJ
2Aob+hxT+0DtnGCHpfiLlg3jCYpZIEP9osQCEd7XI8R4kLERAUYH8APckBK+w1QSW+IdB2lJHweA
UfjNUh8YQ/zRtG07o4WTSRnHXBv+dx1CJyE+htM4Ex40YE0CPHl89ZG06ZEH62SU008C+uVr1YOc
lJQHhkpDrIzPTt7V4iIXoOPz7IDfGYHFCsSlI1neP2Ug/WuY5oAK9WgF49oozNIguvVLoQpI2RMS
UsP70jI50gi6GulZAsorSHMO+46Bng5rtXgkPejITnjLB8pM+Bw9ykQ0GQRdK26YqkHzoFa0TLdX
kylEPaIotepI9fux9p91VBLFAAllwIAzVse9OQX5MP6dYr3VYfFfcwkfSR9APX3jmDe+/jtx8y86
Swg+cvdV2INcwiENuqsInjoMdyZTN4ywzbUvqZdrr931wez+W5/ZSgDBQvWqHy2nBMKsihILXisx
tQj3ObZwXQL2Nv8/+BPx8hYdgYpl1nDfFSk0ieS6fKRD8/jX4IukKPehskBGxmuqrxcdnOGJwAxY
CDMcj84bf8Vz8ie9dIwcYN5/YTkhRvqg2wOSV4a9l57TlX/5A1l0EaPL4wI8IswhYh7NVn6BPMfh
6o/VCeGYGPloJssy+P2CmX0Ggt1jMIxqxKADhcQvuVpX3yBjk22yWDF+IaqzRW4N0YRa3YZKsF/I
EFJHXq4bIZMjhN3B6IscNZlxcGa1EJkyD4Jjt72zZfSHaXjHdQQTm4PBT+58ZPQYBt8ypy9WHcKK
++mFIiKbuzR4TZlGYmKyju9LnhxYTCRF25TnFXeJzLysZJQkoHAIDvSx2MWio+lIK261lTETdrPu
YngYLwAhzILwv87AENRH90qlua2673Lx/kCorpWu6nzTWC67HCpnOqZiUYQlXqhjoM+3tFs1yx5E
ru/0wgoyaSdnoZmx+5Hwil0SQWkX5BCrq2PTk6gDXbLGGHcURqws66oDdhWG9EKrsP+2kWBg334e
lgVWEQJIr1S+iHJOk6Dbub6O16AKaFeLfHkKo68hk+/PVgt+WghGxUsDR9OTm3CFdS6DhXnl35M+
e9HhxsTOJRLl8NabNFdKehDNcvQ5+3KvY9qMREjgxoKnJVy6Kvj4H/bwB53DMpCCUMHpjfKmHtRx
flnKrLW1N/stNB0tpi1VlYbe+PX/J17cY9QIx7+354i8SMdcdiNgovNdd3d7/xh9lMVnM6vBNf4q
ikNjUh8WLiym9dhlXBCufu8mSXd+A60cQt5SuQGShQcIdVySxbT76isFh+sL/+NXgo7mkHu9Skxa
Wn5UXmjt0FPMzocC5T0SrNwiC4ovOdjR9NYNoXApfkwkYp0hag60inY8fWwMPwcqTE+3xeI1n7cx
CH1s1Q/91aG95z3qUIcGOZmBvpqPf4X8BZ4zCqNqAhinEJZFtbIuXZ71nP3zooh/lCfKEjbi9aFM
VjXmL5uORSnjBodmWksG6RHK+MNjfeBqNIsfpa85x/W0AI1XWTVb3L3ehcvI06xZoT5ilQdFEzDw
idE/tm3BdJoc/UyBAHVBK2Z0oHRQj055r08Pgidw24vYfEz8yVG5TecR/JWbqVui24tXtILy8Nne
5pyquXbnElqgjCSr7ji7hWT51eSHNWMBc56GvUsJDGQJLTVhBZdTjQVk8A0D9VcxyCKxv1vMI3lQ
sKw+w4B5LvPTlwYjhXOgHrw/9vjyocvR5ePjBEgmwrZD5d3ElocdWB2ChXW0ZDJ/Gop9YKlYHCdY
Jeq63qVC9VJz+kD1wWjhWtN55/iQb/yV4H2WS08CccXEsRKTFpaUD0Wb9w2gb68Pv/RUhQhZQ25h
w6lUo5VgDko+5TAfLp/2/SujcYcJ8b/yfRf35ELD2E40pXjweyAoZd/EooCec1Uikwo72xjgv/Fd
n/V86nx72DdOLxL7Nu47C5FHxPZYoVYehrc3GG4ujFOXzK3kGyfdOjHjbu10r5zWlnHTUurL77KL
tbb70ZUNhVeqw3ZZDosM8+eCyzUenqMgxo8hdAD9dtxtJOBJoi5mn2Tj4XRfQYakus4jVI1SHJE+
qmkzj9ReolxBI729ZJFcD5rGGRcY+hiqVXbxDjA/dqYZ24SKFi/QOJB83qacxILIWZoDfSGZWrws
X6IMLJC6rwanjnJ7tFMq+lU16CSotAfTN2NKv0X6avqJ7wqbW02Sj7/aRl/MRybFbVKGRuto/9Px
cB5pVj8B0lE4hZwOVdWgOfqaawnv3Jz+Y95eBaQB2ALr0CljrOSw0+4JEwTj1oFarb8Qb6wiwFzU
8rByM4HpdSydqPQibd5G+MEPqJKQRWt+fkHPcJyRXK7JkxZ3/YlGrPBBbeJvYfwSJ5/dr/RPHMef
KsqrFNCC49e/5wZtoVJ8mrM7r5FZ88aKMHOXNHvPUEF6DfD2SNgBHzEJUcB//fUs5hZwnUSqD0ww
CcCMAerR5xrbfcD5uHyIlMPCqG2G/KCXK9U9DN53CSISUfkCMs10BiKNn5ekhUjTn5IKVJSlyXnZ
0LJlXghtVta5qiORhcPZAMIJKWo1/eI3FpKtB3VSQiUPDeLsiWqsyFJkO9RFJsF/hG7plZllDZXf
Z+ZJU+VTcSD3sbD/pzKP9k91haHxP9NLousjWF7ZxrfqCPKM9kks5Y+1qnrnhYk8CSeASf3FKVnT
PLvA6/K0vhXdO5x/PHF3w3uTJsisG5qiawPcWv7u3OKP0aAexCKFx5nmnBamWxpgBDNOQEygttkU
Gs5DIt928krfSdoyAXStutfbixF6WYki81fyaYBeU+7nLhOQxn3W/xEuv15Z1jiIfV9gDCOKq1L9
s9k5ytCvOKxtje1PYdprEzbDQ13SzPMAmRpLlfuZMa+uQAa4ouvZ3Lh4kKAogGfA6N3q11a4ulf6
m35YzIOnmrgWXNyTEBxQ94kMOIITJBUhCDkdath1fNX9yBKUFB9Xn0BBjG/obUgk2OAVzd8c54fZ
DZNHDkdhBynrYNlxfpjGbBMXoSfvnE68PedXuGpO/Fq0gBU6RjtLCmoP0TADcEfuVuo89v31LOFA
C8ncQ4QRJoeKWcSYRFSxlIJSZVMOX65uCJnto0OAUTFUiC+aqINJTm5LUX6hrqLboxpA0Q0HEhjk
vS2MMWbZ5jWnvL2WuDDGwn+Pk8RQJQkOLFcBvTmRO+fq8X7dXHQ080+WWOZnPY34Y7OsPTx4Ahe1
nWOPbMl3M7YeyZXCvDBCjrkNt57J91l4vGCSmE2jjHeT2+deI9MnObPIkS5OZX8KM1hYwPazWtI7
vfMAJPhjsMsnSuoAiO/Z3l4ThYGQPiyGxIv1od8+9tWEBsrN+1HCVbH1iOp6qMEpvlZCt0owOgTt
miZ3+kmvl2GpEvBBwnMWPeUSh7t7l041mVU5xNMgs5TRQjx75dxfJyO2jK6gl1NZbCXlXni+mky5
pSD/46k1s3z1zX6STPjYXxqG3ggB6gI76N8xlMYYl40Y4sUguN578RoQkLPH/TYnUs12PiDjjzz4
D/MfK9SJHKC+rDkCZFHaXMhjoJ3i/CnPy2/amTYdvX8eal+rT3kdvTGihwQ+zI0fW73xzdQzWdHg
1TSkpjhF6WkBCgtWnSu2h9oX2WhB0brzhnK1RkEUQ24j73hMCJ9h5M7cwwwDhnBYClsW2QiynN7N
BPULSZFfNRxCBcTYiERgiJ5mJlialr8nDIyAHUhMwIcqID7eK+JyuKu03M61LYm4qZMc/VzVJao7
/Wl4Z+d6el0dt0tUvjB8WPzugjqMODfeXhezcJCd56JguxSRTUWgLaCwiz3wJ7b1JFnhyHY9wYTd
4BGlKM0BGB56VZMWH0oFuz3WPR8mT2vU4Ju+dYXwpUPQqVR7lYxT8BuZ76B9fIk1Q4RlTpBEmQHt
C8nV6oXqt95DDD6+taidVaf3+BFdt7Wx3GY/qXA0rXRPEa9MoIslja1rOsmoYq0TO19tlgEoHvGQ
DcIumlKqkJ9OyBL+RtJuexKWe4EyCm6mzPcjzilSdAUFrCbd1f0kdHVw9tlvcuvQO8JhyMQzicoq
/jwDZ0+xJ9LSZcqDIsJjROBzVLTUe7jWO4sI3XP0eCr8OpXb9wuwDCuX69Flt1kbbyGLRyntRApY
+gAG2QnoBy37+fgnLAma+MiGOgloMVP5jW88SOHoSG2eLc07soLii+0L3YVpxp5sVtVYaD2bflms
Ow4VAHKvHsTMZFRZe2TqVWQnshJ6qH6/KvNhU2iBhmeCl9XFbbCsKa0GHWJvxmU4Ed/gBlmq2Ekk
MetOAQ0Lz0Ob/cdgor0cyT0JVxciyN9MAdg8n/EMS+V9FMiKInLdsgyOxAm7mn7PI/RdVZkIK6Lh
zJNieiF3crJdUMXp7WrrgbPCHw++4sX8YHjqFtJ3840wIkg2njb2QHwyEEM2hNDIxzTB79ZZHy7R
dd9G1QWyJza/STa8FQWOJaDZauNvWHHyEeutRd3SZQY31sN7a4rGZuT3O4N592o5erT8rdMU7QE7
oLOb6ScJoyvCWRWcp7jGWuM+uKGkrRLVnmH2Zq4DiQd02frSgpkWRwNsuSCzjwHbvS6OPuJ/dmKn
EKJYg4b5Y83UBcQJmxUdAvKvdZwUILHuXpfiqhNOoRn1GBvV9wik76Q96GNER4tuO6S3ecUdQplP
W2yzbqwKatw2yV0IduFmlGwnStIxtycPD1gM1YO/vUI7i5V6DGNRbEXK16E79G48K8YuyiPwNSvd
QIJEgp0p5mO2vFIKE71/gM0cENTaVch5PjKlRahcdxnebRecJm3bDtDbgFD+S8p0iUiopWH5cJAU
oi8QnppODNmTvCe2j5ik7NUKnTcy8xK+2XVF5mNsS2xFJuJo2fMeWGxB0YKyypGMdooJ1F1a1WtB
CdjbF3Bnrzy59GuP3z/hcHPEKE+Kb/ju0WFA6cEuiV+yRX5SVaZdbta3S87tCk0phT+/w0Zwny1P
kyVBU5L0QjD2/eCjZ7CH1jVsoHjiNgxSFoQlM/oeiSiK7kMcinHnvkUnpauJ6B++5URGp46zjgKs
yzxr4cnskDFIMc7QvnnVuObV9soH8Q/9kqqusBEloG4URPvtHxO+ARIUWUNbbNb4jjOVamaa0G7A
8KFwsb0VcmDyYFGbz8vCch6Jh0Xz1ilZIFZThXpaH0OHIbx5jTk9w4KdDlJi3zRUfGrcLK10WcRp
38TuRfLeZ8vPGxDdQZBkI4D5IY4RUTitqVq/m16x//7Hte8K4QA3Agw2QSpJBJLfFAKqcOPFOJ7E
pOBmOU1qPSr0EhGaXeGlNwuV7ld8cC69vHhMLQZxmNergbEOejzpTGiHmWcA5GIMEHuFYn9cfAqx
i8tBXFjYlp8Ggd82tWMAwgJLTwnn6780IdCUNyQFTH1nqV7CHgEe3OluBxx9bfgcn/UTTyV0Kbcg
Oi5xVuljk5ZsBYD05KHZsPIxwP8+qBfthHJ6cvNDOBrouPf7eS3NfmV68/W7/MG66EWsjT6oETLl
gSRKjJVTjshHJS4QWULVEUU68AN8njZgjpOs6VgK/XnP26EvTDedy/nAFZNzMVqPeAtw8lqGO5ER
rW2IiWqpONo0mpjOENsuDJm7OiicwG1SRgAl4/B5WSGh6o+idKjEQKbwrmIazbtlHKlNIvyDR0Ib
Brpxkq2Zlscm+WUWmOR3KzD48jm++oNehskOgADWkRpYjOqb0Yt7mzoVnin2lYc8OMvcymJ/zS7p
/SPz99mC1+whjonnJFgzU+zNh/sfx9LUILVuIdZyiGdt2kVLeDEcy23LW9o/E3FrMRpLeQE5jV74
k33kK/7g0Ha7OGcNORebsseeS9R+HgjYHBDtPWn0bs/91DY53X/gzzy11VuRaolAsjby0YRikEVa
2rbX5Uy89Bf2UjFlLpuLZe9VNpqhAnmCNQ74O3DNv4q3TXnLAaM8NKDkl809LA3Bn0zI4qc19H7/
FH8ODkzehGNsLszvEWJc2CTdx0N3WCjouwyUxzoGYYX+g2ou0eRKfXklF77ZNJMEUH6MBzW/7wiD
zOg2RxiTSTT88vhDyeBF+n6RlXy+0Qgwhc0OElF09uafggIYUboMaK7r8ck6buhmHsg4XQAzDdty
ZdEqHVm7yaLZoVClX/kL/yVtis4wyGMsAXwJGkoVU9BmaMWP5PkHg1ixC8hEuK1C+MPPiPZpsbkN
6Ob3V3cocuIBD/TfcRY8pt4XxVTtK5zq4MM6YjPfWk93Yduj7NOb1NYHMqIWhkRuEqrDMS7vRAs+
SjPeFk97YBVyyoAYfcMGDv0ZMbJB9Wab7tU0YsPTD+q06YXZGAH5S9+zoGPE1YLe1WP4KkovMu0z
mIqqoZt4do8nnN49T7Pqmu7mDswDkWczzdZ0JJqw/WW/8BBiI199BRFrmRqrD29BafC5E21BuP5l
z3eKCydpKwNxTISA9HBjL+VzkEQjrzOYcHpB0DkRNS6zrvpM92FbMTeibAMbXxm6itP8x5uDFbJx
Lam0YQUM+7dIwYoYXs+7goHp5G/G6zPjDE1YO9a/cfGV0Rh7XKoC3JskFXm89OETmp8+OsuCg8IC
IgfsaCUz5zBNtL293M8A74lvu9aLnCqiBFMo8/axKIKaaG1yxGalZUHY20Jg/hxsCLqbg2pmPLhB
Xb8BR5WPDZP1jDyIaLrsVcEpvKc3LahOjlNPjq9dU8tIYCauko4T9ldaAb2Dz95jejbEdQevdk+d
C4faBXdroK2UxFdsY2NBHV1KNTZQax956F/xZD/QF1gjHT5bghBg9tUcxchP2GwlZ+9QBZslj/+e
ikdxCrsU4VfIvtj2V7h4za99gd4VfDEEdL80BdRCvdb2/VbserDUavorTAC03IEwlVm8dW+bmadZ
truR8eMj7QnECscT3X1947cqxmlsxYGfApBdIMhtHSGzdihgMQclF2L61PirZKBBJVR5OxMDJ7WZ
vNUcUdggvOtlPfzjMVVWqHrgHvtkruI/o2ocUNhqxPV6N61zxKkmimsNCLY0atS6G/0Sr59BaLXc
09bOhNSA3kZhfoyNTI85e+Iz7SqUeOcyJvRNv5aNExrHE+ZirNh8s+tVg4/i4gyg9mKYZ/1TVlU3
jepw1RriK32tYeH2Kml7sOmgm8FOpVOmSOOqAtXzurNjYjv454dOBa+o73CA4G1LicYmqz4Xd6UA
ILFa9bU83FRdtPBEgWdTGuH/GhMXomKOhxxGw0sWxT5aoqIKp292TPoK6hrlDgSHP8LCo/QifCh9
0YrkyFYnpH03tTJjR1YD/Paq4jPN5Zl0c42shTtEfLYhGL9CMtYtCOiSAmKFZAPtDK1kjSE8tr+x
x3xR8sgt+MJ+ldq9R1K15odzugDapY5A3fvwXn9SkWDo4VYoI96jHbJmRX2bVdbUtGu6V0M5bEu7
OaAMyMVX3TDtqLsZKYz/l/4el4I8LlkDPPSvUabou1DRSGO7pQCQxK+dzI2zLFCaZsnHE+z9vMhO
D5tA/PZHVVxJ0w+/juKjN4BXTB6p6j4t8uoHLKF5Bkx3h19rENLZXi7OyONsnm4Z+jy1K6TPPjnQ
7rTrJlF8gU0NrXzBGLHSSkGjwKslrWjqm6atgHFVlRHt9U8Y1vkLTwGJ0ZffyK/vKHfeBGUwj6Tm
0AP3N8v3JCNKqEeAJLsnF3s5WowGB+NoOKy3HS9yRZYIEQ1m8LZIFFUkWDGiQiAKEIevKyfOi86e
xnZiggK+iP4lQ9e9HbNY9RgkdCmYBGcjiiph04NQTJBIfKtA2BTVg80HRrxvDre7GNoEteBT+LkU
rciXv5xMstnyc+o4WhhTgPHVweShE4jZhqCfnKGqcYJgt9ItDzDZbvXOVnYTjaZX/VFnVaXYlXEE
XpWad9PHIsNaEgv5ZwnISj0wQfGw+5Am0d1AxTx7ckmkhr5LKAhF04mvHMRqG06PM5AH1yLL3jR/
ZTGwIw+KAFOsJXRUInRP/B4MyCJOI74oHC8kQDrpWGigljmgegNXKK0aiWqHBsXaFXimPFWY6eTI
7zgvYrO0RBQKa92wEcxw7KhyhVDzQhw07CQCTpm+vKSsKkgXl4GsnP1Yg79W7o2wbbnPCdzJOSpz
n78+uPSLSRPPrTCI0otWPQ7ROsSWj4yZfp4jpDCCGUc9otc+e8O8cvMg+ZUVO4uWt/Uznw1RTeSY
rZ6RaSYaRgXXNjZ7FQpj6Ftp8+0NYmrV+xipo3s/yNZsbpnqgx+u0h6Y60XJ8R/9p8V6jLVxKBIV
3VTQGM30RlQ/oVDmfH6UeKOYC42MiVsA/BKx6IvYasvHJ9bfBTlLTw46b86F7uMYGh4Fbw2dXN/A
j3aThL40MsJB9JQlkJTT4vLRkR/SO7ymfeW/x5LiqOGmu3yJ2pMq/Qwy2bCsFkHn7VXLI1PX+XMm
EcKLsp0wIs7w6C185Uj44FkA562HTHodnFQhBdFyUzg0NpLGrtehzdxAATu9peoQUsGL9W9JDTUo
Fw3oaadN1qku0A9TtxAddhV0MkQ9wAiq6lEXFLaqPK0H6ywnhcsSHK32hSdCIDdZmFtFvsm+F0/8
snlvHXjlOlpEVnfuc1qyjzw2/D4osDeINjHUrJdevZl4gQYV/Wj+xxf7i0oOFfQbIAKUxYUoz0ur
0Kdgfsx+FCtxR3fB0BZRj9BLuMqb1+lUkMFoXfcjLjD0gwUpeD9q8oMRG9VNY001iPW02JE8pzPx
sSGX+LLHLP58PpH/LbZm2tlufQ0CdedN7FXqHdKmefefC3bc57tQKutwApGMnCkr2HN7oeNuGDag
2DLQ1z7dnNjP1J34HGFl5+EPZrcpalatRRtoGnR0E5pYBLZkc/8WeEvqLopIYPozoxhvFLc8gjG5
oecR3lL7pVBkzWdC0IE5yue+yk2kRHqdAtewPRVUKPTrST46zkm+klOxwaT6Ecyh3vcbdCaiUGVK
fJyZIsF7tikehLdVeGyoYGV4r6QQslmtmo6fPXzjB9Sq5pNtyhoB/sw55bKdZVHfL84sOsi4SXxU
0Gue+LtE0fYsu9QEH0tU9EJEHPtnCf8bZZWRyAL9cNwzCMDh5YXYK4dJbC9ztgskrRHoVz7hlfZj
N1Kk4vFXR4vcV97bAEafuC296nXfnPM8Jet82HDpCr4oNoAB5M1Ls/6QtydxfoFoAA9NCFidqxrU
/I+Qph7qL67X4Fr147SOIGikoALgjDqlMFacnync2a2KQ6eUpAbuoBRwJlYBbvz8vHP4J/Cct9PV
iWx+xdI/Qc5WKZun3LwOnG2RdPwBIj0ZUN05tarUgISRSMaT2w3xKzsMJvdDWUu2HAr+5ZmQuMup
QgwRbdQcdJECrKz5emLD5QK6DG1JysDzy1gyY9vxP+DmWUuroyhYEax6+lulRU+T1VRWTLh4VSG3
wF6geuSixaL01HkBziiUd1ahPsdStUuA9jARtU8ZCsEor2630NQoSi43V19T/2lNsIlG9x7w4Cze
zfPOz+AfCIEQvmy6LeI1YztYDs1+77n619R1+UKzpyZsb2K6GnOseX8+jA/AII+Kh8n1qiqXqHys
Th2YBvZQbfawmuC3CfKfDUqzLB/tEUJtQEWyhX5GavrGL8FJw5AdG42NXcOboMwp/LCquF7dOVMU
N3w7rbqbM7c6pdGsozx486062Q4V4sO33jsTrDLeTyZ2ne2mBBwqgi2S6ntusq/aHee72gq4ryKk
8ElehasiEq/KhHqSP9Rl5z0k+3Eb/sTarYaEPqBz/JIhI3cjJ3RNn3QBI2qITRc0c3jlT21FohD7
GLiOocLq627qjKdS538WQH0KVl0eHGLFjDPse3qmE8lt0aECJvJT/iEBYhtg6v0BM/aIma5M7YaB
9XiHvApmYHl/G4ZjMS2BkFDbafMb1MnEoIC1cS1sfXifemTrcwZo84gm6DB4lMPib9qe66xOWdM4
paErDdAoxZBpoerPltHJ29WZ2CKU6vAyRrdMfC3ncH2AXw+p0Wojxxu1yMSc1vSzV/BsNi5GwiEJ
Bos8rCtjP9bT6ZsHvsZpSyHCCoIheZXBwC2WAXDowMMw5FKYAWTrnzrnhhMcfGmsuqlfDAblQ1jT
OQTlt+vlsiRYls06QFNdy0mkzAS2MYTFgoHTwogJdMpaOt8QNRx7qByerkCV2iufmTGBY5xcwJj1
rh9MQmHhtS3S1K93hUdacDFRGQZEK+2CaPUqTuy9LUL4EnXAGv4WnWtPK+w4EUbw5VEDH7s75SAb
kSeN3tmikt4Pw7qQhTvw4yh0GfAup9X6FNXhdhj/pI04byOPFM+gy+JM4U6akmJlawylQu/8Q6zA
8bXPXqq0q7UNsTPtsbw4pb8/AwWp0VhC15+S3mlaeoPPWkQ/WFSrFYgzxYqX1cL39tMt375U/lio
+ot59rPI/8fH9s4auvNiJzrc21ZpaxOxFAq8fhMLg/9XlreyVDZgbaACz+4gcOBImBkRMOba8k92
YcGIeXbH+dCA+OCbTRwqwGtNRWkaw7G2GWpPwr4kAP9paJb5njd2yCBtfT7kFFstPQnOTCPIgcHi
4Q2jcywmeiY9E3t9Fq9+/bvU75z7AXGgL4Hqw0+1djkt7ZBqd/jnNPQlW1y5/AIcgdHl3McpZhSa
mLf8Xe7o/ovRNamyZSPykRAogWOKMBFCn4k85qa+xAA3Z8PYhP0tT6Tqq3e/fHRUf6jemI68JPYc
DIds+vrzTuEoGr9GGTEUcIiiGsUIt9mhYS7uFC+HJT2uArdv0CRGkPSU62hE7ODE+Yw6PeNDlNfb
lCh76pBkLhqYX42Hfc34R94Z0ATnjmvFY24+g7ObeKPrwRHYc1gKHHlT6SCITOdEs0y+Y0CrXRBs
ZhpX6wPQO91xq6CdjLD4+n56EyfljkfqiibiVtSdBnnV8/dfArUvmZNmNHXMGdJ3ShcfFaWeqA5Z
tooKWw0RxW/J9p5a1ZFR/tlb3CdZZusxZ3UsZ3FeAdSbbkog3a6ifxBbQdcNvENHfCtn8cw+BJZh
KnPpQPEHqXbk9+mXb9AJifNkwo7P/aZ+eWXuQfSeOarsBl1bDr0xw96GgkjKDfBHdvb1NxArnhzJ
ykHCnpMBD+YDhAWoHu6EexUFOhrooeaVs+Wc5p2g1CPI6iFh3gjDMZ9hl5EBOlFOmG5BDJe66YO2
/W8pa/1ORkk+CNPdiXRwEgb7Hh/VfZqaGgzc6UoBjuaSddODYMAUhvRJt3AnaOIZYGA4E+5vGZO3
uVZoDoTsX/RGFep/LNRYGXgxZcUfkFpbmdpyUA3cpk0fuxSF6cwiJzgPP/mE9/Iip6KbJMl/Kei0
mMy7uVkTCCK1V/25y6UJw5257WqC7qZ+Pcg2VUEL1yvJR5+olxpBwqlbKEIfkTNzwilNeHZiyCEk
YPCo3lF2j56ocF3g0pKw2vuiMMCxolcHksKHgQJ45OCUj4s3abQLqN7Dxq0YrkIiroEae4hHbWpe
zdlujapVaanR416J6NaKwwUmWbt13EcVRo7Hrn2Bb6Tq4KMWx2DylsIU6MbBPKiqTgS7/tG2YNYX
IjCS3s1UUXui9pUSKZzVCM9Fv1x4jIW6tPcHnsG7LZO+F2yAbKxos8woPCH/bWvOCelMxR64Tf0O
MouG96TVty/yXRewc5jdKEIS96EqBIblm8psMSazGMEPpZAQ1T6+QHUGPZbu6e/zgHCqLdXWLFH+
wSR6Fn0+eFVIG498hqJe5Xzqv7PdVgq2rNFZtzeUVfPDY6/7E+WLa/C/V8Mws3H9Cyn1pk459aVV
tISJa8tkpeCWw2Y/oXaTwVMw71ZmgSItvZSzgzx9Hbs72xip1IlRsbo1SjRg9RoW1a4K0zFpEaa2
bd8vVqQqjN1YNJH9AzfXRxEGZYVul2sH9ZKtYrAZifV/sccYat11E9SlF4P11milwY4W3YdWl1om
E99avBgzvtuWoZZviKwj/9Zb+WT/h/Hx7Uul9bg9aiVPjqLWNtnM/61jQYI/qbW/2sVt7CnhPeu5
Bn6ysKCAx2Miv5/1+IVrbjhX0NrjUG4OD8s4UQcZCEAjig31UjXvp4XrIs2Qg+5mTD9Cle1ICZUv
Ah4MQ6bp36E4+tH67cpB/pqnVYyp8IXIlM6lsJdG6zEbbnGen8rDSu31DhTup/EiAAyZKy0N7DEb
mun3i8OnZ3JTg8oNMXbFKSoGna6WakkGyRPXIAkhtwf1BClUU1y2lTb2Pkn/19BKtYOoU7/kQf4f
fYneUrC5lMPE3fW7qUTm12aKRlINB4uroru9Q9NddxjrCRbjHIdMEfR3qvaDgUxzU0SsqZniWWuO
YnvZNg32NKaV2paJhhtjc6vEPEb6I5LqJvXc8JUN27eYmRRaHxj3RXdJJ+MYkdBlpIjiQ5vQqAme
6UHET2ZblA6basPR4wfCaTX1jqtCCEEpQGwQvGcF/1hH8v0fFxlpYgV+EtAumOl16ZVWRzKUNqaD
ne8lTcauyW2vWn6POzk9Cu7yfP1iaQtUy+Jm8APuzC4pErcEi4M5+esUQ9dNaBtjfYTXBqpwYlra
kRa/aPPBsbtp0Jvv64953j9NiLx9CmqF9kQudpE1utrgs61vFo8cM5vebHeO06eiknYTrVI2J6gY
eeu15MEnlqXgagesMj8lHmNRW4KAO5VVI9G0PhGXiyfsW3i+9mT+LrIDdQEGSOSQA2+07/aEudIM
rfexswsoROFPm50TF01fpT5y8nDTmLrjrJ7AIFkFH6P7mz4A7doWjjqRAyH9Nd1TokQpKjuQ5Kx9
LSm8FChAKa1uTQvHQowpv/39ZCWM41Er8jSPOj2R8Yd8GY51o1P+/ehGaDzdElvCv4yPDYfIA3rI
JQr1gVCTLrCPlfFj2K87e+Hg4nfBKkv8vytyTKAmVWIkRDlUUZg0yRKVP4NgQuDOJ49gJCVoXBj0
u8wAZwEvyBpatc39CRkfwZROAPbZ19L92beKDWM0XGTmGKW7qy2wwGrpIVPepkU2wbTIVHJjRtOp
+UGd8BcBZuWtnLF6l7ZyXscH0u+zOnar/k/Tc8sJrdLX4/1tjxRmSilTNfy1KNbfuEtC1n3tNZ3k
3oEVcSRMeNlKzqDgi4NzqThNBG/d46CadqI9wdxp2R4kfk9defD1S7fVTZY21zfZsciXflyPouG5
g+1iwrmdJGybT73eYcWSeYQ39EA12oHHOGdiRt2hBxKoPubiB/fF/mKIZhmJ+/Z8WAv0HvtBB3Yl
kfQXXX7D/kv9UKovppTD8jgycjarfATFiiXZ+kJbt3NQcxwftc0nO6pYszT/8LFYWWoZcUgAL8ld
iF5N0Goy84qBafwpFVWnMA/C6MvJe7zW6U1dT5il43TwUpumC4ihnlbb+5WngTpmFyOw0R2ZOhiC
M8H3VTJz0pbhMVR1kP5tbU37lYh/8AQkiQh42aaXvBdhb9AREBrMYU9aoaUnuGoGakAEpuona6c9
Ooag9StAm1nj8Vih6hw664jevPX1wN7z2DZ42iUhrnKzZ+bxne/bYbaVYBYSGB2xtOHFMC/Ut2xO
XCUr5x1gqKuAKIIey/xov9fIbxNva+2I0spAugIVDdFvgXIHwZOBbuyLFqeYm84MB8Nlwf3gTD1g
P6ahqokpjO0daarXK2c+avcng0ow3Kj5kyFZElgEDlhUcFbqF+908Nec/2wShHIpmCVGfeseJR/J
r+gyQcR7smqsxR3x+MCyVSf3ZAoQoZKHvqNcxPirQPavNS9J+uhiL1Ppo7KlgPChcWpCnfCrl+Ue
MoRgV5ryJR0+wMh6j0WtlO2SMAIo0/UJbAwixyi3BgOW5t8fkParR3qjtJgufDEnV4ImpIPRm1HN
dbXGJbWI4CWZEERPl6VUILJtKURfy2pDbgihsYrD6nhrl2mV3YiU1u+fVqOtHTJRPr5JavY8mxfH
kVmO4R0rmsul5G8J/VSkeXFZtaLhdNcM7XwsKVtcA2Rw7sng3Yb9yKGVxojAPFwkhzxrHnxxNvlW
moBHCE9oY+/mQRQ1+NJeKGaJwNCRDnKNbnci72T3vQc+tem7AkL2zjOcGZfGvYedKJE/ufj2Y1xZ
T00tC4eTacHBysJfCKuxUMVDYXJP9DG3B1vw/MCPnbxHczHJhw/8DNfmX2rhrjbZ1WpQxbZtkbY8
0TbXEJDCtQSLRPcMwHxP6k05bIYA3oY+DlmXJlY7jIhIYmOMs4G/A0jPTrerRtAl3ogs3DfJVa7e
8r0K0qKvRp4TV45Pd5q0aldAJOrcgmQIAeH74Jl6EHZiRHvpzdrmNLI03C8Je+kjaF1oNtlYizIz
abeAuw+Lxygz5B+9XxRHxcaZAPx1XMzg+YEqmqWSTIITImuwaBLJJMgAOy0cNFKRU70bzgfHVqnz
mi5CVqIflPKk60Fp6UE0waR4TGitJ6IySxjevPXuhJXyMNDBlxc/L1ohvVqM+Rt5C7FkTT8kZbqA
B4tWQec2IXtjo4E0V9w3xiIBCePgMiqKgz4C3tAoMitijcAbE4EREThiOPr8dKdm9mRJ79DMWNSh
Ons7+WQ+s/C5GEIy9MPGUEQoDi/pOKNr6uiMvv5SUJNGR0/wS7LlO871QwJenx6oocD28nDuk/nr
s27wT/LK7tkhfV0LXRqbI90ixyuWpJZxrQsy2SksfybKZp+/3yt86LsRfTfRByhYfKPH30kzoSbi
a0uTrZSxtbi5CdigOVzXoG3zeCctcPIIuV+WUfOdRjKNe/ewd+OKPjoWVIoExR0iizv+nifE9O3d
PdgK0ksstbsQ4kGouDyrB/F4Z6+mKTgY+TlvPrZr6PORlBPrd/GprwdbKck8C4Dp/+tON5X7vxSc
/zhtANMjA7nRiQ+Ejl1O0epH1+R869SJRIlPWUbdKzBELyK4fYJX1MK05Q0rQ0KO0fQOJBmDBs4t
pIHpOzPEoJRkwmSodYGkV9HH3Gm8iTiaMP/CNnab38LqKhsdr0FGZRS0c5JdkSFJkAZo3549ERV6
81YPb7vynzY/7A5T69r8jyC2cEBC13spCrR4aBVoBCZJ8qTs6g+xnZx+/c1jASI9s2vKRLd3fYL/
zP0DR+2oNd43H4+wZYo8U+tH1TOW0sI6uJXAN1CHfxa2dimG87ykuqM1ihGGLDSa2U1xBOhfkJWP
wWKGZtEKHlvxgQjDmIph7UU3Yowf8a8brpK8EXaREMsKdZwxEE6MwfIighvmijcV/PyFearz1/ai
iN3+8+86K7M85hWMquRIkOvng27vle5fc9gOTbT0ySc4wUFTTs6woQY9MijKpmIxiyIChql2sL1z
Wch9L7JdPndq3QxAELsQU7u58GHtr1ISpi0/93X1fdPH7bRE2hjb6YfBDp8jKQ2D5iwGbKuRkmpj
tGR5gNjkrhwcHkp0EFSEQK5a1L6pqLJV6afZ7jKoTCYJQDtHBlTxsCtNBcs8UqDUcVt9OPVdU0In
/IqsAnSQx0kXtTUSwSUkJrb0MPMOMqhpKubTkbY3awN4hXu9rVE70b+F/+wqfExhGnwWl3o+o5PA
oe77WCcrTGRxC2qo2kGNVP4BU6+Kam7LZO5IQj0sbTRHMRIHJ621Uw/8FQFsB0VclINVRjYkzP5l
7f3Om1A1gOxgmWEhIltkJmD+1mwkYliTaOppGRA9gsIOvvjwHoSeBNpWbzMVLFB8ENhQIpWCynhh
hercZ9R1IX8J9H6SE4gpae3C1lstfnjfESkQpmMedF/NBwa8NQaTVkOtBUqkydvGTsM3YKHfpZTm
cd+QpaQdpSpw/V5vUE76Dr2HtnnodiDiC0dUvGUdCtt0CexCEo3/M3sUgZGkIVUXYM2OOGrFffk3
5eCV3PBl6fM4OxVZ/tnfHTQZXZ75xjr2x2m8aWyA4516v1ZmV62NHSUIsZGMZLaO/RnGDWIpyS1X
3T0ieP2fwJ7jg2/ptkkqUVQ2IljtbsXwsBu3CzNytrLJl1gRwILhANauRr0tObHiWfOAf/lp7jEN
wB+aWROG1bcWftSVOKmzCfYDcPfkg1LM3Ylp8oxrkbI0A47DvuKy+TrN8IldzNUv6H1Hbd5lFE0T
/8V/YnOiX+WZtO6MBzrIYMlHqXigGS9rTg/X3oVbZQ4nD0aaC2gSQjccts5BnVyAuA18AU00mfkY
GciQYalh3bAOT0NVwof4nPH2i9vqxJae9s1foDtg+keWwgvKY3S2JAMWGr6drJ94FgE1CFq7paCl
2LWa47zytTwy2HQ14QB7GkVA4taaud0p2XTrrmYD/SVJFImFUfCwK1///He+VEjQ/g/g1aaoVlCg
GJJUixVHkbxourRTHZfQTkn1Ds4LbaplQsrd+7q3KvkqnyGXLx3Xfzm5aOeKEx5U5Xmy+1bKaKw1
dOTpy3eqKk1i3LwsDgZLf39inJYC19OhGgTG5kDv+C4B+OcmHLTAVt3g8FTC5Gx7VhUotRzvWvbE
uY2AvmmkveaIE8u0Jq55qmYynPszZtts/ng6b6Qg8CBfdlbLxn3tTpJDcks6u5yCnm+bt0Y29tg1
h4pgBpXVeeYtmHPf+UupJUveHmPLF80bg3gNCmNgvbBYYQvgS+JuaA0tyYK6rgiRpnbL472QOEMN
LOXOtOPYjfUlcNfVejkTxqZRN4ZnOA7GW/I7RxxRCYvFpMokAfV8oLD+HAguzQ6Q3nABsQSOTl3O
UGKBFjfot1eTIk/oFp/NwcizdlV/W3ADez3L4OctUtKsqB+572J3sSqENn+kXxtzrMxAlYPt5GL/
pbJbthQyi3oMTzG75HuSh3fE5QwS2MdxjPOLJnjThgUWyCW5QE17LaYeSI/yzfMQVODJkzSSp3mS
k2+VIRHwIkcMl8vvQsV7I3aibFD4s112twvS05E1k/ijUNMlZQJGyq3m54wPT+wPdKndFhOiXvik
RBA7tmLQf9Im27aanrO0GdnHfTCT6V/hmQS47fACuHYhgyS9m49ku7c2h5Wbwu9gCwwoAqJfq/aX
51gZUx9qRRtQdyVVuf3U7uCGGwvdVhOECakaeldsCoSWXWzYuWZEz6mMaYMdZtKKS7Xm3XdsG2b1
Ah9foiwLMHSmedqBP1jm0EhNzv86y/sOV11mDtdAe5qy076pjeinmDuURRxg+b7NybYjDuzsUG9l
I1HcuxMz9fsVUKZcUWJ7t/VruFkHzL2hR4ote/k+IiWY6DAnrxSpno/49ctkJUaNsi6D54ksH7mr
7hWIlbKrV+xCo1WGRf4o16JMGDT24AeXB6CfOQse0R2hlvED3haJEJKgn1XY9YRqK+qzSh+MwmI5
+An/2HMHYP/Uuk15zghrewiqLU0iV1VG1IY3TZ97+THk12MMZzPBXas1qNNkZRlTQr3GZVmR+Ia0
unB779lFjXRwvQg1JfsDK2v0VXJ3KMT/ySHqBS7EiFmo41fTA3SzHSKS4YztmwZj0XNBQPigoeu/
Wk6dS0KeEcmLjMWUfDaF3MfQRuQEl03IYi4WrqfqYo7dPuvr7NbTKnNBcNmC3H0Spj9sHLNwl5/q
lIwk7kLhBbL/FrcRuJVFOHjQDFoibDYjMF+CZcBDsQj/WWkJmVpAPdqQosRMTlR7bxty9f7gtIcQ
Ym5yY0eEVEDx9Bhe8h927XCJUpIJNB9CAY2OGDASlRuGMghtVkp0Dwm6H12zKqNmqZgfBZ0mpW+8
hmMNEL3FN6Zzl0LIolS5F2EqhqOXst+LK3wcnNxX0k4OnDHiQQi3KOSLWhD+Vy3JbF4Rlz2mNbNJ
MTX+4vpLt8/ApIQHQ5CAnDyQh1MrA5N+/Z4bD1YMoDo8OFOn4JcQLHG9zNZQDwVxPY14SPTkag/R
X1qsibcQY9md9NjTZgB+Jga1aofpW7h36AJjPUkQLOiDkJ2UJKZ80oMmjr0GulKsdeO5crf/UV3v
FG/bRV0GbX87O3S2Z2bG/3uz/lM0JM5qJhRrBzIYaXJtlPvC026xiioi2vGkNUkgbOInpjUGW6ym
gw5eyjdv9F0J2NjOiFCzERJQaH/7Gzn2lY/pQLO4/8hLbpxDuiIsy1ux/bKAeYdSykrNLGHynBA+
MXeOZkhtBRRIaocnaoX3iYE8x4BXh/E4YQa9ad6LbZpO4t9j2QdYdLNVvj/E9W2oZS5vwri+Laq9
uH8ihQjvubB/t2xyrxpIZQk3+WUrgsN8eIp+ZTBWqMEaE8SVH3M+L0IQvUAFQLbNWQ8FESkfy7VP
dHRXQZVmBvPSgGW9LFZ93JFs6wv6tmZKiDxCA0Gqrd+XfASECHXZN5001F2MghqzVK9U3dwyVbQb
Cw0nrHTEM5woQzQMlwnx4b5mEILs99gYPAK/lHjQ902DbWX8m4ToHyf7WLWg+PGTFliOJp+6T+UP
4/vWCoNP4H4onL4JrZLr+LdnlNTloiv5W0Zggbr8z2NdLhqp5iCXOZJr58PkcIpr2uFu+e4uaIh3
M/2Lr6A8NBc7Pt9WjFtyAF9oTIkcVSjVKxbEobJgskyf4HNYELGx0bGgNppAryx97njJ2UciTBd5
/RwK4XQHlXXRyotwa7pfpbbq1UnFLRH/Zrn68ZhWZskxK4roKtg6eIPqghEBvYFFuW8ngZU2d8Mp
PpWEhXKGnLL/nccx6iy5o4ZdnyWOSAvuD0zllAjPkpv8CbxQye5e1ho4Wiv0JEkCdveONkLU7zLY
npaHtjKKvu6s9YChPUPo+EsaUpRuGvU1GHdvY3EaophpXRopgOVypVxZsIuzvW4nPpIoCVpTp4mC
M2le+5hq/eRKm++kAXYQLjOIq8v//r7/ydabscljQgfiH+R+F9e1sw9vLxNbpRZHpgbRs2085qZ5
mvnt/z2yEWGLcSKdNZZU1Hl2ZTqVjGeDFBNhsHyBWXlGbevS3RAJXNJQ+7ocjikHGBodQwuR2s7z
+IuqJN3846xN+brWinpQrvXybqMUZ/JutMXE0e6KjwG5cQ2vyW58ZiJ2UN1VFFTo7uS1dbUXQzNV
OK3gNrXudUcjjzVFw6KvMzn1fLhyMXPeW0jMwB3G8lgq5E6+aERtS5wK/P00UqNZaNOA2/g5QrvZ
1CNC4RDHu9wBIyFLcKD2BMwfDAGMVNGCCHN83FIV5mOwcHhH4iJGpZLNstmeoLmY7NyEdQCeuSLi
HOwdqe0gb2/uWFDTGbJeIZtpVtrH44t3PBUDIT6Epo7Xy8nghMbfF9OIDJK/sa5SaEIUjMzXagrk
LdZxwPZIM4QL34SMVhYSWbYVRrseHEVzHE3GKJ6nZgvDTQaWmVCrZHxSW4L8IUK4MEjNTrofLNTT
0ehn2YOGb9/eHHwlzMCIL1nx7pKRl/xm0RYa9okToy3MD69aulI5N0LfK9Lv35diSauhiWB8zZvB
HFUHt80/8+XRl0/QdOT3N1cZF85Npu8CGi2vy0l2HuK+qcLbj+fJS2iD317wbKpoh7SNLsv+7JcF
29Wn6vSuqdDgjr57USfLlvewzteuwp3ozO9R8BUdtqupU0CL32p638e782o6S16ee4HzUB6IyFTa
QejdykvPRLB9eONCWz7fPoU9GuXDwiTttUmnL2w8d52RfvUkrZQK2V/epO86itoW324FrA8db6ar
FK5rFAuc87alUsN+MFFb2hJdZ1RF4xMZ/5Ve9yQvj9EYYrOcevQvpXZp/gpTSPg/20TWPz0uROCm
2X7xMlImee9qL7sXFH6dAAxcpC9Qdn+CqSZUrME33qTZmsdkzWWd5QmKp4Fn/+Pn6El5Vl7CCOpW
EUMSWZIxQU+bBT9tRZOBrWDW04CL57zJ5yrUtv78WTfzFTXUMkhnwRBv1VE740De2aAuctzCDhau
NzbYNJJxo+bEjNCMOMFo60iX+NdpPsen0LWiXBrKNIYB5UgMq0nxfS+L/wclfOkvoib4E7s1/6A6
G980elzVZeGF1vTPbjqu1/O0dyTVo0iHOIJZhG1/AulNyFprnKQ130Mr2KwdAgkFaZHES0PHlF8W
E5C39sD5Pp1/lY14SrtQ4KDDkd7Kf/HZyznbd0P31G/gAC4TvGS7ejjsmewh5Go1JMdt4SGG3yq6
63pPo72S1vcsB9ustTCKBuLTslRqnVNdwVEjWO6blCbt/Pl5m8k1q6l2CJXwCseyzzm7PX0fKXG8
fO2llAiBjdIYkx5RQI5P0LMFHXacjIs667CnKuvJmPSrMIv+ULdAak6Zb0cz9kJh6f6aUmADjbUe
jyNPvgOocsl5fp98I0RrYMPPQOYpYEfEjMT5V2nqwj0HLGjPBwiir30tktSuf7UcYE4EZfQb+PmC
rTLAlL2ukNHCD9Shfrkf15itppvM6JmTvkPLtEVPD0ZWlXQAKkZPWxL/9u4akw/snDPZG5w0OwAK
z6VcPgVdMcDUwFgSpbNLFv7vjeYPpfUOwldtyTm018pa3Kc+ev9IZzdSNAClvosU8rMqNqTwaqlO
VXMbDNitV7TXoSDDX+gTnmD3uB/SGfOTznn/AsrG2qKa8VcosL3aUCrKUupVT1lG+bjUyB1cLx/j
zahCv+Zkt9e3o/6BlD6CliK+KmqUzBLeuo8WTD9ECrDflRz9yKfkrAMP2IaH7hqgNDq01Wj/9ClD
2eAtRga7yCWaFkV7VJaz9CxsOq8ifDFADUr8DvDxFG2nP3L13kETrigdoAWQk2xS1hDwARmBn1Gj
CK60+2GqudHHjT7c0vXAbgExAKIUPvRkKUeGHvxH98kPtGdlRsgPTOAMWreMLtPblx7buE8QuFyR
JMEk5yR/T7uEPxuw/gSKopiSbWnmr2r7uzbBZN16kALaasZjT+/kkSWwT2iTXMWQtK8XgioARBsO
m8Hv56E6wGBAvndy87HWvMni0EFVAqQnOIwkvCvi4Ok16Mwe//Pi24TEWLr/5LcCYEM037NG2c4Z
6qM64uw1JEzIU+axWo/u/h7FfPsq9mzWESJqFt4w44nJGHZCt2ejvI7WUL8E+bkZyKv9gpb8tGxA
EbJv6WgrazEsblOEhbGFHIlFW5oIHV/QAbR65wGfzJmt/+skf/l5DRnVEg2wxTFLv2KLq5u3x8ny
KBjOyQyeRc+sd53iF6HBwNP3ohR5PhK+tNFyQOwW9w/TgZQjx4h6qK3OaQCnmZ+a8BJdNIYgJonC
2dJUdK5TZY4i5MU7SKKiY7atmnPLodBLyT7d5Do3awYQDiuW43FYjUAh466N1BxrLjpQqKa2/vGy
lq5kPbeUCAMtt+/Vc0tYij5PQNSMbL62V4Dh7alh4hcMOCUcBVptrdkze0zOlOlaKgHZ9LQvLDLe
yjI864TsKlMlVdZHldVFQx7KNxkTRagPe9M8NenJ5VLvKlSPhANMH5tWnF4bmDJlIXpX21fMD/Gp
sxEdo8Zg5KWHXn1sjVRRHRDXfm8WyqA2fnMHRvuIZpjQ0pPG16MuZtYVFilvOTwsJxCuV+W72xL/
f5KGhF34ehj6+SQ8cbwH4j06xSgdblcpgIGDRPl/vrrEmH17cPgkxiYv4kLu3Fwk21vCu55Lr3vb
cZx5KW+pANcZKxXL6GPFsnjkbAeVsOj9dxZrqJEu2+a2fgIMnmdO1CSgIosBc2WErzaeMwRhHDK6
ztHxJniCXo+Fkse414BoAelurXg9YGfe0Ssl9lBnqBlmZ5RVDDZIePmRWiBxKm9Gm6VORur07A0+
soxl/HMK8Yg6YCO2Y0KsOMEbNEYkvoINm4oltfyCz4GBE4DQgcKImY+BKMjtgezc7ROlFP24loUw
4JUku3Hs09bRezQ8Q7pJseAluAgyhXmP+HlVanYoerMhKdGXkluFBTrkvH6OKVbCkjOJpEthmtIC
OiNoaTuq1tOcIHDLiqQCoXOpYJg19Sj+/Bzg5TVWbvlo4ZUtIJq+m4b6tHM8+QdyNYvi0glm/s9b
xKZVVBrPUgUMjBOdTaQbYTBuzYj4J0hJUyDMpOjq9OQzI9/L1cVEN+2t04q9Vs6BLaF7Rdhlgn86
7Ax+qus8VcPsyArvD1FAJMAjIg3iFHh6cB7fcdFi0f1LHt5yZjFygoypqp0NRuUV/w2QXSconeUP
U7/aZ+Z0DwL/FjBkRdKVPt4NwG1HVSuGOfXCC2W43ntQVJ+37te3bFefJzMj4mbAInZNtpV+scBK
VzvZMrszyOSE0Lwp9CzSNv5xJqLgIEk3M+c2lDhhjxMuKeIgnXvniRyf3Ls2LSr0yXT3ZwULKW/t
xld3hzQPY1DiNd//MV4kctWg3I/+MGyiyHIrF8okxJnY8y2pw3wa3RoXHz0PMl7v7diIcVvxO7Ub
uiMX6/WVOvboDJr46keTHYc5yf/IzzE39A694jwM/H9vJ0snXwjLjj79HeNekOMzdMajPw8n32DX
JCGfJcwPo/Ts7i1/Xl8VAGkFa5EwepFeYXDJUIDZFmPV6md36tlWzbKPdiUsWw4kZfnRiDMvyEt4
dzx7rdcHjFPv1sp/J9dfEdYZ5oTuwtuMzdQRvGlAbhYMaj/Np4A83lqKRamhQ/9Na1nkT6ikmSlL
fBPgu0FmUB30XAIEUFH2NjJA5LN09ouRPPYvmcLTJTFe02ZIrbBLnFsUBP9suzZ89mVcvzjeNHs9
C6H5Pj5bgDBxXtYVuaQR4rf9KBwgBnBzPP+amKvR79ANJWz/j3XuBoPuL/QZXEdQW7TL5VVUrMnd
V2lc8koPOF6ArtvFmZHRsG59d5+dWxG/G4nX3tZaLVlTLsrX3ZRlLljxuKeu7Fx0vNMYSXNglJAC
QMnqcVFtoc98W6DcRztpqEnmuj4aYL1n+S0iSkbJAye9zDTzi5IewpRhaFSUYV+l/cF/sgsawReq
PcDvWKqpyV9n3HovGX1gsPkexS/AlEi0OIUMMnOsO/aO1dKAS7bs0qttLexOUn4vYIJdikzIVcs/
QZSJhKhC8y+iYWQG5kF/0BlxT6xvOCliCl7UljSzwoT9YO49YZZIpuG9DpVPdZPP18ECa6jfrpc7
4Gat72zb9DSbcSzee85TgTibTfOP33vyh6hCwfIQ6H0gPO/bw0N8BdO8z5BYRtMhTDFWINai/4cZ
SIJDYgedeN7Hw1VtXNW2O6+wPSvJJ0rmBrNTX6/sBNJ3tSA6q+ivs9yt4lXmCJLG31bgYZdJmSbq
W0uIZhDD2QEfRfy1MkZeamZ+WKOBGEJGDtBdZU24nO5gl9si0xi/sEcECxr4LpbNAZKAh7xLwtYa
ZMUMlZ/Gf5WtawV0njnZxVenebm20clIGjBFZmnh6aQQnBr7CsJ8ySNO279OSqqd0+DFMJ927Wyc
31kffcDmRRJnsHGm28EnKQ6vqfrHVfW1Y+gzHYs1u2zxHN4+ybQ/YR/R6I7N08jGMYHUlpNs9oBk
1wNQTUPNXfxZKmgE7tUREXXteTzpjT8LfOvRRBgUeIwGSyBCfXUVYdulKZaUg37iEb4U576uvVhx
xBA7b3KY7Uh9Dj/h0NKg40iLxy69DniWC2c7he8c8gY5Y4++BHxuT0fqifXY9MULif9ZFH6KOaot
7o0X47YrqZyuq4ZLOMrYIV3y3hsRUyg5FcPCBVgfTzcsRKbg2CPS83+Mywyi09bbC1Uhub39V0KN
sb5bR70wu3kb6GEFL0RvPX6X/bd0Exc28c4jmhrEGrju1nfFE/DHJAkWvlXvZWs+vyIKfqyMoMA1
K1md0ckeCZEsCaIi4ZJrwAgjtgs++UGPYf8WFnyrEX1QyE8ARCBgA21NUZ28aMQg8ExFyrNS5fsJ
Kw5hAufXpOtIMvwOXDft8gWelUBRpt+Htl9If406RN1/OY8zGt6JZYe5hUW35AnzevmjV7vxcYUj
98msiWYYFdcNjM+p97XiiFkBflqrK01LUCs4SHe0oohnoZ/RC0GUUZt+FtnUozAqBwA7YcDF/KTF
qsOjG1GnFcFbcVEVY9DJa++eed2Oe0sO7Wp9zWUg9lg3fDWrWSf4D/wnxxHiKqciIMj/a1Pu+sbt
GiNHdZbNNgsV9v+QXCwJUrTKv7mtCoS+FZCrKDH7l281n9TDxa9SLaOGFu+muOETQ/fSKfLA4ne0
JHtjU5QSAnDnn0vNRaaP9Ll2Esx3Nu3BSnvpf43/qSVc+H/4NTyYPVVEH7hDaSiS8fgGqmvZhXaU
IV8HC0FsgnakhHZoPrA3/GX2I8BrRDg3mhsTsFiNeZJbtHzmjuKrCnLXKKJZXRZNIC4gSXOQqdmw
UQZ4td0mByFrBvyMlS26IzfHb6vfL4VCMFnEunzJhDc9S9OsA50t/3rLDRu6twK5kuUsr15iHUK/
4CtVmfKi2cuKKWJC3PHh/H3KcYrSLiqLSLX65uHGdYtq912BbjRIF0F2Ac5+8pxPyuzYdkXOO7to
W+CFyin6CdCoq0ifY36/TmijgjG9AGSbHVEMDN4Muzbe2SaC578ayWaHDXXrfS3B87dcvoKRybo9
9jqHjaWPZcDAZPGHpARPnLDvATAxCydC8lqIgruILk8urulhAXEyuT0BUmy5g8PNS9CbSoS9VY1W
YUUSu2s7ZQ1PEcbm4HCihSEpzzIb04yxPcs1Dn09XxLcce29yXDWP0OnNNQdId5MmMw/10EFIMkl
ndG2gC2qo+SM8hApyHJmFdMDKhjeqxiffWE24EQ6q4XhIG15V+C1NzsRCxWnMCeT95gQxdML18KW
YKUI6niOcFbs2P8/TvFRd4Th497eC8rriZzpkSLBrLAZQ35Z70YyJEkrUv1CKmmMzZz5H8nr2pyG
Y73axwEp9cfw9u6Rrr7pVGzH9Beohqs3913M/UJ9OoQLdYHML4BSN5YyaMSJ5kxh8Pd3zIgRaaHj
VUeNfRdEaVTianKdlK9SIEIrpqZPaQJDYh8zzJaFZBTkZBtXDdcHW44sn7eOpcNqG8G6L5eL8OWo
2EWwo7kNtq65+HggYPgaPtXoBSR6Ftc5wgUUEYSya7IuNYblQ+JAwq0vL2KU0mu2j1zbjz4P8lU/
3Qcfql80aDhJW9hCzAm26Jolt48CSeOIaS2SnllpcZhe3P1tYsVAbBK4CiOLJoG5BTLLsaFe8ZiP
AiRgNw42/nZKXqRgGcLqFGKACiCeLwyPWAb5GOWnxL4w3lU6g+EbKuCv1lkCQppAKP9DK95VWKFk
cdygCwC/n3zhw2SNpA/FauhfuYbw0eZBLEicHz09SX/U74WWfHCO9nu2PjliSdWCHvwhA9wJuFuh
UKmBmgHjjWZiCijI8nA2Aj8MpbvUaah67tOK5QeaUFVFxYJvb1tED4mirNgasiFves4dFPHD+0hk
3N1aV1JpNHyFDCseZwdf1FFt/Sc3Lg4/D/Q4xLNeaHhOvxgYzYmM1bNA2ix9oEivdxMMe0WUsB1K
bI5qfUL/7rzQhEKBIiP7EEXiqC76UweOpZnx5YssCdRUAURHrKGzqrxHW1JkQN7zqiNrzS2PXkMi
zESAHmDtKSDFY7Gd6CfpSRWw5gkSbRoG5l/+wz/+Upfipu58MDq/8RDwZclE2cW0L30xw0+2yN7C
dFV9xOupI7shzeHiptwXJrDlX681x3s/1qcJHQk9jZIyvK4y2f1do8zM8wh6MQY+hSIgiSc8gZ2Y
+99wmIJ6JfwjKJr/DtdE5irtD78jGh/dSHNQx71UzFLYXsDqUxVZg18MYfKqZKBD3FZigGt9920G
VIwu0ikrHcrgTBr19D+SXGDQJN+sh8IylXtkgON/uOmcvVLYefnddq6vCq1+lz7bvCvxx1omSD4/
2UixNbmUswhMdjiTjM5gztAIp2FwpSS/V2+Lz4ej+Fm5FmDRI3v55UnORd4BjhK4uPOpIjlj/VIE
DrMiaCRbC1+UMbi3Vwv365J3w8IYJelijbYUnHu4Bo/QCXySXWh4+emI0gzkR/q3aQlgcG8Jya4z
J+HP8EqHMw5RcQCNulQTTlbo/u1Xg2m1HHJtOrXp9dbHQcR3dtLgYizyHhtWZXqryWIf6+WVfOwJ
vrJrSMGWNP0d/ZsMBtQP9tsL8kSjakzKdTQRTAuJmWvOmCnN/c/a6VQrHgFdksxnORFE0GuxKx9L
yxI4tw7FX6F2AAzci3SrCHVL78NkUW1KtSO1yoRxaJ1LaAI+TdgnRWeW9zin1+Xi5Zk5UE0xmpnz
Vq0D8VKdRHeb6zN1Z3dH5fCsDNOCsB+0Bgd+EGQ1gFSo035ks5h35ZXGXhTfHmzKd+hzy/qs5Scn
BrVow4WOLdlNXI88W3K/Jv/v1ok1y1LZkpzWxYkjxZXr2rcbDjBhdP+lch5DEijJNXUUPpfAWIPg
zKuYiB4GU6+N+JcUYeihovLWTYyUT6+n/I82xRnnHQP2p1y0wSygTE6NwrZX4UyYDk1/zfp/+q/r
flup6Y+Hu7Z9NudItPQ2ZeNiHgIo479U3Q19IlvHl4K8pNdL4uUPLBcu55+62ZIrKc/4O8RHnTOq
KJIww4j3VvBtUpw+VcZ/kWMDxRuVDMHbhHLT86YwrPAVN2M8fHoj8ibKOEW67gqNagjKUhJC6xBd
Irh2exGNeLk1wI4fYTfNHdHyDLzy8/iEpFYY0Ev1xr12R0r6UVl4+Q54S/Yst4kySjnXlXoJEIqh
5VFsy3Ov3P6uPtSHDCeTASA/ocxgSnuU2SiaAaJ4nSKjhqrbCETsZnH9bbNlSnMuY2wNZbhov5P0
ol1FNWy+rtHGMAxWwyvfjbcGYq4aC4XCDuyMEMuzv6qfYeGXiCeiGM9cdmUPeXWUESigXh1sfatT
rdDE3zHFTggkl37kM1Y+e31BW/9xT45poxhdZf1eZCkn9PBFY5CX8KyUAOrKFrMGZWVTZAnCaz+e
Y1lKkepj1l9mPZzikJ/ytco6Vb3/j8rxUcvk7iZRQ0syOceak7rS1GrfxJcWIUWZ5+KGm03hW1/a
hE2gsynnxOkJRKAec3whhL8DOfhBgrP1AlyxMI3tCeIOMsNPE3AIADUlHxL595+2tBzhqxPTMeeR
G+FL75iisfRjS8IKQ+pPARY+ZBNyvJE6b8Y5aKjCmKyienUhTYAlYJu8+a1m4cbr4YOMvOtSGMaS
paYsD3BN/+YJmcf+Bs1v51qVUwTUlxj0/c7ZqviXPVZvHycgFUGberNkl03PtC7FvC0br1uAb07a
kgxVtxNYMIiWNpl24sowfWwCs8qMW1aZR6E1P2XYQKoTh7M2s4lnfpJcW6oGmJFrFs/q+SQ5wtlx
bQfSs9fSymBnDJm0hE8mETa0mKhPbE0PTgA/De+O/vJ5UqeGsfd1cVvUvPb48vvW/puZXZHVO7ss
ziMe7lRO8BKdwZd0n9M9brmVnDwGrG7b1Bc+0cU8vdq0hTvM8yiQYmSG4tfXk2G3Zq4q7qWy/6e+
D2WrFADlMAymPe5tzkJjsgm2Fj3QhSQRGPwU2ENQrkU3UI9ODqUKo/U34jgFiLI+EaQtA7Y8s4+j
lsqVejbPOQOMEFzxeEyn6bagtzxzhy3RZXLdfBACFTY1SIc9lieygL9/bZB9OrP3Fp8nc0pVH0+q
7bOmtZNZqi4OiHktdBRj6ad4ZMnvTVAtRTuzW1AO+0d+QQzzr4IS4qyPv28hbrCpWP+d5NSdq8SS
Fi64dwQezklIZViosdmaTzqMwKK3xzsWC/5uCc02pju77rkPIuNVc8EE4VbUdIt09YlieNgNfRJJ
hhKI/7ptT+BdYwtO+LxwEiuFUKiVHT2onzuv43G/+/0LFGEq4C6Uk2t12n4RkJfM3LDy6C+iYi3K
kJsRNxwGrmL64pHLWRuv532iIsbot8K/PUqKRf+H2x/j4TOhfBmlJ7E5GPeDISpXW/X0PTTS3iZr
nIHlmE4L3fL6AJuL5VohxsGbZe5bKtf9X/GD1/q1tom8ugkgdIdhhOn0feI9Rxt7q5mXfaOrF8ns
sAas/2Wzlnf/sfescwtXoarcHf4JPQYIHi3urrW2Wf9okns3N8YRrh1IsJ1yqUbm/QjGykeWPVZM
E/kT+Ytr4UsNXQnQGFDYoLRkjN+jqqs5Yx1cAqHvpg2SCCwn0IyYHe9fyQmrzARFFpVpWUsAnyy7
lvAGBAh1YEKR9ulK06HxjLKIXunliRRbD4ertu9vnhv3SYd1M+43RMVMyeyXmL0Kyo4EeT2MGq/8
4IkIQjQCkeCR5mKrWVogPpWPU9ktchstqk1HZK71yst+TTdG7580Ltj4bzM7jAlRx3n9zkhD+cF5
HdRzd8M2L/hUacpE888tJFLJRYAMHbOy/xWDgcpJos1QJjNFhn6wTlLB/WRJwb4+D1yznZ60JYBz
yLK0Be0UOi5MhqOKCKuw/Va90OxpE6ndcizcbLjMeRLEhUeQlGPUoPPuFfG4LUpGzh5NWUBMoSxL
D1BtRwCFQOkdVXzDuO49PfgkIdYdk4qypxGi+kDcAjmhp2qe58kojNul9SvMs1bXqKIp9K+51MDN
YQnA7UnKrKP38dpDrvbAC3tRFPxu4Xg+Px3M9Uqwxp93EnBxEgGgIUVljhTTLZ36laQTSxDTeIoA
7+5mjll9WADfrJra+vqIh7mli48IC9zV9Wmhr1revPCFewGw9yzzJII5iuBFEP9NcXvVv+A2Vohy
7A8etwPb/op8BiSxgmvCt4ii2ydA2LbnSc4NRg3QCENQc8clWr7NbTna5tv6zKuCFz56JVzh9JGn
aHBneT/qRkntk6Xid3i8zm0+0oPyfZ0DI3IKvbcTpwtM+HX0OK/+Rw5Qu0dttZ3BMPQH01p8MI0Y
QkEyLcYa/Uew5wUt6LHSgRXNgyaj1DD6sHTqStHxMukgxFGiwRTIq4ok7C0T/UHDrFX+9/+crA/v
KHABZUv19GGd6NCAzK6zYJKtFdFJxQQ70WPDA0YA2csP+taubaiLF9nmwMygDjofpfN/l1vpiGXB
2RfK1VIRl28kwuFLPJT+neuvM1p0nuhIriwfbtg1k/url2JZFI+YDAiUgsd7rMiCgoi+46XkAV8j
P7NzXN3uibhjta49vAWEHmTlRrZUDZcTe3ASYGOF4mvOglIUnlCJ09x2p0KgUbXnDxexjJRSiQRU
ylC+XaRTOQc5cw582QjTJPMepZZ3mWdF2aguXkbLzXPEQQBDcEWEkhTYDdNZnVU0rfQRFAJ/AKEj
jsgdq5HX8W6hWRnDzMvmR7imRNkzCnYWzWp0gE86qctBtnRncMhcj5yM8g60XwKGx5LnvzGR3gS+
cUP98Q1LB/T1/ZFHt3U8IsTiChi5DJdNHLY09l8OyWCfv4i+iWG+mQhXcLiLHXfhuagHP+W46giR
fLBVKcjUduvGlvTMo8RuLjtesKCX++Qv5KOR/rZqXkl35oufZOIWmLMEKujaaqm7t90wSBBVPYCT
t2IC6+WZLl2S0KNWqBP0YpJt16o+U0XUbWU/ujdEWO2tFVnmP+IBrEAXGHT0ABp2k7FnN8jjKxT9
9yhfzNMfPjWlp4nQaTJ3IiFuua6kRpxNkmqjktner0WAM7AqnpUP6JFCbhnNh2RlwG8UDVlAMF17
LTuAcVpSk83W4eOjUnfoSW1Q/6ygiK9daaOmcIxGqlOkQOkO1hAvuG8IAjbgsCwEh+r27VBG3l4A
UaaV47V6YQryLdUNtYVLCTPmDtSFXqfzB7GSpjYpvMZP7MTXSZaShzZQ6KROpkhHmz2GY026cyiP
TzWXJ52i5ohSCRCWQqtoF9wr2guOw3dg/bl2UCD+6jm4hr+uYDVyHlL0iLB0a5OtEt9PFN6WfKqR
iDMoS1utzM2VTxozEjEtoC7s0CQaYxpGPr7sCLSeAvJHcDV1eow3e0nuYbh34T34y/oeBp90Q81F
yN7Jwz1gNLr0UKa6Jwk6Y4+67POVOlZ4mk4nwBDrahsWAXizqTbC5bAQSFLWrnS9gFm/gSyGeWAw
5DrBYrw9pWOZ+DMahSK0ad26ZOGq25h/ncgaW97txXM+T83L1eHU5tOs5CcZcJbCq7g3yTvQ+lvD
RGeLM8oS9ebEdCCjvivzmciZPzAzjK88jYPlCzKDAjde8p3T1lB5YN51JEIod6qEo4Ybbiktwm/B
O0PkEKcqdH7HrnUKxXkIm5n9My0cxK1WUAf/FnDeTxJ0QsNsgtVmCfqoDJSGhY0konOHyAnBdhkB
Egr56dX4q0FBJjyBsMU9Fy1Xgap5a5Stk7Z3E7HztDIh/5pM6NcRvDKaSxOoDY/uw1kUcLjRzPDH
DnGweM0QY6vXS3kzbKuLKkiJNsXKBqeBS9w5b/j2GKSx5nsUqDZUpkTvYfXTcbTR1t/Ml7zdKv54
U80XVilCUwE/L5qIu1Os18DXMlNAGMLQPspMK7ePshlIz5tzBXl67quz8/aijOIuMT/BunY5mBck
q3jcnBLUmnZ6AGzhCfVxgvs6JO84qbXt0qGnMYjFc+kNTrTMHNvPZIA9+jpQfKbs8I7l0eJFHKof
0ZOxlle49q9bfkNL9zFyKNT8/yDM67KKFhVdrUMZrQkGVwTQGjcxhO5lccRSu2GCN+aQSnGxgwAl
Q71QZWqvSksE9vNf9ToqWteqWwKR7bUqkiN2qh593HWv4LrA4MLzDzP/Ocuh12X/7J888c3i8NYD
rzDvdvd5OWgNYbF9EQZrBMWxXgzINe+ZXHHhqz5Iv+ptPZIpZJG33jSvMoI1yIKxZ5l+oPDted4c
CH3Tx/19zJa6xrCJMeVx+nXab3zpyhgX+BBANNEYRCULWFowXTzNpQjFAJWDeSoxgy5pE5pQpRDk
z+Lh6SqQ8enRTOWUDYISbcodaDuN86bxL+L80xzcaNDggkhVJEyG73MBZmB5oLo06JPA7hjodCIo
bner2eovyo3RSnWOO0q4TM0+LUcoBjEYqPi4CHCYsale81hcXeY40Ob0WZl/iwQdlfY3D2L5oCVJ
mnRYSIWSIrQPulJD6mbM6BheFrcKRdGXEYin4y+UcPveVi08/wHsT/0zmHdIQFhe3ErioelRcpJd
lndRZ0ZG3XWGKSs+DfH3j6tKdvUZKFTJMhOJVC/rvhRPnpJzPWDu8qKrWebo3Qea3wBtHYvRDv18
QTVko/7nDrX6kxb6SO7WZDhbYAJqLp95EQpS+3Ui3AlL2d9BIdR1fk8CC5OyKIkdSPRc+v4LxUNZ
nwPLcgk+j7yt5HKHmmkslDHGsyO4zMG5lr3UZh5aGm7Koer8pnio7z03g70KCmm0qorfNZZ2Ub/f
kMPqg2k0M/DOKSiVJBRVdHefprl5nlLOWufiCQe0n4Crv7UPhbIU5RJThiWjpyrFE3pNhdDH1FNA
Lj+19fiOtuUrO+4WlROVt2skA6T3/7o/f1jnTkbmF4Eyf/hgx0HOuPjguP5P7G+FXZKOm5Q17Hpb
ANOPDLTHV9j5VzBlrFcEdOKcpF1mJ54uh2UZn5icvSYEE9TMlpHSqZVhSIVtq08ofb7Pe/JgpV/T
E2KVuTZpfIt2KJuN53Jgspr6GEWS/0HxoaPbesSnh9IdPn/UmEQQPSRa7Atjr4w5ZMR9uJXmxBIN
mji4HJX64JmHOWneujku0vb2ERb0aTp8qgkEATgymzycuJMwDLuaqqSSKT0G64iqngEEgP/puA9I
l+jKwoYZ/AoPQqkVamWr8sjjMHtVQYZ38Q9O5b4otaRFmI4fUZfgLRYebSs+AdIUUrV9zf4YmErx
A09ZbFlCBriuVW4lP5kI+UN0hOJ7iFg7B/NATGr7RsjSsvrJJUQqrydX4/ZzKOYwdOdYSO6/NaZ1
rop7j+02jANwXby6o6PDjW9no5HifLCiEdbGvsb0UT6AQTHxGT/UNd/kZYENXZLq6b6b5hFadnXQ
VF2ax82Hzo39g6WLG/7q+xjnzV9Sh4ZtAa4P2VuMj7Qm85A85a5wFXJdRpTzdBzCy3jXZgVlx2k0
26BD+QwnAvf0fJ8yRxUzYivRIBkVsO7EZLq6i/EjTsElyBn+c/U2oft968PUaqZ4R50uCs6PDyUY
CfY7/ZLiRrrD+D9BxQdbhbhoXr/d1oef3XbIiKFnYQHavWRwnlUFS7TVge47md8zqQSot7XcGuIP
N89iECqmJTRBFroP2fCFJS0ORJ5bgpLd198NIrDltAwcDI8CtHyaxG37yY82M6v7RvQvBM9+Z7VZ
Tz1EnnxbE/KUgh3xuK/7VEdkAbM43pzbnxrPhQl7keF1vKiGYgVynVCYwzzSjoe2F7ER66KLdiG0
jQnrJ+gNomyMwlPKaY0Ao7+36Vv9Tq1zjU4JjXOwKzqdibiBhSNJ6MxL0Vzk/XOF8HQ8bsW4pw7G
vP6ljEXmwlZbAo7R3qUTakOSqlBF478ZzgXwujc0VYa8qBaRRDvs5GSqmouKNmmdOGFVLbcuUt/x
mWQ0OcMXCwMIMWGomGKn5KwP1R2aWH9TcrrvTBWmNzEWcCfqLhvZy+zRx7R6xhio/wcScTp0TUHb
KPDDhqH5q8+vIpVYqwmwIGa1///pJkUch7IoDBuO4YwGbZklHhkK40UKLSWcZCx5UzQOAhwxwdFb
MoWn2mxv9bE3o+kgzx1tNPoAEhxEovuHgqFZVftKbMVc8scYFXoYlO5yAzd9LK5JyQyWvJbWF+zc
L6fmOP0Suzj/fJXwPYrAJ7xSQ8Jg3ehnQaThgZ16z3NFCswGzMxFmkJUyFTZOLg7/4CA5Gk876J5
RktUyfk5jLkaiyLoQNtsah38teaNCO07IXYpVj8Sfxm2CQIZE5JWQFg6m+PAKcqalX1mcekuLqaY
YMbcjOlVW7azYSf5YOCo1n7P8f3i5wDb1Y6EyaiDhJtadNQObWa3xHBW8z2R8JfH+gnKVNKvnsOe
e9gl7r0uE+bFOC1Eyb7o126E2rF3X4QHpukiZq9MVw8ltAVYMfzecpwMDhPwpRdxdmf/hMqF7PAp
nhB9kZ4Qt7v6T/xdBE0H5X0f3sTXjRVeqzMej//cSHGA4YqlKAIZRCGDznPC3AKd165ms20qWGsP
l1P2BUfj0hugp2ErMialpxPFBc2QJ1EQXey09WFOMFZHtgf3qqd/VOTVolwWgvfPQcGPVy+hxrjm
ycuZr/7p5bFNrgveyxQDxv9BbX3COWqKfgzFHgOcl9uqomvSQ/ieuclgHrOvUoLS2njYw0b26uA8
uRyp6+iYHZUUxPL2kbGIa6g/FyUXUm6/gnTz2FYg1oOGfOg9/cxq1bYiHExt5ketF+pLj/058wxo
fdbB5/1oSy3qKOrXZ36n1aUeHHfoiJKJpkwzPo/NYszAAMirVgL7GkfMFpJ3Vf4LrJfEvYUxUXvs
2MQMqcELUOGySDd450DjJOSNhKeF03iqPHETY+cbYevrzl53RKlLrR7PZE1i1l0EntEf2Hhu2bAZ
9r2pLCUuOQOo9lGpAo8iX803Nm0ieRHWk5cynzx7SVhIJm5CFR5E3PCbM1baqmDjC5GMdscZC4Ix
fuWtVx2xj7rAVfaWsCAwwMbMeyrlVMCKncVXS7H+tKs/9r884KgtG8uuiIyswF65zJCOAuiFbYwB
6dCAXM1+xxL84IV9n7xlupbUMa+wTopaAZCa1s/Tq/ngyBwrUCDPFYK6WJefEzU070VtGkDd5jjB
p1YMKvqv0WvreRhYojsdPlInXCMYeL527c1Lw2wTujQQCjZlCXNXb90yZdkBCNBXvjOBdKyprhEK
6jC3YtxNlH52auH0O/L0h/F9sBdLnqiJPUXcR4WckQDx+jgPc0MxX5DAqTsj3NheierrXwvdq/Uz
jXEifG/Xx71UWFkkYRLJ2fqURQCef0clwhO080IehpUu0zYHCZ0BivvrqKW5IcxUy/1l6+iM6jA7
tOr79oqv2j+Z8suworAmwUKsBfmFTJi69dMYTfoF7hWktSVZKIhWeqs1NKL2ScAZXpubb9nwfN4P
1Qd9XHIAqA+anBqW4SA4sBAY+55ScboBF/7Bv0nlw6UR/2m94nrwf4k6+gu9Msbv/4Ui6E33D8Nz
lo0rwQFuebJg7DCGheqYcZNBUgUNfFw81Q7dS5wkjPVEQMpVC3JBhEHdeM9pLFg12ByIZtVCjP0C
04qWyU6Dj57gyc2B6dVGcuRdO0CINrTKjwPLTsikS8anrf2i6MiDWHADVcDpfLcN+cMnTiSNeO+a
MeNiN6kF8O4lBKkDLDRUfFB9XDE0PXqCItbCgHxb8XyE/+8/HHN6ZbkDXbEVaE3lMuupF/ZSzfGl
/kPEk4IGF2IsA0a8VKPndB3d4yWxLcQ1FC8OKahofJqfZApzX9TAqTqJnb03L2LYUXH2oeKwbCmy
IZZhkJxo6mVdk0qiHR6pS28AOtrMgB53YY9y7blYEUTA8m914fsRqO6HapbDo/Ai1vVCZkYtGDka
H0D9s7OLlQLWdoQu1yIE0A7Pm2/1jXtIJ1XWW+OVmRb7N7pgFnUtU98Zpl3xnfwAU2ck2MSu2Gqr
+TMOOycW6XbvnlI+Bym9lt37IzBZYL0iy5VckMayxrRw9PU8tU1lNtKSwvQkmSlkh2QAtiabczsN
jkbfleHb1psrPkYqod20b3Ld0kOyBw9J0LDxw1/k7UDxIGM4Gslfb4OHCBJ5IeU2cYQ8JTDYNC7u
h70jSRLGjElnYQJ6DFcPPRXDpHGLgtn9qysAL66vjBdKlvXHRTpVQiL/4genD2NI+Q6xJZjdSmKH
EhVDzX/ZiSa0o6hLRr2QHLof8uU08HNQvSPVMgDilVYvdo0Ykn8pbrIcwU/FLFF2EJTTZRAWAgv7
Ft99u4bzl+gUfOK9gv6IA1DnSbbnyKsW/yOXTAzpig6KDho7lHX88d4zkstJi9ey7tz/VJr2ehbP
tx6aofIlcDNxtaGdOeQq8fqPIjy5JECD0PZp2U9ZQBYN9oGbtK8VXGlJ82qNuYEpGxi0Ws659Mt6
0m7V9bWE5usltE2MEOTJPj4Y2hQWSabLiNL2WWKCur2LYucx536XA3WX611Y8n2numO04U/IiaJS
AerS0VYSW2Pxr8wX8j7eiarHSXVx1J6sYC5UwmY4JJImCHmKsJ5/0FclkWX81njyT7vUUVDgJzCe
aHYJt12iJAD7iz2ojlcCGRG5k7kJpgUZJSaJQ/7ugwVZpFtB36TyndTodJECR+KeL9fab2rAFqAe
JjYod+uOrkBOw1YrUUSHmLd7z5b5zsP+jzcosCKFpbEDn/5zsSigry7DlJDdSnhfZdvOgg8HpTf/
w1t/vbgscAShFq7B4voaQPy4CcJirISo7pHUxHe1//ZFNt8fkkds1AbPZZjoF7p8b1C506oGI+a8
cNW0lAzxmPFo0iXhNfzR6iPtHs0ACQjL3zHp5wTJ92rvcdUcwj+BtiTK0WrN8ASVKIo4bsI7Jt8u
1syYsxSdLPAdcT6yAGntkDp0tmSG9ogJmNlEJnq9mPIUk86BX5iyQPwhBJHYCHxvOOA/yGoIuAjv
8aCb+6ZeB9gjdFsGUQ0phLa4WIz0MSkahEqmQ+u9je/uj+ucgMl3tfOjlvIDcyOe3+xfuRNraGAL
SIabSVVB92w1LWDqtWxgrf9H3ewJlDIgW29VMq12V5ven9C80ji7tn7EQwD9UX+r3mom1HXI/XaD
lV/Lu1x57IES0Em713pUnoIsU6zv2p3oxHsyK0YugFipsp+EFXKx9tcTRgTny1QQgUhaniKv7W0y
hv3CQh2GekoijxkCb0hXmlgMlUZLnBc6gFfIiMmgrTPAVUaRx/jQkXAVayTZWwPeAcB9XLfHnR52
Rvk6kMIzyZmsF0XaaT8O1ZNBm2L3p3KZ7wPs1A5fW0AZDDWzq384Gc4rBuQm/qQTBgCAYkstnA78
L1ufmC6zU+NvVR7d/yXLmYEZCWrIypHm4W78PMD4LBYqHQlIcxAdjIi8+MDFOaSb7rl0S2rZLUGe
TAphu0hI4imefUe+nA740+Pvc4PtwsRmIBH996QLIekVNpyp/MZUbDBETPzK/AzfMa2QkansHQJw
dpuFDre1HKBArTgwdtiF6tYIIPJguVXEioZT30yHa7EI5qmk2V4jNJkwntkOxymSVEipVi2OOy1m
FOxNdx95o2SDK3v7vi9TMdKx3HaUhyUWfUSy/dUjkgVL5Yey8n7GJQfaM7Go/P4tGmcxi7PUUZXY
jkqhMs30Pwtkn+w8NYSa0bQUsVfbXoMJqk915Tn4UHPAW73HhvbhkaoV6JQA95r5WhqO+8Lg+r4Z
nuHnTcGUbxaBQ+8oq7wWeFt0JuOK/90GOVt29gaGftB+ePvsugRtkEj1CcjTAQboEY1v028Lvght
SRKdXxoxWoG2nP0TbjtMKCuVS3+lI28gJjkdfK7TZ9DW2GgSGJm24KjX1bpFhMq6gdc78pDonZAP
jULZaRpL0otwU3UmkcTtsZ8SM5J3w5NXKYj0WTZ0dwIfA2Qtbotl9R6J+xdgbZ+pe49kmPWvV0AC
SU7MpOcTwO4XcwuOtErVhgsVD7yM99VEyiOaYaa1LYUA14vpo/305mm0lUfqq1iricAUtw6iYPfN
4uplaxk8M45Y8O4YVgR83LqR4xCDGSQfv4c2iRuoAlxQYca2y3VE2+BxGxWdY4instNIftZLlYSB
8xx7R+CSFVFa/F9PlTu9yojmkvKM2nzUCuoh5/DXKFrsAVXbK18YKoOd6PFsBfdUZbpRCIaHmvI2
eTyblmbQS2gYo2J+RumDIRLHOoYG7sYR0Ku/ywjGzQHRDHccJoxE8hL2lGUp9P1xz8qjwLp3TfcB
4vb9L5L6I7WOQ8a3HsnO/TSvGlJlNcDfSVXlZbBRdL59pOnSoIYiKrUkTRKutyGo4EMhMdbAuAh1
JfYetW7Nic5GKr7ot15rkr2ZzkH8p7utO/kN6UHINIpTouS11OziqXohLL1rmbclnGso2FyaISUT
iGytJn/jCUo2gvsgD+xsqRumOHUaXACQdWpR5S9m4pEn/sG4TBSVBZKIova7JFEOZCDsXXpunIMJ
KYsTcLXWnGo44+gH5Jr/z1P1FCh9U7vAN1Ek0uF4mLWj9jOtb+Os6tJlJEddgpeI86vIoZuZ0gfG
bina9uiQQlKTmEDSNMMiZJyLTdbR6jLvUs5gIoannLEGccKUz+ZbDhFx13D8X3NaMSMZzbCnTs6q
dAz07ucWPM+W7ALl+RA7f8MeLR8Z6j6gUaMVV2gD5yA1w468ET1NCrz9tpHKGEijTwB1TtS+Un/S
5aZHiVJTjGJgsX5C35TgCD1u8pTroQ2rav17ZckpVzdmaDbi4u/R1dB7Az/Z5BwEelQ9YQoCOxhk
hH37Gei+xBOrk+l01jiiTj+P3E4JGpDq+ZjYMt/4faZKR0KZWw7dlCdt7Y+LpJ/pxEryd3t0onoq
75hfrmF+fzzGtrRdn8Nuwe2IBvDlZEPFMvF+soP6eK471ubIokpQ1du3Syx/6jvEcs2FaWarhRaR
8xqnx1y5liFd0HK6k3GoIjR0CCbSZ+faP9rVp9qgA70UBkY8UWsbvYC6EPnJJPA6BwuHmC1FRWeu
DQVN0gM8Yd7U2toVYLcGizpwpFiqdwByXpM7K327jBO8uyADUGbdanIaZ0S8N7RXbw5dkFdOSvTU
BkeTl57lmAfY3jhu4Odz5I+flWPajHSfpXt6/ouBbpO0RlenAuG+oUjXYsLjQGNvArcpeaCws9OO
Qqe6X+vpxzxfvq1siLJ6KLfSV6CrSPa001Xl0l0sKamPP+Hm9/MPtQ0Ha3r4x5zIe2/9P6AfvZa+
cWgha2U2bnBoACqzq1OOw0cuhYytDF/dRnh7TCgtEBarUNryXbOMN1b6HVGQo2+uyHbfhuA2mpFB
S3IWOzGQWmnJby+Kwv3G7Nbpwq5zj1ti0iJI6UvH94oq7/zc530/uwnCZkhF1YTzB2exirrlexu3
Wd/88BhBf2SJ0BXvpTam3NBS34IphvxvC7awZGljWhnUJib3UdIgbOzaXN8hT/fVwG3CGHWWxGKF
7PYbNvYwykHZX/lARXt5q995OtuxfOjx75UrcjJU85+rpqF1DbzqFlWDuqY23ons30TpT/ntBWNr
UP0UOwxFs/h8qjO28TNulgUZ82Hrjpxp3vIy+tXE/FeHozkn4Uv0lojIxT64lOnTxnYTDpj6IEHg
k7gCXq3JLmEVfWlWHyx/snUd+qc5qxhGYQGQK5FstbObkfmhWco1vItjq4gyfE+mJzOnyNNpfq1W
dhseexkAxgMjg6sbL8baASlOgYUVK+veod9a1CAAJpISQlNcLwAgDbqFYDJWvTZmOVa7VzvG5ttr
sbPKgyIl5CDCP4IQ/mOtTxy3CgLNsOxQWa2K8cFQq/vrNohprrzt9XCkWgt4c2wDkskOuZ96hnZV
QYVPEJOv+9EDRgiNEiP9NgxrXhTalLBH/fc9XngbkbA855k2cgOC1IXHJOC5F2mhO/FzNhR4pAD+
AIawZbHEQY/vZbfBZHAdXd5NxMceatCWBd2Y5sD0Ht7srOJxDzJL7loLoGW2Gfo9kXebLZ3uYP06
rB4N9nijz39ilqAWAjjuwjFpmazOQua8n85HI3AnwQMg0yKp6XCZsPJ8hONdT5cYGwQawdSVFuum
VIVzm4LhNrrMGepLCJSkzPnfczRe3REUtr+CQlTX6VVE619cZo/1yo0/k1zW0XJief5UfV0g3qIF
DiAfs2Wu4J1CXU01y7KVCe41rtgXzHO25mJF+/VH6sRU0CXSkifc3BpoKfHtVmPZcO832o8X+rs3
jVH86gVJqKAVKvUBfFDkFCCcROiLlOp1vvXs5wilryp2S98HcX0LFWYpc6veaxuIlxq1ct8kcZms
/NI87rl780C1tgHuDlTVs5I23V28vWD7SGNdPWkJbCg+zAYaciLU0IFWxAj9RV5M1Ch+lB71Kfdz
fn+ijyd9P0JeuarjLVgSFC+QJ8n+ivmAjLB8K1JuW6Du7DhsR0swIq/opJn00KvKNbbfHr4LZZqz
dr7x0jn+4M9Jt84A8gKcfrXmKwOwoHl1As3CeUkQc08VgMGJXb1ZLL+55OIbtDmjDubmL7rPV4lm
Lqs/HsqL36EtADojog/cxaLQKHVu0OjbHaPlgPphX4711UclK9xzo/asR54cgBe8/kOSfg502lZ+
BwDZHDOkafzGAcodwm/Z5wfxX8HfLKj0U3VTF27j73PCZFd23iaXf4XJq8y+vNVtmv2aGI4r2S1p
YiBlQazO+cZZdo/MZXu8AQOP/fFqAiVTDuuwxnMU3oynJxnL3Fjuo9BAHZwoPowxES2dfNKoaevQ
BlNElTUhHVzS1+HZLxWOESg66iDamt5LAcpTHICSrBQUR50r80cdcgcRE83N9ll1yYo42yWxAF+O
pRWUx1sT+KCO295td1h8tPYrn6lK4uQ4EVVCAkVdcPHLbGfpACI+tJKHyPzo4Ue7qhPohW22Dxfw
HZkDFs7Zvc6CVWP9yzv0iOEsVCMMt2ssmp3RM8ECXZu/wltza7KnNaQXSCVceJDoqsGTMK54f1pH
v+obTUe4mVr8cZOg9OlRlL6Pa3YhaqNCieQ0VZOoAW8pnsbkupfAIlt9f6hfi7jU41JrKoEKN5X+
rdvi4WGO6eEKp4Z5oAKC7Teq10ctSiK6AJx2ceROAjTXf9pVDsU/MUQBTIDrr7hjNBnmM+5AkJOf
PMfSBv1piopxetFWjcQ3fmjONsuyA+3uyyXdwuueojaoTD4kMkzgNYs/hO35t8c8xK5siOirlA9m
nWgNQNX9QnuHLb4qq8Ly6oPIYYMBLzuwQphNAOBlTio3NxVH1/7XAO3QzjwpeIAt9LsI9Igp7kQc
vl16DMVR7xObpIxouzTzMXE5rsYcsexjCU6AQsN1yucTI+3lB/4sBH+Pl2YxTLo3Ci0QjtxkvP0x
xS/tmMZr9INDkRaDAspMo4mzcfrjgO/V1f0VzG/Jlj0DnFcGU0IG8GWIkD8SehNwH8Koosg4eGUH
Q044cuDiSOxRE4/EI2359bovLyMPG8Ry/4Ds5dzjLg/ZECw7hAY6D7m4xc4mHx5nMjHrth3ir5j1
wzLhy6+XquhLlwt5Bbr+C9ES2QFF9tBUojbIXJO6NhJpRf5YOVv3JfrA1mk9wJejp03vHe3qHNzE
4fVlpehlaKxp7mvgn4Nq+DIb0Cr7e9/oUu86yz0j9K8bg/d5dbVBjgL+jQUPMaFEygGJGm7C/+YD
v0lnqRi2KX7OCM/ORe6kXtexEb0IOAqsEA6/t9kgoB9qtHU9+E606oWz3hfYR3GAu+bnPGirnbt6
+dc9zSw1cxUaX5sogOVo7+gKQdfF0IQVESlvY5H3lw1p7PUpd2uqKjTvy7CRiHywFflxeeRxJc4F
C+b+c9XET3oeR4H+cirWaL3Z2kEwoqbpKvg/eMVL/SL4IzKxWn2pDbnoP+xOLZpwGSq2AqKpeodx
KhWEXL6a4CvebFmw/kgeMtSZA8KnV9azqWux+uQ1QR20HUULQgXtCgw/JGUuGbnEBukyVaTxWMoc
vsLNO4ydlssJN8/QzVL/Hd74x9r90B77dhZJsIqKmeCZts9cHvyI4nJ5ZITfjdcNORUZH93xuTde
gvE3A4FEJTs76dFaVxvvLQNniLtpiGAR3rJprlNUIRrm5PnIOfwU/1zB5B3cZ9lVvF4ALrYgw7Vy
A1Td+daTQoXamf0eyv8kt4AhyV0eKvG24fpv+CwNzdnhRaA3gl+HmSSdnzGKfpUjUdYR09ACNya+
BcsExhtY/fJ3FQSz44GeXReT/Ap737ACY6GkqfSYg+eGh8URuT+S/UqFpDfz+gaaBli/WWQ4DKC+
Y8B+FbUY312GC8SNKmwqCznI/9Xg6g9siTjDBAwVoKi+29slaojPu6WFAywJX91GHHwlwt1+djfX
u1hG5jZLbyzm7DYAZ7ubvoJ+M2v1xuRPzzGA/rAQqVtwOpm7ibteZLBo2BJlnpgl4BlKkgu+sugJ
/zkRfQJfmI6He6JlDKRpAwp5B0HKx1ZlJ7N2fhbrtqm3/RmyjOuGxuG4wMYYH28eiGz53ZEEmXwl
YqwmiFvh/Cwhe9HWPtzQOCC6zTF2s1erxSR7NVszZ5y/r7jfP24D3zLQ/MRwK/cRIhdetPE5ASu7
WcklvZNMcC9ErK6rlwcdiO7/h7Nnz/YP1MlaBk7UuXM4Ji3UuJFr/X5LCOWMv+LJSs2Bau0yesUO
ss/d2Hqt7z0f4wcsvJlwNLWDOQfPfLcIFacMZuT2/itheQ+f5gPwUZT96ctuETNWRz5kWHk/ZNqV
QZhTJCD18KZJoGOgdVtaPGyy3XKfoR4r0ESaZw3ooxXRaYOeaXjbQRZ7qH1DKK8QDqtkoVZR7MXX
JuEvi11dFUPIbNXMcfEYKU408Ljl0b/2Me5oLneiyrFed+chj+3jWeF0i65FcflteohTgcfN810I
d/2bFK9F9jk2uzFYLD0D9LCVJ8MEGITZrtyGydHtFqW7HuALJHU2A2nMhfVNj74VEGpopqLa7s0P
2UPbXpJVp6q1E4DREDtTm2L1N3gh4a8wDSXDRRfdesWYMvdfnj4dB+SwQqadce0DZjUNji/Um6XH
zpssBIOubZ1VgW5R/qAEBTh3tGDcxqB7B/e/7EL3UErZZ1yvOYk8Z7IpCfgJ5P/0rrGExIRgoRYj
Rxfia4GU4AMDe8BkBXR0s8suX+wQR0Cwt2Y0gjeW65/uBMGdv58W78CsvsCtUUslX7xWijb2wHgj
K4sBE1krnlA1XvYg1WEnctuDnNJcMpo806CPuGEWKxF5EvFtw4HlTtTgUL5hbOu8EpTgJIwz8Jug
RLe9jUpwmY4kqRcKVIdck3KQHl8LmjeBnkiaEP3CDaO4iqSzZsW0nmvZJ8KR4sY3DyNzz3WVQIDc
YmnE0zNZbK5B8QhelTHfdkH2pDOa7xT2udbGuz7weVLAmg7REdTZgLzwmlg067yChDvkicCkLz6U
j477/tiQuKpj9lhh9Ltq5YjH3ASg/JOPRhtA+RJzeRvuKYoY5n73S3fhkT6WZWJXVIjluym2bP+F
zHsxKBlCwV7B4e5w0ODoZw4DF5Cel/Ku/jGKiGFVQa0MmzLk7j7WYziHmRCftaX4vYfS5WqU94YK
1pmimoXWF7ipzyp5SljHRwa17vXg0EqmqQsRTpOXfnKvj1sYAuGtfOnDwyavT/jOZepoQFGMmHOd
TO0+AOvps3R0EXyhbZy8DkIFIfaqiK63FCvirmtbGV1RwDB8/e1Oj4Ne4Sp9ZsZWH0lEHNTZ2J08
n2ARGG9j47ikSfxefSetY4ImbNdG/wUClxRiHWoXPgfGBcFEy9j4wEkt/gwMzoqEeZTYCzr2JEhG
I8DdEoPvL7CxYka5pGSTVLzdPqmzRDtKsOADrE6RRKcpcC48dbz2oOep5FDJhkvGkJEwfq0hJ5+X
F4nfPTmlEZooPmACkFPa90NYPfY9pQ7OvJF1gaivZvGnkgxEpKBinglfKh2tPQRvlCgW0A3VBWGS
gIIW7uNO5l92IVlie6mJZFOBCb/yYODbInKUb9Q346RcQeGcuZsMe1zJAm+g4pWtoVYrGNz1ZJda
m0PHt64G7qAq0CK52n7/jVAVewaD4xut5s4GkxGu5R6D4v4KcLac4XPXSE2ikHtgGh1FR5kNvvF9
qzv8oJazZV/hjYI+QIBw6yQTnf8NlIHFR42yXo1B0CNG6PbJBtMIDgGvzoOV1JOJQEdrH5m0nzzd
qOZU/QpxlXQG2jAeCDwEBSZ/Tdid9+149oLcE69J9+Jv36e2KPgjMY7Zt9N7y3XG7Nabt+Dp66Uq
K0ml5nb1nnuX7gOdz9p2eIHuAIC30bwDHxFGGEvef11fqEU49qfMtD8iHuR36ME4PewKM2bKagiH
p4PiZmuxF3NkGZKKvLVzRlKekVN42Yiu2km5UppfS/4vm79rWpyXwNaCuulOHx+6F+H32xGoWKgF
cot8jbZncByBbgUaWOjDQ0yQTxFlNo4gKJvg2bzZ75TskysDegZyLnOJl2pyNXLgovHRcs1KYV7B
wXOF0lkztKTMgkw0V1fkbdIkyx0BDM+2K+qMJod4fFhXZJDpXoQfzd65RyJu4VFHA/pdJXvZkvR7
Xb0L61/F8xuIVXD+nkwOUauTJRkH2ss+bFGndAFSZ+oSsgp3ZxJZ5MOBFV6InLXTNEG/9Qp/cwfb
WikunsTz1/SfVZPqkmCy02FckGbXmKD9dWx0Q+EguYmoub/CIl67kSA6bss5alTh/tvthKDm0NHO
Yz3N6CAlTnkmbb9S2l53W5E/xlaxLAcGWDGI9N5o/SgpzzV+XOvCqsOalTrhc2KO2HL5MAcUxXxI
A/Rvp3V0vYQ9vXryN2FmLGqvurjnzvb6si0UU7tmTJ84gcek4YeX0RDiH43NlolQhfjcs1R0RJBO
wjCHrNYrS7ecOeeN2AH7ssrAY0QVo8huDH+zFMAiQkoO8aWiGhzlKl7bBVZPUCW4bncRtcJrOBox
rKxVHJITiZ8nqjygFddvB/vEGo1/iGGgeUvW2SYlMjTiCooN2/Y1tPbKRnWee1noHBRXh0T3HEDb
zZS6KYEsqpWJTbuO7iHV+Bwz0vcDQQKPR9DcTLCK5YOWDmF/iucR080VpcsSqz0KI1Di/sXXBk9q
OUgD4L8Uvbv7qvrde8bK0hUHVFn20LJyLC7Cj2qFb1sWmRYbYc09xeTF+K3XEnZfheQypg656RMH
zVsZIZUQL8cXFnRnHXrtC3AmiKRN8fEbkyKIujzwxypz2S2Wt9tlksOCWS0NFcZq/jw+xj+rCIzH
QZ3Ly1FsIx0fkuM1T1pcXawwrZvf7Q7QC/uw/6WWAOgNxefAFvrAfFa/t74a2dn4pDMY9nrwi9cS
9+z4pq0ADHWpqJ3nW12+x/oma1qvAKCDVOS5+0YspgFqrCjvIrOdGJLLrioIFXm9kJbGRlP7HYs+
ONLALK74txJqTCc79cMCFMWVaUp41zrDGA974WH4oUmVJku1xNSWm3Es8AoaXpqnoNNofbgJYM24
60QsRSHNQmZsPiqPpeOxT4t/3SPhdFki3l/Glsnj9zKY31ZHLBklla2N+v6NKIoGRmzmFLNtqhoI
iiI4yH/9/gaXYTU2kOa4mirZHN117J5mnY4m9iucrusFdYBIzVVmUfjY3aEKz84b0EqEqhAZZIwG
f4otdPAIzLKIkGnfbi38qXAZCqwCRymcbYafoXZ+X17UpD+FxL1iVBD2NdWb1KnAorIWxhMTOLr1
n17I6I3QSUL0obiqfoga1GPevP3c+X8wiD0YFcuTdsigmyKU8NuIdjHfkU5ah6fqdY+JeBos0BHw
uvgmFs3I+Y9jOy6IhxrR7/cqPYt1eWeZvWYenQyzHXCXFeNGM03El9XYTk8wWEUOUg/C1w/It+XS
1XDqRGtpTJXmiIbw9tfg++yZUlDphjEL5G3R4dOQFHs6PlQcpayYbbL1rM+Y92rZC5WyQ2k8ugiJ
dLmUCp/oVdeVA/rx/SNb2OkJBmXmJQya60IuQTEzKMFwyNKFVOqGPN4q8i+5m9wIbXUVLMTPJQm4
+EnNgqvoBoj0qr9wpw3SV5AH0v/4sfMuC9U0PnguFxzoLwPnP4cu0KHugQ9RVC5OIC3jxTkOrezk
e6B4j+Eawn3XxR/y9GkQsPyEl0PHDGTeSQbCmS8Tqs6kobbO5xiIoS+55WFcr/+DExugOu1XzDbB
4SJABvk0cXVhVeQJaTHz1iZcMlJky6wSgVbpzSg9unN4ri6SilB8Jy6Bzgi6jd1SQGhSMj3nSaiT
uxNU+Gcr2srhYmhycMl6TLO9vR33+vZD0eM/NRjd8+IwTXecJHVkff0HRI5R0oxghDJiICCp8JVE
YuKFvQ49ut7PK8qTOtGB/y4rt04RyNsEOT93TnIxWCsvALyFnH9gv+8PXF8x6GXnn3v4dPCfIUlb
XTJgFIvCD5Vq/KBMLZJTBLIGjpo7Z0l0pgkuj1IwqRRHyo+TdjZb07zRB1on0x/sQ2fo7WrU/fEj
/BMCaQeG0l8xfWQ89LZUYsvEe7qaMOT51GpOmXG5djE4qyMH2bWOezt+ZXPHqHoIGQsHEf9lxD5g
qVYZe1LXcMt9vDq+cIZ+g5EQ57Hby69yDefDAAcWjxUMDW0KBQABIBPaaWgmpDulbXpj+qJkBnSn
+2rjv8Atxt0vs+dSacv6tY+6cJhF1CYwdUsx3vpmYRp3Qni7h0oKQLjkdUDRCCtYsGSi4JJXbdKx
8Me943NhmJU/w7OtUVCu5nY3unRM3K38EsRJx30HhvDx3BN/xAcN+7c8iMyeL0q2dK9+7DLKhMFZ
sQ1l17JdQ5B7LJDQW7VDirdhlE+iLCMniNFMu4XnYhp7nG5Jd9jPwvxuW+sR8573PnTxJcDiqYkm
vdNDSU50hqlbzMj0kUWwTOjXesdHO/hogfYKamY1bodiVuisAMqDJUBNVUIEHzx3RBxGD7lloWvV
DD/RqlvDEqa7AhkLnbbeLvwqtlHzLiLgzWZh2czI8N1KBFGLE03lwvhlnpVuxjmrVmxGsSqrWbEg
GC/LOSSYCREU0UtNlRt+Zcia4TzFwmmTXhJsq2XS+WpNWsE04dttbtzIlQqfKXM4KxnJXML6HDXM
PzKrI4x0jdGaKpjgLDGSD722ry+1aCgkLxkqx5oT9C1z4xYfqev5Nc+3klGv9hiecE5SuYdEspFJ
1oVVpx0YWlCfwNAsraGAHeXeVW51J1/eFZzGcZUPBU9hGJovl6p0X1haMeCVKlFgWRv61FNTuLdz
6V4yEpblihDrMiLVFMmHBJvDH+T7ENLebrYH951leozzR6ZNVfoARI8zMdyw3zliuyDf+EZz2odb
9K9NL7tsDg0Os+a/8kcZvOb4iLSlHdydVmgWMnnMYJw4f1V78t3L9NVSfvc5oZ7ADEmrw5Vz2/DR
R4vfxlKvmUwmXQVhc+kfXkk82U61kOVPk+5iBhEUpcz4rAh6pRd39h3Z7xPAxFkKuooUqaA/TKSy
do+sX/821OpttxpFtJbhspwO16foiigYY2qiUWLxatvn7zJM7qRa6IBCBpKuyekM2Zw1bcZoskLx
K9Bek4nQn4ycsP1Hz6pVdjw2uU8EbAhNCDWp42fiPLMUmf4eMk/zOdiP/c9KtDI/V5iZIAd9XB5w
RKGaxGNPo5UMyJ7X1iX7w0kjGjjGwBX0BAdYqoDVc2F7OdCDrOwNm8jDGEjblNXNFG+bJY+mB1dG
POru4qglxfeWpoHkgE0bFafBkvryHv7tXM/wqgF0+fXdZ5YjtB2w3ad6iEZTH+3iEs3cI7gBfxMn
p+rYp2Oarmxiy4PGiM2TyBlEFl/wAKfM69KaHpSSTI5uGZpANIuvTvt6uUxb6oGpr7Saz5Y0GYjU
av+MQz2JZCX7EgaG8mx83b4mdXVOMyU3N+VNhjeED8/kEVtYGn/ewmfoiQ70tPdWtQOHUJju3hC1
CFjrBpLnErsdQ9oYGFoVUnwbXILEGVv+HNbGaJw9OicZK7K3Flr/qGPXC8joFac4ErQrUES3jqun
zrvleOQ3/rlvMCGMgDv+rGEpTIRL3wqgveW7fxR0cmCyzQLkwbl+P7E0dK9eR0qLt1kslN6vWycH
zQIRk/JxXbfPYlzR6graDUijB7vumRiUA9Lr68KOX+5IEeGz2fvdi1doLtAQzcVGCGP5rofnkWSZ
VwyholGPm7a5l7tfoAZdDrrN7pdWFjB9L+X9vqxuXndR9fZAbkBFlpgD4to6GZXywCYVmdPcikQr
kcxUHliPqI4oQ/FFItmrjgmU3l5DW0tYoxrzl5/P1kmL+Y4Al0zZrxiv3t2iaLyZsgegdqNJPrhN
hFMbRBOQA3FxG1kFLStTAD8RGLSbphFw03SzPd/fXju01dIidlNBFI3UglawCHgiSbdy/rcA6JxI
R92WA4h/jH83ElKOgOSBbM8idYW/0Q7HXz5ICOgei5uyKM9/JSXpw9Dugww6/z0Ah0R6sZwzPDO6
o7ftBncmCzKYItniFThIiN79GOuMJXv/PLDFCxw3xgR6/z4bj4j9dpawL88PGWS5IssauilOGkcd
vnxR38IrhAU4fRbkJj7vqXQQgO1ItJ/UPIuq49rsttKYYm75zvpT8isGcGAzxUeW7xUxVcQpxAbp
yPHpMHWwdUqUg3PIe0IEQfk9V0fB+jAhLugADkuCzf8yI0eq7db05muqYgw7SGnvYRHfuT01AOCS
4lrLPNhfvUzyp1LPucvclthIOUiraKGgrF6PEhrJemPTBICNR71EJtvGBmrL8i1tMLG7qSg3Ahf5
cJiUmlOQRazVsFCev7ZM68lA0XQOzLFT5TXzWknYcFCFE2Wn9geWL9wBGRDWkCdpwoPxA7IPBRTe
2LOBplDB9DLX2Ks6ldVKRLMfUTqtekRpAwl3+JV8iCogErSANvoksA9iasy/vkWPAPJA0EuFpgFk
5MRHAcJfxTx+PcG6+/mMS2hQtVO4zg4L0Jgxw6ckPZpG78THu1QzRbA6UVv6OyjpRRQw3itdVHX0
VnI1EYWaFiL8L2fejiMUoodol2OAYtV0nbsLOt+zEVtxhCW4ybkTP+xyePSJhsEBjLizhg7+HJZZ
0l8DzxpSw3d2qkkI69mff0YKcRXmToQ5v2YxT+iZr/UsGaPiSbimzaMQnpMpSvBDdGM+NnUynZne
eZ9gFo6B2mpNT8D56gRLwj51xlQ+zraxPMXQiKmW/Kq5qG/sWllSeSH6JshSvaGmNPQ8Y0g3Lx9I
6DhivnJjm0nPy/KhECwBWvoSdh9MH779LKJ5Q7nFM1LVzAMkyJoHymSVzaUZdfDOl5BBmB/6J1Kx
LzyCF6JmylwKHMySrKMIzpk9h2d3kyrPF0oxy0FjhAdTplmZAs88xiyZVv0xEHbpiJzKtx943zDI
3fFwhIOk2jfjdbbZCuVDPlSIAn/2DhZxtu9jeD1NLQkR2elbhIqpLBlOKxvp/9ywFAiZslGdFQrG
7Vh/fymxiLHzO1U9NPHrUGLhM3LH/YQn+HonI+05Dq4J35l3h+Ou/Lu1KUnD6oZ62+yEfotFH2KJ
P/k7ymNqvv5nspTThARip52MNkiJVWJEGvDqeGZcan7/DSsVrYQ/dyzE9s/QUhV8tur7o/qzbZ6S
8uCPU5cGy/e4xSwKD9pcEMp8kUeg/QsSLVdyLgx7I0UDBfz9XooJ6obJlzojvglMjpbYU29GWo4h
HtspRiA1AtwXbpg2g4TXgf6ymgxdfpFp9hpmhXHnFVsQ5P1zuOItzmzErCQvP+m2nlRbXW3qUAu4
JawcE0zVpiJguolKlLSjRGZLb/jiUaDW1cZR75KfIbgjM572+oy3LmeRxtf8vWWw6UOniv8L2w1O
nA1OGoRoZQ0Sm8Dm716VrpXES9aSnrZsX7FdncB3Z9KJLbmMKQ105eLMYLK0wSwvbitdxLKdpX2O
HPd702UXs68hXZeQxYtplF1Elt5dZ8GpXCK17Svy5b37AMyyq1WYBlL4Bh3tcCCv0fKBNtRbBxxw
egyU9lpeU8NzRebn/68G1mkLnP3rRkwl89fJh4p0vz7gfV2FH5FtcFz695MlJvX0dwIoaAFtLu8Y
FCJHCXih8wjftwPRN1J1d8kdcESDGQztXCI/NJkxNYStYsYZk/kSKZZ/dJA84i+qVlfNaauoLw4V
zNJ1wa141W4OYHN1CBdFnfQuMRXoWNQiCx4Xs5V2XYZxdkHTNPTmQJUCXggtPxyKiPE/RMlnIsqU
7bM08Uu8AQTIBFuye/PWu9RctlqyA68WzO9ZJkDNBE2JcdflKELkFt7H1c1nxgAM+fIDOcU9xckx
J/XhEN9vlEMCYxL+RekKCUmd90+/qXxid8m+a+GVLfsO/tNc/tULoMltF+ntlXLpEPzkM5bbPmCg
ml/aVVd3gEfF5GHlwCcDcxUlofjY+JWA3mtiATtfY1nKjliLasa1JjTbcC1Brh+c18PL/mY/XiRj
zlbjjajXuaVR57WZ55/427431sw+EfMVetEbnmPqZVKr41VWZSntbx3w7umfmrCsWBvpqRM8L63B
7Fnh3l9iDAPfRKadGLsqE87AHmJUJNB/6LH7i9sbEQtS73zSMkoIv2j/73hqFcGcvNghF2p65YIh
QfN0S3h6rCa+Bqfnhj6EJbCilyXAvLlog2dBMu5DgkCoLcYrkFxAEqosjw2CS/HTEjOmmehV1Wp0
tUQkGnF9BqE5bp9+2usmYvfyBeAd2vBR0MH5dfiXGa6hfNAOiMQdMU6Wr9/WziwsgD6knRsm1WW9
i4GfqLos+Rbpot7tBcF0NWUTwp6Ex9VJSPDpJwUJL8Dw+mmWLofW2fCxbrUkb22yIJyzXxL/RSVH
7T3sbOUpBpV7omNCI0euhAh1/6UJ/mFQZH2yI96KqPMK13twp19eAZG3QDEKcc+50DAYiRNAGWJQ
Y6c7HWxavyMFKzPlZEiioLOX+xHLmH6XxfTj5MTDG+FERh2ukmqFraclmAUlU8SZvWT37/8Wi+S9
kaHpbk4jHFREKR3IqtwS6rlCJqUqPbEOHpGGwqGAdfSyHwbqGPcGfGvovrwUviQgnhScuXT3qIRP
7U7QRZDDKrezwhmUvKt62S5JqyHOtID6cMWTyTms5Uh13Od+RbuTtgEjr+w84eEXCF2MSy6ym9sy
uLvC5XoUDjALJXZ/1LjSwX6SuhnDK9hH9ZLTDKmOhleOHmgWFIUP4to7hFYIyiotdrdMlvI4/p1l
oka1CHb2daHr5AK5MRX/X4WN2uoRglrfZ4O/jQQVGZFXXFpLO2j1V872FcZ0t1IOrjB+a3/q7aae
L57kqDvVIyr/SaHYsmh6rToRgRaZo5eIYAV0xkeR/T/MU89E33CLzYZeNsnl9EoC555mz1SvI0j1
iInAGFX8Z3jWviTR2kcTc1SC3oFrmQjFnwEOFLbgL4vqjXRFq3WEHz35AP3WZkquVd8rDJ+gNJaF
i7SljQQmb7mURXJjYmkmn6vw3JQfyYBd3mICSQ+tYIIcNiLPnItswoaTi3HJxwVCbg8QBDgoBlab
gb2TfEWfee+PZtFIJOAP7GN2bAUr5W+BBwLmSm8/Sjql/NV4KD4d5MOAiTmmb8gHRMqvJgs8eEmJ
jQdkiJ64dSnTFR9TanBlyKvcEoLucy6ScVeIIl8RGzoW8QyClx9QikV1v2Ie5rvWb06tzrAtcb81
aT1ym0KCcFzbLQ8O5IMLhoOgr2dIMemsA56taVJzClx1Hqf+CdjfkDu5LE1BKYUIsDwjpk26ORQA
3wlmuMJy5xNl5qRUsa2Fr0ylAiOq1rP5BKUZcAGAEz5tzCkjojZ16fShaaBuOR8QpLtJYfBJ8MWD
BxQK5Jqhbf5k1LQIzmxq1PIYVHorminDYYtU03jnFwQq03rdjAqQxFmBPpiEpC0wNCl7t4UjgsQr
TqoH4+pD5gby6dFBQuvstReMzeQ/Qp0XSP7rYal6/YNi2Tgb570ZgttIoK2CQddCkJ8PMmkXV0KO
URfCSsGoNZz3dDjuOQMAuffFDW0xheexIAyrxWq2/YyDt42P1OeTh4uI5iO26vB4If7PS9qCc4gq
F+0Obm6LHQdFo0R04NhPfFut1rmCoxMBsvFtbZ4j6Kzqngl0pQhSQyCTPw76CuVWLKUsGyOJjYPz
fezZ9FQ9voO6Ok1Rhy/rfBTO5xsgXRT2yF4Zx72W/856ptMlNms9eqGSPkTfVBKlASL8ov/iVsYQ
t/fuNY/YOymhHqMm9MVoCl3yseldNucdNrILU/j7yOPdOcdkHhLcilv/8qXYpx2jHj4a/J0sSFYd
ZemH1MF6YX/k1vqHZUzpJMfs1JIiPto63zTwfZTQrnHM5vdBQMkGiNttA47ASUoslt0ejFMANHAZ
nzZfTKjnDzpUThIPX9xmj9+RB/7XcTJBvwbQZbGX4URx8LFtfTJekuNrGuNfMvMsbgyFIDxzr8JM
M9bN14Il4I8PWzftEJXi9VczJCwHkcnEv7606wCSVsR94dE8RUemwyGPzEuL7V+EZmcSpCk6jDb1
7ojp/ebKJiX4we/+X8fmQpbnFS4LHRz1MdUZnP8xxEDNQEY/ERU77cA39lEPi5TrDgzw5uakzMat
Xpom52wxdqWfCQBu5ZPlR3I+BnUfbr9J59J76c+SnO2hDeGVDZ1Eo/Gi52bHpcsYDXhm+Sz0B1Xj
0e4WxrWDeOYgwBVQ6tpAKYZa1EesaDbtTxsdhgfzM39wohErJfA/Fbj64risgS0Kmnd0/o4CckSf
AiI2KplTfBovIyZPymUAS1YAVs2ZHDtsb2hGHx4zGzcG83XvcKT9haYBl/7wY0hrhVXMhlC06n0H
lPOHTfkn2T+ZSLKMuA8tq8nn9XY46F+BXHWNYIwC0ozWIlO6xAvpBgj4eRyZU0HEYAvQSLFvtdVk
v3LdmiEFgXGi2N2/SM5lTrhtw2dTj5ZuNGCZORkC7xzuEid8SiiGopKQOjKYaDeDEbRp2Nvw4vsU
mliCNIcCYbz9M5g/s8PhJcivKHrur/lY/dM6vLVjxolmANL5V1h6a+6i2VzZhKBdxelqf7zT8HGN
9vPKNC63kD0dgVS8g4DYFqyITfHbQN3npYEGyFIy9Fhx8OcWaLl4WUYeRWuJDJv+Py+n9inAQFMx
+UbaX9g8bV6XFSVQOF3CUBs1LEnaPOJdJX172VYp6Dlm0AyVAtfMAuxTIkAJ+tKiFs8jKKPorvlp
o3jGtGxrQvvwTFFHc1SoBu8SR8UO0ul4vHSDRPScKhe76AIgigSMJnhm+9IH5vaJzQEX66nZ9u6V
w+Od5k0uQsOBp3Ylq+ppx3Y03ER1S09Z/AadSnmXBIPYZR5+2zeuuKFe0ja+HYXWHoFuHGzEGkw/
rsMZ+d7QGOoBFsfvTL+Ur078Y/R0wngSnfDaItSfTz6quxwYvM1drhZADEt/Wtgnlu9qGusr6Hzd
FsuMONUwAYqNHFThi6txVAXRQ8tVShx6u2oQuYQwpnXF1NbX52jiDjJMgGgBjHHJO28j/e5aoWsC
KSBFHCMPkHaFU5F9tyHKoHNghXdAbLQ5N5e7m1/vT3A/DYBBn9TcQqKNP8m7qt6WhEmqw1sukudW
erqUpVHCOnZPWScP/LPAqqdNXV2v5+DkXZ7d7uVSJ2KNyDRwAXY6hMM1GJtywG1JTBqmFrRRl0zP
j4QE0iqykwFNqNUIf++Dg2zyqeavcOeHo0TmM1ImEnjuSkZ6++1F8j7CrUvm6DRm5X1pwrPN1MS7
eG213/OZJkMcEWmMMor9p2BIf0whoZpfWi63SqSA2D/ZyNM1qAD5/c47wI4h712BYjeAxW8O6+Mu
5Fa2dfrRSLOfhEyk39xZ3n6ElZuEQLTclzzPNENynykusnaQUDImGdw7yuikhQRuAEg3xPkaXXtU
1N1MAptAQNGPHbYCW2ZDdtyW+OWicLXvj7Ccfmd9H+3DGuAavpcNQ1ex5UU6XWW2YhcUnkNMeRIv
BgEE8oAFuVrANU622YlbGzb5GoinDb2pAMyw6UbVShlE7TFhJOGYgDaCO+Rguj9vnHKdKPTf4kwG
QTnxShbLiJI0Y8tSFa6cflKj8NTaMdxFUs7tJ8+S5yeFfd7xIU0mbLoDJ9WSHJuTtEKXkQ3jNtwF
V4GdMGpQCiHMGSvEeL79GVsF4USIudP38HFDWwmf5POQN9b1pEZu5zcITPUXLnZe0cagOpNTlS/O
tVoIqvs+/A4kcit8s0XccSlV/+i4wCKnhNyw+bYfxf5AhHmcGZY3S+X/jFtzMZRjRn5ztIaM/jqw
eSxJAXxvl0Dpt2xocDN0PEmdJe/fgKVz/OazkK2A1IZ4TEROjbumPWUtipyeiV57bHmSyW2VcC8s
btio4MDKCquJTlAVww0TX6imJeGHo8poJegZXA1evWkn6Eh/edz4DBQFXMGoaV+pEV8QtihRSrHm
rImuxQHhzI5Sx8tsEBNCl9yw2sOt2Ysz3VE827SRK3CNk4YZD38KVimyPa06xwFXT8uymGeoWXwY
dImRml8Ql0qQOoEHHGbdYEZCLmM3zj8nMUrmGS9uxv7YgKzDKWZ8PH0cs+PgunjQRU2Rzzc/5d8W
pFIE+7EofAzZxVWvqSFqB31RATog6oO2p5CBq6dD5n4tD7tdyHm48l1d2rx+1Y+V5LduLitCV5CW
A/T5okAMj2PbFOGsznk1OSnoi/RxjB3iFCNTMvo0WXK4lDbu7h8A9OczpHaaEm57548T4Ai78EHu
9NC2za2BQicYZJLlMF4o4/0BBU7WLn3Mwk0DQGvqOXw7N0/3UPlBoH/osdg5l/47sRyA8K/CmIm0
zPNmCa6gGj3+C39plzWEG4A6HpaU5levcR74Xj00paf5SkSzPZN2i1+xfTSon4pLdoGXoz1ul1iH
0b8+0vSe8Sdz6+RqSoVK7ExrEp6/wBYRGgYlziHgLmYS2e5bBjviK/TJvVOLS3XhERjddXc+1vFH
UJ6hsS4not9unDjr0qW/an2YHlvLcB672iiu/retGKjmCI7SQIndOzyGr8miZ5WR5PjPVqSbEN4f
lnd1KzGiGmvXuk6GCXGYucN6Jg7CrEX3CamTeEsTohq1VARzt/MaCkOkELCEmXAZQQBLyuTimkbx
ukwQmmh/V27TOsXsoGOMxWu/c6baez+xFSjnmjNtQbHj4B+Xj9d1FzwbSKPfa69B+qLiTGpGMT0F
xaxdG+8HrleOBHjuG8gMYWxWvjK+yg46vIo44b8Oftrbac3ryCjZ/eaS6JZf+SGUnTbrz8hv6BjD
WwEX883oJsex8+TUF3Q0+YcFd9otxVH8JWY//IHjVRp4V2zNWGGpGBWZ3b9NTy9vYOU8CZj8vP3K
TpVRWFwqMB/wcT/jojIpQ2H/odWZvmlPZXNwW69GZwnS+m4z9ZcoGoMb85IB0j8g5PZ1eNHI1pcN
esuowNuG+FqofxUNXxbTMtgdUQsyGpyTDumj3nx1HmlMoL2sh2wP/5Cq9PTSRtGSKR9FQ9hSdmGD
pDAFxbYng+OFqjBOiqMmD4s47rBrv06clIHl5l6HsOJvaAQRf1yxQF+Rg+H+v2o3j158Xxxc/Qeh
CXyYMnnTEzicMlnkejFj1a2V47iDWpIIDhnoWv/AY5fjpTfNJlTOU9Qed1BiAiMZA6H1lVFlKahn
D5xUGPBKqzDio1/EGz8zaES1avCdpVJ+fgsTMKTQ9NkSGQDPN3uBRSn/FLjAcqzESwPa6Tjy9/kY
H0Zi9jBpIso+xpzteU4hBT+C++z+sb1nEOCn9fejmx8Y5xZ61FZvoSW+rzidgpngKDCQOA0PXlAo
wSEiq7DhAoyvL3RE+E8Ewn3dHlUGAjbNG9ubFA2R3rDwu2xIf+Svy4ebPWe3pz/yRId17gmetPC9
yyxzGRIBomF78wu2xI8u//MqWDugw3cqLLAC+zPQKP5hfDp62wroRPaZSHW4U3KgyTuDVGV9Doqv
CfSfTXJp3tE2rZFZIbABqh6y96R7+ydQBp+Fqjxb0MnuDme66/iV7mbZOsygV6nhmdQBxU1hNcLl
38d5TpdSzmSXh4o+T83e07gFsibtDewK2KA3cDrb4m0A3b/9xvLxLy9eBYS4okLRINDrGv0XHM4M
hbPWcaz6puOcatfuDnAPPDIcO50+H8iaiZB7GsV990lT57PGCYnsTS/GOhb8TogpoaHZbsMFLkPx
H+1eSXwj8DwIKeTHOyhEYWzeJ2WiJWjRzbGW4+oi596swmBV4QRURj6TFgoDzv6qnKKZXXd4gwc1
ybIB8ABxkeFPmDEiUvHGend7gqthBscBeYuS7zpoOk8NWd+yE3IMMuiM1kMeLhY34gWiwWXN8KW2
R77T/YwzsXcRsmYwzWpozSpZYMPo9lXYt64BqzSE+IJy2lSByMXcrqKu/kMXrp5LbTisDMO5xozb
fUBTgS3ABaDb0KJkArTOmFf5vxsmGwTDRrYq/GM6v+qnWGnK5dPoQ2xmKsEyvgQK73hJnyhwcvAn
K/RXuma1OdBfh3aRwABsPywOpGlfm1KIoYjtPjnoB855cmeOQWWdNFDl/leFPzMgvRMEDt+rhqWU
5LlM8t4x+bxEpQi6WF4UnunoWt/aiTE8N5tbUTK04LUCCfd1TxOj/ewvZpXkIOlZCqgEi5JogMnX
HKimMuGAatJgm8BdrgLp/b6zQWIV9k5jS/hlTbwjdbdMj7DILkmUbjm5IwmdpfXgyrxquKuTWTyv
apDs3/uPsB4CQFUO7kDrYfIILMUihZWfAtRJD2uF3Y4jgoeBRo6i2QuSsH3BEmrDEhmjRxNrJWDx
ZiQboPjCaGNNtrbn0sfCyfJW1fyG485bwPSfnYbxDeCEEcNmE6uK11hkwOCo93Ohs79M7QSS+Ruz
fcxinR3pfD3Ih62X+jpXiKUOr9iTARf58TMEzZsmAF5qrifBB8vjTPh9JdYdLZm1zTLuTsocVgV6
SgCYiWd5U/lM8pnR8YbhDk3LSfWB0gJCJTx3PBTNXopgjtQB/yKh8EHBpmPOuxAKOsVfBQVG//b+
OpcONpBmevrPFmy3d1LiobccXsSs/1Wp2U6g8Fk2x/EsRDYcGQWtQ2Cm5gP/7refUqKitf2yJlRA
xu/z0DB1cpEz3LVJ+OAEkgVF6Qu3LutYCCmIWxy13KGhZLRBeiQCPHQxdbBTSYbDdzW7Os2wUjJb
bczfvsu3rSU//BoHt+Zp98OBgBDRv+NPaxq0MoVigtnlBRvMVovOUj+3dtzU71Q291PdOxhvPyBY
ttBsVrEzfpwr5/EkcEv8czT+wC3KUrDPDabOsKLZsIwvastz4xuSWqjDxsCxFf2iPhx7IzjJccyr
X1LtufZFY4zMtS9ek24Ay76Dd5dqD7A0fVYz8d3Zlr4fEZbp32enhs30NYvXFNLBCzeAk+wzT7KH
hMEjHDLy6J4rRi7L+QW4FNGV1KyPLbUhR0m60wUqS2I6za4uqZC7VrdgmMPQogi0cWUmr0AULMP0
S45eeiGQ/cOWupacX2JN9CmOA3K3aZcdvjS121kzqZCXKFFTHlyzPPprChAdX/UNEd6mug0wtfZO
lalIiw7LEWCYfxfwJ1IIhpC2TsM+Cfqv4SXI8tq2PE18p78TJLs+oOQurQIzoO2ajMy7p4kLp/hs
WoWJJHdWFSISZ8r1XjhDWvhflc3av4B9ZhgEYUY4V6i10uvUb5BWliAEDQJRjEsfDn71aEtI18De
UJNO8D5oSZ4anPEgook8z+ACMubW51/BoH2Ptj1qa8syimm6tVM84ymm7zabgMxAA2u5pDR8GowK
IVBMxWt0NLSPnmNLZtOiF0OXP812Ex7C9HFt18mKz8lFI/UkrCEXDWlYwCdma7cwJS9QcmvaUx37
eqIiwmpF4ZpVouJBOXE2GcRTRwZWHKimEOIV6bzLq5aY99800m1QvVOrf41JLj7eSfeyfUvW8I+b
hHWw7VbGwXJAvBXn+J3YDg9nQaF11ZfRl6YDe1Pldk2uM6N+eFhR5a2EyJ8Q8GXjTs9BNIk9JyuI
gq2ktzEImDauUfCFgv7l84YKFnmyYie7l19EO2RjIJaFq8s08kBQPLSiNoeNTDUzib44VQkLeHzf
stVRycvIKgbay8a/nEprLblpS+BvAuOVMBSmatnNuS15GMRU3SYARmPGd81NdlsciCi0ioEDESeD
L7a8lNP17Udq50u6RdZZNtQ7zzoz2+d8+alYutilpNjzOybxoXU8Cb287GgNrBlZrJwQHBKHopXb
nsSkej/I+d80nc/N+PAAr5znjxl6VAqVUDup6VIeo299SkZ1giLpJY/MNb9N4KyKjY3ym4o+dovy
uzsVWXNP7OmZ/0Fwp0gvVQo+IvYVAUOZfaXGcIX2RAhVIj783oUYdWGDduKZCxFjbmScwSdlIf7c
TLD3UyVesqG+GSHUyyIgYmc4OKvuO6/UEQzq5PJMsYEkomNYolmEglvM53cnhtaCSbDYhqYf6Tw7
T9ZBnioo070dRriPIJOWPoZ3fEbB6vLZNHJtJkn4+k3bzQwagcTU6/4IwPEIXLoXpLycj9QwRVC7
XN2MmQRprEZckC6S3xIefm/1sxoL/mNOH4kzS8sPpnJco4BXtOlPqbqOn8eGGV2hGRZQh0fGr+n4
dHVS3JI6q1TGN1/W7S0EP8qTMcnGlcxsmrcWHl9NI4spywTg9fELjDogNOZqjDB3oarU65fzeHp5
9PNbanj6SY0qFZDxhMoOBdrlH4ts2602UyhBBjYks6/PNJuRDOdHbUhOMnfkX5uwpD3G/q9It9JA
mdxtdSHEAOXz7NQBpCRC8PaD66ggyfEacMwqHEXj9cQkVLKEXrWx5qnfI4U13dxz26AxCTDE6qtP
cCmdcZLV5adrI1sazahczmiRTm/z7CURVya+1UC3UETonrI10qUXK5cXZsEpGDKY2//T0Q+CFqbH
V0szEBXZgAo7taR+mPvWJjdcEarToyHowfU240Bfwd9sBZdv+sJhwLOkLq9P8DZXHFLA4/ktw+Pe
tv52llHhoJawWntvPLgdWM/cmQL0DDcgLzw7Z1Lw2lSInHWe22QckM8RWTuLdzhRU5mnJJrspgu0
iWMmyO/RFKxFrbgGHZbl1+fj9KwQ+xVTkSpgu/D04TUak9QUCx0V/CNPMTTixOLSGLNmCUVz9KKu
iuFP+9gi3b8/Qd5EG1DxOtPpVjBYqmB6TM9aZGC5FkSbNRzcAeKFe+YhvStTUOnEhAn51sDEXhCI
2BN72Rw3LV2uEGomnCmvJVVweWzIjU/iyhye2NJqmd+3zHCoh0SpRf5OrdGemNLZDTSzukx+DRLf
O3bLEnRRy5Aq1zZEOpwbndO0uzE2fGvRJkpOyFhv8m2ZKiF2zg+rwhBpsyOFeAThuF0nXbAtyzts
bgX8Z3yPUsMBP3h0LyXm+wRAvcFfWviSkD5LrubFej0xXNDEes5HlGMoAupAo9WoWhlD29iO24Fa
ZtvTelRv3wUIjcpVwMVEzo/3NQU0Gdgn+U7WwR3212HYQgvf15pVCMKQ5ksSz6nqU344NlZfmkz4
rV9tO2esF3/WyITrd8zXR/p5CNWvz3ofiQ+nh4jVLISoMBP/MAKxtux69EgHl8jrpow2fRyL+ABX
h+nIBcR6nETX1dbWysB17UII/a9Yo2+6FVP6aN2py0meM1VxEvNYX96Dh76Sjr3poEtORYYCXkdG
wdXxnjQYEgiia3kmTlSNwr2VMB07RqWf4lYwvzCakAcUZsLC/p8anZfURUKBMYdNlHvsosjLKvZ+
4UbRsJWYO0sob83vGcoYOWm+yAQZ2xY3Au0Fl74dopAWwKBoU3NLzka0O2/2WB/NegT1PrUU1EZR
SCbJb+3+GvTJKTLZZrbWgeilkCBpgAjlVi1jiD6rF+wgG+nSmPwfaXel7/Jz21OZrtBayInTt540
9RLpVOYbo0BXK4QghLQOFIUGuNPwgs9Tq+kd4PqxluTr1UBkpB4BaznICCHT+e3yM8gPKyihCv1M
1i6vdih040kTBecDGXs3HxCmsYarENZS0SjyX/jj04EVTyL/Tb+TIvzSAL58qI224sQaryi2hZ3N
CEbRZ7cIqHlAx+iC1alhZE2MsunaW41CLwWY37z2Repgc30M4WIskgAwtR62o2d4dtelRetrC3Ov
xK1FNz11n5+5GVZtkgUaCMvYFiHkRUy6t9uo20tAC92eQkU4SDNPKjH3zT1kSxMPw5lGHyjY0NHr
2ZVU4Omfaq2TzzIBXdW5FdSut9x4NMyMWL39Bc2l7g5jPYb/pzSVoANqKT97AvB0HXFKQDCAx9Tb
/CrezfPNqvYcmGsz9WJcA8h7qaUxVluXapUOqnGViqa9l7YXmziFnSaw/U0Xcf1TwhKPWdqj6krC
zmFY2dyDqVu8HODOdkmXT4zvnKcHFHntTUypxYaoQ5yrh26eFHQcWV9RVI0U7VdlzAVwtcLWXOPW
OEY0SakfTTO3mQPshY80d0uJ2Tmo4tIIVsummN8tzLBuXDUgjEA9N4b6n3inz99Z4DWEmQAblu3K
tiHyJ6YE2eqFt+5LDE6DpR0JDXmHIHkw/VT9+1oael4UFBeoRlCsoguG6qfjKyZeQ/C0pkCHriXm
ytTEy9Sst9CApeigUrvK8boZeyabsLZQYIrgnAPDzQhZKxfh0oUdU24mgA5HfT/ge6+qPQrmVMCf
gRv7thPH0AKwsnXKeNCHQvDb8s/MqyeBXEiLUyqUAh5HYzLycwCOHHczVSjAqLnsCJYvg0boCQkJ
00Gsmk/1yQYBV5ye9LWnQeajhPksbOoHRg4HToVtHnodbgaysoaljKQ5KpZRzF7LoO5f0zfrVBwK
zo4zr27tDZsoXgLhcPImDobRBuibiuk6GcBPtbzFFbb4Kq1+uA02EpM/NNxGdvzmpEnhVRIS3RSR
sEjNvWqinYbVWGGV22rBzz3eiAaLqP015/tjwSJbQZLZ1VG6U1G/N2JKHtMJEuzkeUPixKMfc4Uz
iURXIY6NUJ2BnmvgeBtKpKsYLv3disDnenXBYJXEZCgwN1JNzjKYlPAmy7REtckSvU4EVYOwn2Kk
3xkhIJIZtEy1B8PZQsCyh7c3LPMVw2fVxrWjLIg6NKmsXTxJYdL9wRes7iTOwPmR94Z+oouPoOsa
DXmYnZDDLrusd/CR/RtxWq9otWg9UzyqDR03jE5ahgqCMGjepMAQCLDn1OSt48LcXJQyZl+cheK8
5QwU4E+j/yIkBvD3yXIk6DYEAelfpc1BO2Yhkf/m2Bhb8AXFZejlB6iLP3ifgIiiQptTw5yuSf1v
Tbbvpc4OaJul22Vk2les57ySs4raOduoBkP7n9lByQRS/EVFvyjY5Fx2rf/0x/sNuNSLsaKtnr1M
XD7wNBvrlDLF8qEEeNVS9ouuBJfdfNrTeC1KDqoXCRPh744HQlmv3bmyLlqcQm+F/5hFwFpWPU1O
D8s7vJWGxcEw3xZCy1sH3sZAocNT+LXxIPs8Wdayv+c8DxCmi7Zff5KVFc0uLzQ/qEr6rQjCAna4
rdFBQqtdJ87JNno/IbgxsuFfmKqLzJHvcZvFXc1ZNPheCeQpX79NlOBzj3NOYyQDHHTgA/7vux34
ZFv3Vo8oBt79A1Sm/Say8U3fq5SjuID0DSpfy15WB5qu2OJlWbnWwB/fAl7PwYpxqtf7rDuTMIIE
3QNIe7nUjmRTlEdtKenpf9tFHtdHIitWo8NQdeJmrBcRzkbxSjhQCGzO/EiJ5x8xSJJDZoUDNNit
70LTVPKRjLciy7N5q4WBLIEkY7+bq/4ijySuj9Z9hKGhuTtig9OBCeaep3mr+Nkj6uZgdCZhQ2jA
j9MkzorNqWxUa0gvp+YFS9OncFMSjMAYjaAbz288ZRVHrraLUfx3IOTQAkwl+T5gbZNoeS9sOEHm
idm0Lm6vOpBMH8wKq+0URZBJYPkH5C7VnrbzyC/ZeYkZdAJZUkQdhLHJ6yqWuayUEjQpwyV8OKQL
dxLZJMbK0/eJpRUM1TH1xvI2JsId+bMZAwMUaX4hHzXTo7YqLLWVK2WijVOYInRq/DcMoQwkSPt8
0UfHx3RPfgffVS38SX5kYqpQqqAe4PwBOZGOTQSV3UCLIpb1ZjlSZQWDqCWgl3cPHjHHyJ2Y0dTE
BB1zt2Rw7vmoAeDBURGVwJcdD0pD+1mazL3tXco1HGtRKhFNbs4rZc9y7gc+2HVRLhO5q67QB6Eb
P1nOHzq5rGlQmOKIaSlSrImCF8r/b53YeOdz40HDyCuwVJHP3NZFUgfVvZrEN/y6kFgIMGNVVQTv
pOkDnE93OPvRr+EoHJR8BL7EJdtVV5HDItAKGtWQ7h4+47aO0Xd+imPpgfyRtAYsK3KmDGcxg9x8
/nfGUtiPVSxv+EXmOAYLmWIi4m722ofzN8SEhjoalngiDEhS5KslJdvzLU/t7IccXQLVP8pB9ouk
qCDrSH8j+6tJ9j/vAadBWUlC0NdBuRFX11QzGs2/ZwyNqJJL5ZTqbhB2BPekUHxvy5Uu50g6tqTr
3Z/KJxSg6j9eUKhacY7Ylb4NuPCQZs0t+cwCUW3ePVmhXGW0CBJnlSJxt8dqn9eQ/CBr6h1C2CdZ
leMRlfoYUuwWDTqq396zkXZoX9bpaMThvoG81nqzwhnHYR4s6eWNx4mkGst+kZ4ON7dUowYBZTQF
cTAlphxEAVPnUQjknbztoI1l//mrG1aLythsBx3qMl3oQ6vyD1NI5hWuh1psZJmbRas23hIBCv7/
sSv/SJV0VJ5oi3ouxri36UKMrn1HSXB8K4+uOZaiJmhC1FiO+u+NVT+rZMiG7xgb1K2Bn+scDbuM
kpsgHJr1Fijzv6U0U2K15srtJkjjJQLtaLmOtWgqEEvtXznyzELQpMR6lAMDoPu/DjdHzVo6Mnf8
pfqN+0QsBLZuIEiwmKemCXxzltYf/rPwcAWNJGJNXmif210nEmJ/la9aJNq1QW7SviBSbVYK4Nrg
EBbtKouREY8pnzDTTVC06gO8B+XXXQikGy/DaR9YpWnZl4tFaJh2dGjZmQPsG1g92HqT+TiR2Az5
mYtDFtJxEXu2+HVSxaivwCFZZeezSiCxb9d0kOFxC7twWc9W+JBWfO+26d/1O+NaDVE2fBdhU8l1
8jVJ0ZjzZPMFCBAHgK0kr2lI1PCshJfSuZpzFyfspmWmnqjVl+qUTM8CAiac3yqnaidKnGWfI2uc
tuV+R9GIvAbpxLz1k2aqGpM8neX3ly68Y7TqD96oFQSrsLXNMALfIP3aV3vNXBzaEiuGENqEILOe
btIPbhlsMfd4WNKlDhnTcdSipSLMV+HosxDNeCi3f2Oc673+b021hxHDFvc3Qc8Au8X1Quq7vkW5
IZkXzZro72LlDLOwX8fdG30xNAUCVZl0w7lV50TslYpe3UvlvbSlKyKh1T3i285Hj4wDM/W+BPXr
lobk5V4NydqQ1NBWVSCpb6kTwtm6dOSFdbki+xe9PKtsy//1ROSfOEe/e4z9M2AEqxVaid3p8SUo
Y45gfY3HIQkMdeT36eVbljYzL624So4vakFqdleGWrFqEV30nUy2l24yA/t2KT3qX+Vmc4fHmpCx
ZFoC0xVfRZj23vXwsiw6Sz+kRFd4UDhFMcQECEJscWSehnOidOLgt7UG87F6yN5Q94OO0+TV5vk6
j/yeifpmVSmgSo7p8sA34mwudyot25Hng5JKegcu6N2QdHlsjRWYufUkzBX/YfBeqmi899Scmdrp
HNfqt1mT0tFk5TFc4pg8gtuIBAId9BbtIurP0TKZoV73XaZy4O6XsD/SSsU5bb4oriTgZ2dHomu0
ATVQplSn5qVJdWElfni7p+OcRG93S0Bo+lxzMRpYv0GwLmkAiKvqnAxP056BZ36ddZ8sz3GGhTGJ
h7VdtCsIdttZF1EdcPMHtlKkHjUOi8ewFDZh0pddRKQbsPG5id1JX1zvzs3btL7uJDyM54Grk1qy
xGlwSqUuBYhk9heWWb+yKWAdmsV9mwvglklO6uNSfaH1w8e2Dq9x7LRmbXL5mxgjpUb0aPhh2Fpc
Kn6zYTHkxrn3WQQLqBX/nOA+TLA8nFGCdlwiAvl1yIaRQjUSE1bSF6jF4WaGIah4PGcwb/9EZXgN
SSrlHNJKqIg5GDVKNjgzd5zPNbzIeKIDGZ+W5HH9A0hqbKvE/h0/8JkknJInAVFslQxh8oUx9TnU
ezilgCXvniX7YRNpYYXRdY/g4ynu2A3ZXMnYG7UIMOkTIp4j9CJ5wrarVzuXKf6HCMduVRLvTRd+
9LtioExfumTaWucuQ1HGy0EoHNCGDMIVwYis9Ins/QzEEpa+t1XB5JUhl/tii8R5UEShfDduJmB/
P9CvtPMZpYYRgtBPRcqUzHl93q/vXBTa/fZ3OBvMaXtCApUSrcvwSyMbo0OkHBuT4rukiqI7uBfB
ePMz20BDMkJtUzr1oFYflFHRqhztZm1/HDD2DhOQckKoiM9iPmEQx1F4yM5+1BybJ34Zt0q9s8J6
f+pDLcrcqeW1/yXjRf4FiZqoeWqRp1b+E7h8kKcW6Z5+88jfwsMW3/lT0tfDHdJIXB5JqFgVUvAt
qBdCQI2L3whsnEK1H1PYGyTQELPilPa52fndKYhjoySWCTAOKTs3Ru1OZDmn03DQnnJ8IWNYpd50
k2+CSIriGmFH/0uAZAUP4n9WWz1+WkTc/xpUQ39rFgSXHf+zZrHJF6sBmW3yGVeat3VAd0GcSivi
lRFwZx8u3v+Akkzce+lc2mpCM8vH+8KFIcwFfc1eIwIAZnlV/uHLCKiXm2G0sWQqp/+++C9vPylL
zONniCPK2XEPrKAkBPqKzrOP7WwDxZg3rQdldxasdfeX2r9f3aNkf5aeBv9kXfJG/UiRgHZxhX6q
140oJYgBFXtTgpbIbIc6b4K0hYbEeZ52SMqkQaRKm6q4OpMS1JTiiGop21l0mL8soCaSAM+7So2L
EJMUCMttHX5x74233nkWYH7ncZz3B9fymq1vC1g/obTQ6LkweaOvI4yoI10L6ADP2P4U6o31Xifu
d2wxnr/IXLFzMZm/Vmixz4qciPJ0I+pPEBVWf0Hrx3Wnvlk34Ma5OCEEcsIIpdKrkZOmaWLL0zmO
ho079/WKL9ORm1S28xsSduaidoElUQ5U+YmrccnD+3sxqRv7AXUs/9ARnotXGJ5gLlovUMYwLwee
regESyx8vvu+YW3Wze1mBY1kcE2dvaFb2zlLGVaNXvC9MPwohND9/KmyQ5GUVlA2JCqz5mwdZc+N
L4Rt1mfthlzWdvQ3E9HDIfeK0ojMYjIdbU0WSvddmf8EOfcJHgdlzDK6lkpjF7yp+lMLjU0XSBZZ
+nE/YO0arid4FRY9uxIM4tfiscoltMcbDNUIyK/vZlzSkQvUn1q2H9Wcra6oUvBKC7SgYMGLWJI/
j8umPtZOPc5HJLNXImfw6AwPK5RZUHC/w7qNKTWkcA+G1IUjt5uthSK3dL6VDynPjKjPY69gFr9s
cSDdZPdJRBD9/9z/ZVqTS0hIsIBM+D/2F7ikNptF456dareJjH+QbGzdrPDH67q2ki35bdLn6lJt
MVOK3lrVHTXJa0VZEyr2/ikEKZh7pCRmb0EXcSh/g7wc1INE8wsi4+onhyDKsdU5XRb863+L98j6
kSMvEGANWx8XS2z6bSatRsq0dVitMJPo4AD9z98OknYUJyA9Ys2n+R0i6uqF6WQ/WnHphStvsaqb
YGVmCbZ4F+DS+FNFk+DXtSpldOvd1XSmH4RdzscpqZfwSSZKQ7PhNMEvHkQin94BpF0meKmxl4mi
IS6LehtyNwGLirOt59zURkcUOqPZm3BbiHRwE1HHue3MkMNyPh+SfTBhuZT75VYWkbSwe9S2iQUx
SQLanZvdODCk8fUbmGX2kA51ChbUt5LpFgiBtnBpj+URLEfNXwt9/LyUb8etfprw6XsUEAiNqUqz
yvj9WuOdTA1oHpd8Fx8yFCcgODgi7/L+cHYBBMsNnk/MTBNf6nf8lfQKMA0+VqpwxW+OezFCWBVr
LAFRtHJvV/scQIIIMyXMOf2oqB8N3u/KBrusbzLAlUlYyHX2w8eXNX6aHs5o8ttusW69m83iN6KA
fGkVnUkghZ5WkdVOy9izJT4cd1ZXM8dwwBb2EGM3qrt3XK/GAOWQXtJ96SBCbtgty/KupBHbST4V
34ca5t+9s0dU4X6xT5Apo570ho6VteNsGyeaXuN8t39lSmUqQuRpS8gjc1p9MNcvBJMM1Q8HfeJt
8cpsNq1NnZ7v5QZ0sZ8rAGmUcntaiQ/WkVVyet7MksFERunZGHJu7Lnf5z+0CzsC3DkHEOd3lLE1
ZRmgzxJTOB1dK1wL8Jht8sPjChgSGrVAxGsDx4ZkRgE9jjbr6XdvqCbWGhUdU4aFmyGfuln2SmJD
+wztF/8AwX12lHzoeXjSsBoGnq4blFJgmO9JPrVbhWdIQRi016EvlKMJ+hlUyHorITbC/XyaCJdO
bI0+lgBigUyOeKAOu/WVlDC33axSuhogzUmorduostHeqQJE3Y3/trVhO/bh3enkyaCX7MTEP18V
5rK1MuU2BJ0I1q3pdqf9tXhfvof3MX2YxFNDAs7K0yT0Gofuh6QIV6aEbPDDhEiL4O4fP5nlVj0O
xHPNmlqbg4TwvN4RJO4eAMMgTD/81Y6g1wA8UlJJcMHfZp4z1C0A9YGyI3cnOGOJtLveXDk422Hl
Gzpxuva8E6IY5EU43nfJ0hpNdSWQauCM1811HRDDJyCoBjeMGt5i1Ds4Oow8uvRvzAubyS3duMnn
vl9FO7H5hdNKdzghOlMxRGD9M8CTOhxEDVuwMUMvJEdAlC08DWwxhyS0eGRDpZhE7P5B2IYhh/u/
MnHhXzmqhq4XDZD7y2Jn1omswcMG9RZ9EbXIL3hruqnBxQo8GI8Es+DKezeB7vobRjpeHApUy/vZ
1g9wWYaQ7FEVzPBCSCDTZJHyXyAhEEQ0I/EkPaMwUZlZY4LQN17ewqxFBNq+u1h7EPdLB5BG4X6N
zpwRO6qw3fBlsZ8ZjP5oPNGxOOXWZCyE1/vEK1yR6Wge/Poc0dGXxDX2p7pQjFakweUReGfeLFGE
fd6R5IhKmcHPG/VBBz840ChZPQ4ubpO/uEi+2jLN/aOz5NDG5mWrW+fBzKjj5/F3t+CXVnFYsmks
qtG0o4wQcnuGSYZR3HRJDRDAA8JwIR82VQ1deQgBDFEfinZtIZEaefyNi/0gOzX7r2iXlGPfY9o9
GWvytdrsEo/4F0vnBfrr4artUvPF7w+vfjlIEbofokfgz+kX/FrBVKBm8CNEfZ5LMxTorUr36ZAO
pqMtKq+mD5xm8awk8yWDT14KUCiOUoKzuzwcyxaefohgRv6p98sRHnbkSN1xhf5dtrJxLTXRPj3D
rNooItB5YJbM4gpDp/sxKOZAiy17Mt1sC/DC6ksKiKAk5/3L8Lw08dnhuzQp+7Ubd+4bICrKTZIV
AH83USsRIfXTsi2N3ozmfIZI4qUGJRamajRI5VLYU9ApkIDXyCgkTYlho8Y8rIh94fdNXqApNIDW
7JMbjoxWPdGr0CkhYF+5kHjmkMrqjHmNjS0ErvQhyy+WppFDjOShJjBy3QUKNPGYPmQnXwaFQjqa
5AwExFqgb7uGNvLkHGheNw4Oq5unAvCaRRJpkx+w4uLPxp9yM5GtJZFV7TdyzFBQRbO7BGTSie+u
BEksjYlRLOz8ivW/EXUcEewwyH2/V2hDPHwAIX/QimDgT7RwItHjrifLg+bwF1+6dpPjTCrTAasV
O97w+cC2o845qPsQ1IGhrwco5xtapDpUkyzu5qQT9lUo3H0Hns5+1XSsoA+JKV0vvQ/TK7jdSqXx
T89Wohe3VIi6tYgcombCGLJyjLD86gpirvsPDZX8StHy0noi4T2DcvI3efdRc0TzqhIOBm/QvzIW
m4kYaPT7bndQJ5l+f/qiP+QKYSCgZ640ILP3nkl5WYjZlrW7BCu+ZuWeCRUDPaFWAigG3onqNIjj
dKLI8RM47xuJ4gvBvBxoCrauDwhsw+V3YcFnvNylGnRXpkYV2bklIe0/M5JtkOsfHw2hbMp2aFI5
pyj/0fH2WaowJwLLtSbPF76E4tfDrA7p+6CHXpHVwP7itXU4TLvgPZlyicfdw0Tdjn3RGzQCGrV/
npMnGWkomSuGnfs/HaMhkbfaTOv45Rl3rYV1Fa1yw/iogPTWOrWD/BZyzt5Nb17YrgqiDq2cb/T4
i4raT9ZurKPz4lSJ1GjX1imd/b+yxum1z7Umz7+DRgITkkEJI2jCxhj7J/LT8VVKIjiY8gzsuBs/
UsYlHEIpcKrcbR+n8w++a95VkfkpgdISsXXFvvtlJAlcNpkDdAABH4QM2mbav22un6Ge0mY43IBK
GHJ9fMcqkebAu0IbY8dzG14DEyZ8V2A+hM3FvmmNDr5wUWeZDhvBLWUyOgUsCEjJli9d/0XYRpxN
L0MTjkgsIG0PmiXrAhBU+nU+zw/FFcQqP+fvV0jXe0E581bgZIFuuALHieXUSgkvse9hR4E5I9mM
fiflLYzL7eCH4uqUtoT9xuJ1EZ6fiAI4C1Is1zECGXGYuzV5NMfM9wA18TIJP3xluy0OLiQu6WEH
GuzRihGpUMzno/I3NfjxTESnVh+P4WqOo6aChjZdvD/uRzCg4YIaS37zcfarj9B/YXzc2u/tTYId
IkGKHROFoyxx5jiWK1jYUXpiaT+oadk71KK4tn7nQ9jC6ZC0KnS9G79EUvSabwzSaZszGvb0JSwi
Q/fS4o7TYo+Mdax5IJJxY38zyyRYfJj3293uMcYHxDJy/6aWFGfndtB3voJRIfZGrmH0h3w0B+8k
GOj5bgkJtt6zMpIu9efGJrLE1EaLf/C1S8TVA8/u3c6WdYcx59bBZyf3IsaHR5CCtSD+rcQjkvJR
sP2UX98B0CMUy7sgOdrU5UiAmHNnSIWCOuc48t4InxIZ4Pbwde2c3gVwVYo5AbiucUPd53CsBcQO
pS4/gZSJAY4NuNPOa9ky5pgLDtyatyeOCtCvYIupbJGmTZcBEHW0AFMXFKgjVrMag73AA+QfMiST
+Aoj5PVgQDgl/Suc9zva17r7/0nIs/auTEdkW9VOeQcCDQfV3QEFQmn09sinfVFjKaO/ouCjlJo0
hONhxUV0ljV+3S+1I++yRneCCRzvI/LlhdKT+SlCW9G4chBwr20buDiTp6CSKMaes/9ZcMA0OWbr
9KjNvn4UeF96OMj8ZGFMdsQXZdCADA3Ba3IjhjuQGci0nHiT35rLZkALTyZmbA+vSrNmaTMsfxvq
jZ2g5awp3BYmrgj41IsLf+H4cXgYCLSX+MlVUeXCzr23+wTzLguh/rv2VA3r/A9goRvzDKq6ePzY
aHStiWz5Al8+2Fhx6efotblQRWx+0IdzYbeHTuXbueOAWfE2U+EBbemZonqyFR0HCQVC0ebuNle1
UQtvufhsNtC2MLKPWyYCDQo0Uw0rMxiFkaEOZ+eA6bmYqsKWoVK1XK7J69VJEOvMMAqCg5p3eJG+
14Vm5sDpsm+a2IUbxEs7QanhxvG47hCl2Tezk7PI/6xzSstEeUyD57v115e+0FQhVWUZ1eaA/IsB
9A0jQgs7lBa/1v4kCyTIpw63CmJztvcRcDI2+9RjomVFo5VccLtWHUsAuu4O2m41U212LHXXr0uo
vYeQLcUpgDpNZ5pJGW4nivLO+kqmMWpQ3krJxPw0li5yWgbo/n5nGXUHjQyoXpuTSZTYvXyiOKF6
dqvQqtY91yNfTzPTIerIvhAQ9Ah/xaD159IaTq095RnGoj3JnJ67vs/505P3ni/4pupQ7hG7LeYr
/P9AYQ8DMaYSM2bD906yTFpVEH9sZYA2DMnQIiI+VBF8MnBeCzEsEUZOMJTXMeklV1HHC5oocUc4
e6gYGhvCZvPIEJ9CIsmm19WKmDx0x8tJVGVbCnPeVUZozCQ5S9343I2fKl3qXfIDdScvnsV463g8
F0n5Txvrs+VNusj5QwhPsfJmpuBf78sAwJuZ4Smujo0aBhLAKciXj1w7MLfLnv+oIsHzLF0pnptY
Z0R0pwguyjK7eMFnhGeLwGbtTZlpvA8Zg9jFpkpuHZd2ah6VEqCXAsWkEkJV9RGkWph03VChlhmS
G7Xa/xNuCCqQOyFRh3HmLt6Jzgv8orNyyXU4w4imSQQLwf22P0Lnfoa25J1N4IBXsgUf72QuWRA4
FE4WLYT2jrrxFFfDtcyVHF+ZWZZ5N9drcYmJzO5zgX1KHumKTBqg0lmyjoKNQ3HqfPvqCPd5YD9Z
NO+8ZJiL6RYzDSo6ZcsSA6QceSV62/p5ArRrt86vwW8sRbEE4uNFqgN6/xTlBEqmUP8mJofc/nr3
0SM66BQAfkfRs+PgVqEhW80MlV7wQiUYzo9KNTmJg1/dJDZLE/xIOqQmJg3/t7aZy/XA6y4LAFgS
huExz9cFnzYeU9Llt6XOpnJ3yFcprDbwS/vYpp2uPRqwPHz8U8RFc4wCPx3h22aQ5Y9NaRZT2pnT
JS7JvZMoCq06aw8XRcrzE/pQjvO8dTx4pt/wVgx4Pg2bQkZ4/+rzVinSA5dnKyeYcF/RmUSj0dhQ
eKcVQM+si42VNOifwd+kDjFS1ECPUIlw/f6nWSylZAC4gLsBs4eoUlG1SBeIU+qN1bycq2apJApo
cflPBlFl60yb11mEZv68q6wvl7VLFkXW63+Hozy1SqhaMY2PC2ay62A95iJY4MRm3lj89oMCbE2y
UVt6FiU5G9tPqgyx8m5o8CRiI7WgOTfAhWALGq7tAPS32Bc3RpXEXMrMLQ/29CzhjWuC5ii/nZiC
Je8pcf55yCoLlvXisqxtKAMLtvF5ArPSrfNsHtyrzXuRVFkNiRgIvTagv1yPo0z+OGBu5l8jMGZH
HV9u6SQeZ9x7FZiz9xOPbqqDr/OXfvb4zy0YUrIUYX5/To3dNJ1hIQURfKQu0jLpU3xFzbZETBDS
o5JXAxOP5KQDSzw60B6rq1bJqDv3I84BIHvL3B87X94t71dLr/U941x1b8ZP20zVxizrSFx8YMry
TLJe4mHdgRz1ch680YAt/HC5lw7TkVBWUo3SI2qMqakoBuDwWVFCfXe7y5uIZKryKGPdQWiqIwUy
jOekV7k3T82nVyz+Si6VGi695D6ZF7RX8GyjJnsGiroxu9PB3RrQWBjimNUClseHMpT4TLenRKAO
4bNMhdpaXFC0eBjqKR0HPB8o5IY1BXnj3namOKxFVVpRZ36VyXM9Li/uwhGlSqgXSJZqSLunG56g
xxaKSxPL+1WeiC8oOJwuKNrmh4uP6B1QoMM0PmVDNyVDWGqYb4KBTgt9LiROYQ9z0UTJtzPglc/8
lSsiGkmGqL6GBbB0iXZpVqqk3kzyCj8aMWnJBPzkrG0zIHjtoMotaFtCmnmJkteip+OJoixzhRdk
mP1Q1o0VTH0GeZajHcVBmWhzcTBGJelwTdgXqNpzwnk6qNJiqRu0Az+mwDuknslsrwc/3mky3Xik
nFGoCMKVajyDRGfJktW0JBmewWak5cqArnq2zPYo41RCmZn+knh2oSmg8hXzaG/b0gLBZfSOHw1j
NV7SvG9Mzk+HKSc9mbZbILbprRWQl+tdWy3kMAXBB/+3syjUSfdoGerIH14D1fU8ClAr+G/FnT/N
AScQ56hXg/msWZDc8CUpj1559tFCcqL5zTwD+vOUMJhrqJ7Z8V2c8mSljO8VOIYo1IppzXetq7aG
YMZMtnfYVa4TkT76q5U/WXfbx8qeTlNJxVw4BagD7DCJlnZ6K45+cmm2WMIEFKkqwbCe+4/HrwnZ
zdbG9GRHsXJBR55hSAUWmQZz9KEnffpSxf/4EYwm1+9xBuk8U/MIwFiBfL6ul9/TAmXIhRSroL5X
oEYmmcCxrtzjMzSwv1J+zENf30PDw3T1hpONyudbJw6JXrhl1D5KMQ+1ixU0g+5bsv1rZ3AYxeEE
JABvnq/CMGIgTiP2eQBHb3geZ5Hq4mZ6tjn3XQD+hfSaaWws4CFGtzH4Enp9nQPCjLqNJajhk9ZK
Ayu1TQk8B06/somBrHutOrElJF5RqR4kO/MO0izi9bNzWeUBvz2HOcGT/K2Jqt/pVbjcXzsOGV74
mwexFArprUAdLFbz8PrKLqFBYtpwi4weX50/Kn7e4DHST+/CLbEOGJh6WZIAruug9tbEjCTn+vDe
giGkqDjWSL75y1Wj+y9phbnZ2FyJ/W/iE2LqJm6fi4G/tcGzSWj8lb0yxXxeI3aTwkar0zxAaPGU
XQZgRYGoa0LNQZ449w9uDr9dHRsAM1c/R7OgNFiosMq/lSkeoHBFTaV5SProIHva41jMHOREXj0l
SIo+gwFPgzBzHamQDqTQKWrJSociRZAzyB9408368dyEcr2pchFqSkIsFhnAH5YCctP01pV9FBdm
f5P77ehTgYAcJpDz21iQPVGS7o02z/Movz1wN9oCBuOOaj09iMKnY/GUryMOIX+5bOKD516yRddi
Pz5Tk2Bwh1FNqtSLUnA4D1/85E65Sk2O3s71iug/ZUmn6n5ZvgUrD2E78yx/KPvm51p9Gubf1nDA
4idmRvwxDLq62alIDdGYYNztq7DVfTmUHhXOryLXXJErZ25Ka/Hqk95jSmAPKlDK4d4DUyAcKaad
l3FCJLw9IeJ+h1vse5QhaN3AYL5WS2nq7wUvkkGAViupcZvkuaYLPgvbqcdhVSt+pBsEIU30lryM
4KL5lKdjNLBnPlaT6CDjycraeX9yj0mJBLcJpxtL0jULIvIWJrwHkjdWl8yQfMeTr6IIuRi1gt/j
BXAtSk+fVku3tgih/cmzyPlYLpiQ/GRVNz/GOZy6q+ymNqvJ4YyUQX1JoZcg7BYW2ro0gY+OXA8n
qsHXV+pcfS2HRMdCwbrX8mqEFky7Fb/kcjvhZG/e4HDIs3Ior7LF3QsvfsvIjF2qIRXeqHFrE+W6
LqABxrC/n+Qjb4xJ1csafbjzhBppL5eru0Ra8cHCNEePuD9b4HBkbhzTf2NoMEfn/nl7Rm7U7HIT
6+9n1kw6fwcAi1CqNudC1/z9QHawtCXICJHnOuoxH78EIhiIdkkCmuKiSeQOODCT884ZJKAmPxVQ
DpSTX0mmqBux5/60K8uw9J9jAJD3odhggueuiq/TdbdB0JrUj4bC2Tv9ZL70kSfO5sWjzBbFRzNf
xyXLyYWTvHlp1Z0puPFzQy1XsgzpDHlTJTPq5nVskeQKUCnJPmtepv7jHoCAerhG0aVUTqOTIZ9W
XOcvADrdoNp4De/tRRFnyr4oXKqSjVU7pW2jP6dQ0ICN5unRFin1QBMu+FwDYoLHrn+lnTm9dLyK
oV7Rx8LJIywrZD6tgdufwlKWIPe4SwwzLXgd8nmOWCJl88dCUlJFLBGr7a+KPGhaVjp0nrBQbXV7
be3WtOMjkMj0Lfr9YCtLX1tba4olXPaKUtNIPtKpYCIDCe07xuuzG4T3mB0mAzBu8d1IqoT4CwJa
TRAPUgXq/j71WHlKWtOAu1KMuLsAoMczCF5waMtE4c/64HpaK9p99y02EMrKFnVYUTdanyqibcIn
JozglHbn/S3JS37NT46gxgrZAYlGGuCoff6US0lfrtixVI3C+jHF6HBp/AU2u5Wa+Y/omnvTr3/r
sWX7M3OWCV1OA4hMLCCl+0tbGWkjlw+I3DDM0R54WbXjIn/CUokZMZdj3XfF4V4E+sOj1QXz98eA
w1o4dYimAMi16uGRKO41wG33zWVqWKSzu1UMPMjkJjSigOB8hnGP7OwclwdRgbHhsPGD8L10m/F9
qXUxujoBuvzvEAxe1fpooOlATRxmI2UuUmLXzTdn8bNxTZ8/12Hqpxo8haIu+haJCjwNsMMKE1tu
VFj/90WqLNRaCx86mcYbHd0hApikH9MNrf+0LdzjkXsT93gqDE+9fxkwe/QGfmZyjWGo6oU2iS4H
r201yrqCD7CXgQBNyuLlQGE5jgcDmNGDOwHLEVEDLmk6Ca8/ZxqtvJfGqxn2JUA7xQoBPaKwzvS+
7lxG2VT1mzED/gKSqZy6dUqD84aVFqIwEPE8PSaytSSq+sey0B3wR10CnLMVau/Fk2NgYTFMdpj0
S4d8kULZrmQGzc7s4/robu8pfVdSOVnLlWrLKIDJcZsdodwiz3jF3FBi97pH+rzQ2Ze4wm+xvIY1
R4PPNENLlEP6w+WhxmAGKH2xO2EW6vAd3pZF5cf99fsELWc3vPNqpRZixbqXPvfxReM4io7dcgHD
xOpNwqiifZSKY6hOyVlsbwnUqpeiPz/f1bMVDzm01zq/nadRIE9KO1zj0Yl5bqXYsz0nVW3jCjoj
L8BpB219SnnnSpPuNH3M6W8o0pMjm4N37X9ST49mMqt6nh/gF603/zGexG3oDXrIPoAknpLVymBw
tacMU5Mzw/N7eeIFP8sxZAbXU2Ccdq3fOWWYE0JrKr8U1pi7h7wUvXe5xrAhE5HVCm+EkpTCw0Yi
/DjipGDr+tao20CBPP3ietlqgNJi8Uon8kkwmX96t1IznhiTS9V7v1H3TbyCV8CCzMF0mIuSYT3p
Cdh1U5ZXZ4D+m0CNEsz4WtqRcmgCZwS0cbaDqjcLeaepTRoT3DFeVHeNxlc8etf3iA1j+B5mcXQd
bjZ8vOdfgxR+Zt/17LElCV1Rn+VMaTLv7mB6+tK0hjuQL7Kdldfd8N1C/QiTK5bOqAuKLTb6U940
/7qxdiBbaRkQIgEYKVSwLNDoImbPfdrcaVQ+aUlM4qinfxU/GA3/a4XtRB6pn6oLYN6WnxeLpfzU
ZW5fQuC/QKRCjW4M1P/E+GZeOVZ1AhE/KftG43eekOivlt9nlSTfB+VGrwQV8viPeizmFb3KhOe/
r/ZkUgg8xOYK4gsK+U7pAG/TdEMMQgEtzjV6QVmrMbn9TOHmIxia5XCpsrSojFxI0X2ZIOlVAy3u
OGtdZqcpLQphL5VOR1EAL8xbZyImUZQsgZV4gyj6nDxfaatod78ImLm+RzbzFFgb/RbbDqZi+z2x
AYPWrFWYINYmXRylxtgY9MunA5/JgKkk8zjU9i2sd+fWfIODH563BqT+Ntz4kYMhgikx+ESi74VO
O1tiSuUNPz2vz4CHkHke/GGNS+WMOgpKetgzjRf+yyrcN6fmBYQZTHbCsiYJG5KG6uc13vV3blDJ
18+YvdS4a71/IbAW79fQcWOqSnXmIIl+tUtfcqkUuKJh1aJkwNPeVMnTAaqmhfaDDjp9IRNJHF47
zqJ9YlbS6CBmGGPnkGUJnN3KWEW2FAdcIUylDnobkEO+LJQd91tHwA3J/0/Y5lNH7/2B5CkEL+v+
v0fY8HkTpySNDKi+j0YaMUB/7J37CNKRfO67lYoNYe42oyresP+7ZfFsZjwXAoJJMm04NLyExtdl
EfNe5tAedicw2rJ+6dNk0+3EcNkQHfr0ABo+h6nxqjQGVIFKN+7PbJektxfVFcsqwKUKAFJKmzzP
9HhU8twL9yNIfpOZW2EYDGvxRlUrktroZ+/DO+AMnNkGaBY3YWnuYe3RpiDXG+nIHzsnzKrj7w5z
peTzIpCsIBcP8kdmuJdc9osPvBZmf2IADl7Yh+YEA3wkbq89lEXic0lsx7OZvoNsR1M6NowW8h1+
KM/cMfhi2IRBjVw01/yl9z6w8MBLVGmMR1uKmu2Qc9p9Zi/Ot9FZYKrUpLYc++B/mm5w1IF5iD1H
39UxQoDLQDyvStYcsJbiAJfqPDpFK1oxSzEp3ddt14b5qy2HC/rk+CQ/7qmP7ZfIEqIFWxoPDaqz
8Lfp9E05AqG40GBqw/EEQVxzoAf6fAVlTFVnESioWzTpszzjJ2Y9ZwgRoLmp5MjKeMXp/AyzzzR9
GknHlDT4PG1/5M3B70WJSFsrUUXqMGlUF9JkIgDmsTwiY/Q2bGZ4VNWrGXbZ4p0ezKQeoIJmyzYR
juUAYQ5Bw5xUYYhKrBCBat8aJ4SXfkKy7UhocOFlJKH30/dc0uEDCAghAi7TdQyGkl9SuQSo85zT
GOVOW3C7ql4K84TjBtGcGUIjKJDuTr/8NESU91XErc5L4nGEekk9xMsF+Y9JN+RJ/73trqS8SNqp
VWH8zvWmfUHBdF8JgLpyfscSDQQ/kqO00TiiyGu8JdE0wcKR+BXuy5lRwVfEGdsqU8flinF1hCyv
ILKMZclE4FLJtXml/E9LVePSp04eR/fhk1n+TfYEFA+7y4wjZtno1D2xQX0th9b9/Wa7FdoEWpMN
6ZXY+ljL83oLKeulsP9KxUbIhll5IP31sicNXxlxdSJnoBVB1sUepsTBTsekclhnO2yoog43GCHb
eyx1bHpFDl/r3h4YTcQwITe6XEdPd4hzi5xlr9t1f5Z5DJlxrERd04r6r6US+WezNfRv+nQIaSF7
J/iGLnAvnvjDz02EoU3sZO+0ii0uRUnZvkujUcIH1pXvk2UwT6u3okw209Lj4XKwwauPQ7wIUL37
9/85ITj9J5Ie+qXHjWrvqm1lW3CIb5gVH6FmBYasX32ZHxJIhtr0aIFvRFSKG5KflAd2wv0HVysf
XD+413H9pB6xWR4rPgQbCwHc8D7lpJFi8JmfAiY9HLzNwSml4tiGI3AvbLXhPuUMnHqPew1fzTPK
tMwV74KBJ454l5fyCn3Svz0F8qEWPVZeeAencHQJE4VlZplTX6tZj5lfqhx31q3h5TxegY/XM33X
yPufqjJ33oJUqqlSzr7TS4T7n2sShmFrocX4x5fz4vwBLwnuN2LZPRBu05KSzbpaH7TaXuGQ33H3
N0dj7l3KUhdGfd5olT+YzDxJDyUVmaLiv+U64DO0plS6J9J2Fnib2XsHv/MJkVY5bkndkPE4c2Yq
7HILm6Lm0zJa7OPVLICHaOrc1tOe9Stnc0zu8kYQDUKCb6CtAs2tej+6VvoAN4WqZdhpnPjveYEj
+dXqXinLuStgHvNBKnoArDfV4n6SogPncdT7fXOkSdAGXO86W0RhjVoCMzvfoDG+P8twq8eMwpkB
e9rBxqvRxaGfNo4AXd5xqKJ1ROlg6AxsL1Pzw4uwk8iualbvlb/g7/rlJAHMbjkYKnci95B9nW5i
FrlFY+UShVuUQl6Xh9xH56qGcVaTcVURxHrPZsMudqvRv9U6vwIjDLKLH1JvqZJ0/EWxVDuH0Dny
H47Nw7wk0ohoUc0MFYWL5UtUCbcP/w437eWA5V7ZyF/JT1b6Q/ZmsNIsahBM+34C2iWXR/tchSee
Xd9glc7orXhyUuG/1rpM+Rr2gCkBa7o+y5hE4NkDEdaHsIY9edz8xvBxqfX/LD/K4mvACpFcoAnz
goQsN/my6mUlgE3FBx56jrON9QigKzDzASKhIq09Ki2faetiOk2QZzm11r/FHh1/bcdH7/UVUb2f
5Dtyd9/zidHxPHL8Kxiz5y6RtmegQCrvrsvZRQwdyg7maEiOLVctx4tbPgnP0+0gR+BV7B+6WQMG
Nz+v0Ta5cEDwX7k1G1XOAsPKdk8XYO8ASlQhHgXsz9dhiAjQPXXPN3mm4aY80yPI9m6F/erLwezq
KyFNHiH7YjzTW4g9vL4/GVU/3vZQBVCWCkEKl43dOWPcK9baTLn/a+6379Y8Baezuyrz7Wi/0UDY
Ikx6RD8TWAxYQxYOfGrSPAx3sBMk/6QcqvwEUJiHLJ/hLl6ZiFfGSBfsGy9B628t1FCgQwx0HAGc
CmALwIdZGQBTjwhrVWIZi/Rkt/tH/jfByPgYN9eHJ8jhMuxyDUyfsV8p6rezhDQD3h3/0uAZ+xbK
DOuuuj/PThtw93oHC1YkeoVaGdEJQHgGFIn3h/3b+Wsv1uceE5syXgF0jMcvsvUuGkA30kE006uM
UwHp1B0m2FKIBOdsV8gQ02NcAByZbSgRbT4eMyXPMPBKvwdMuTvsx2F/aK2qhZj6DddhoYev0is+
rJWlEKyY+mkYQcWs7MNmkEK0cwjoj114/AtDLnoZ0KqI8v0xQond+BsxBNRmZ17SWifUt3hDbnxh
p3fpMrJzhFKs2AIIjyXNlBpWBS0uVz+ikE/2y8hXUR9TUiMByiJrsDuX9+XzR1HkMiYdhQs1bQrY
JrdNYIcnIOkSEgmy3EafB9Mhk4PzQ2zFWagTd/+BXLpgGJOfXTP4K5/lNEFXgZOuE/WDQrI1UGOd
NWmJM6rgjcj5Ox40YNTUE5tjUxiKQTNQeTJfynXHCrPicIIUFRDZqbxh1MntvhLiglSBPe+43MHA
7Y0JvSAhfUbHsyfBciXRPq67CckR7R9WyxVGY5IKb27poqjHaf79Pve1ytl2P7l1Kt3dUqQAIpp4
O22Cync6YxW3f0DVUnphJZgsVAQqeDvR86sjGVP80rUjRZs4JjjUcfoLraHgTkXR0AyKRVSUsBLu
GqXLE5GOUPsWzfs8XEzyM6auPRICJ6F/3FD7xEAPk1P1FwTM5N6K2yKZm+oYGbCWcesPwf2zlLRY
JaEyUyq/0mbp2oCKe75UaCJpVMPrp7a86SAvxgY73UTLBSLMHAhZ4l0CR1YBEoxIpt4lHLECNFV9
9yqz5W5LgUd9rusb9x1zwSK/hSKAvRUPrFdMV8LppGVBk1Nrd467SIQVg/nT00Kk5e2Pba2hvm3D
Py+zPq+CVp9XgrXtZ17b3xevqj2II3NBq8ZI+xj/FRtoBeb0CdPUQcVaHir/JxSCpjkt6C/Bfa8C
mGWhFeWOYcXDv3MkuzoBB3Rp95tsFAPE6D8E2BWIBYNb7HnfjbytJPOdylI7C6Kwun/jmmPB0VYF
AWSMpb73ylwDRl62C2oloBFa0+7wkCa21/GwJxYKT6OSwooGzdIgXhLcNfy04qOmqbZdj0tDqnMf
bHHTUTpAIO/b2mjp8jks/QZmVyE2zfQtaGitCdr7RBwQeW0F6E2ChVGE1UcQ8pmxiPUxKmJlhNsK
SdKaiiE1G1f1+l6kebkSeqd9ijbCo2ORfbC/Q2g/TtRhq3IRIv0rbIRrIwK5wgrczdJSGsnCJCUh
bJJ5cygfmLvEXoD5PW/C/8KBVPW1PE24l2cje/50KRKHiDeeG54u+ZEmkpBDvX6vn1wmND7SuoQz
DkuO8lgM+4yAH3E+mhGn5JMSlIuRuDT8fdAM0RyYCBSY9Esvb1I9KDB0HVk4rbWeDMKFr+aPMvZj
AY9+YDd0v2daaoF8dnlXXWxU70yMO11Kvnz9oN/Px9ueWV7VGWF/cCxaVSoqj7h4eTYkYoNxxi7B
dQ6d+EukNKF8lavzvOsLsNqsGgqaJCFAyVv3yRobmXo3P3dHOfEfM5aZxkYjUt5lyK/S4aqfnpPX
/jxsU9guSWm75jmjYBGt63e29QOI7YqwfYUyUoYP5iZnJaroYXlh5jl43m3U8M74WQcSs6AzSuv0
/qWptWAFiz89TS3cljq7msn3JTdpAcfGwcQGINUT5EKyDQ/SVLuwItCO92CsoVzwKxm+pqgoW+qo
MMIX357R+m8BDZ5Ttu+Fyw0z1cJQNHVe5qzYjmq74nUjCwKQ2cs/xSnnLlnKa9qkgsfh7ODUweu9
zm6A50A/lbGXO7lMNS2MwZVIvEhxwr23g/OxeJZHas7rxEd9PjcdeEu83yAxZrT31xiDMUabRYW1
YSVDEZkXN7xEwLm0hlqUNVzHPazWGLPnHrFXxmXEB4TBHtGEXtxTtbx0trFvdiYVi5NeG0aH7CaR
TibfQwBML5mIRYuklNhltUzFsBNTPhTDhaXXDQjQJir/A91jznPLG/6O5VVu4j5E9iPHBSohmD+P
9jd1JCR3SHXQQtRLSFqJ2pEVxrTKBtyTKVF7YzL3NaXQH43ePoDmD8R0oLpu7JxcC+CAwJuWzGlK
7acQsfGIl+kiysxgQRouWPsNH0V1u9upPdYuTVKncdJURIqUCtO2Ym6QxPt5rU3qnhr1woHf/9BL
KYz7/dGe6bkketghuBFzXvwTaU0toPdFOx8SbYo0WlNkm1BcWt5hs5i6Dw0n+Xg5XW3YXAB8e9k/
Rr308cWkyosiCKdqwNzM+KXyTa1i7Z3chtrRCsluCZv0w/rCpDofqPlngqlfvlWHdmflIf9LZnBA
tJBExl6rXRONd8A5wTSiliXn+5AqOkmvB8tHktn29EyRuSvWsaEjSFdNo5PiPtjcXg79iqGUgkl5
JANPq60kTc9vrDwEYP+nzWtZg9P2TL0bkHO/WrSJrX56frd9gbflrd6Iz97zN7F2Hz/Ei5Nw8zVQ
P3aopGBVbnGieyKWvteHuoabj53KhMONg0KaF4V9aU77sZZJIjT+NTEZe4ifTag9+zhVoIoteV1y
SqOBvbeKGcaYoQY5sRnMFgCo55v/Z3IJ9Yo5cQ7PX0KrO1bkyYUs+yp87HjGFSdkuXD7ji7+GIQ6
idYibRRL+qX97GGyEIwChYHDqc8/96Gr0wARcBzoHOgXKHuj43tfm7fg0k+aS5lrpCmfFjVx+mz7
1tRDHx0dWOwxKzX/HhPgXzNhcMooXVKLzg+WgMf7tUQ0Ni2/j0CeJMx4tEo/faVmCNq2Kx1JEmpx
Z0e58rD4DX3W73XtcEezYgUNcZjy/ThImHXNIxahk8WA3ntr4SLnyntRV12mwAxqXRynj6EFcaVx
lgvhqRT9hrgl+c3UkDGAO8o9lg7NL5SkVtsXDgW3qZLzYAbdxU6s89Ff7pzEIxPYMlNPnpJ5AW5K
Y5qyDCq3DLCUv17hlRVJZ80mTuZNDpb4vGENXlettBnP7SOJOlPSqQZYUy9wbflklKzjy7NDYLBh
tZnI90dcB+esu/zqXivIok/YsGJ19xJ0r4v9JzIhf2ghZlL1YHOuhyMa3+uZd3gta61HEGptd6Mz
CHp9D6PpFl6WbaxIpY7L8ZarPlq2/TU8bjb0LyQGpfxanRoAPa8wHV5N6XO60B0qUpL9iWTZuI54
r6+Kld44J6YcXVLe4tKhVyJiVAW3gFNUJBIM3EJ+svtl2SxdCr2Wzc2vkd69RRwJ31hFsvHJN/UT
dTLPyG8RJ0sa9riivT+ga0eisUttLUWdoa42Q6yypv2p4SNf5VSppsQpK0pHUu+pEX9MBlX4MEGR
TAW11rO+Rq+9r6anWExSxJvgNMVcfHsUmcKNujUTxMf2TJlTYH5gJq+d1st7DyDugAUWDfjBL3Dw
T/jFOqUVR6YxQ/VcuhTEGCSV1RRD8FBUPQQZ0mGWM4VQTJCHK3o6oZAOwbudP38bKOs7Lw2gNkgc
seyv2jpjSfNSfNEkj+HFUshob22v4BoXCIA0kdzHT6duOO+VMcevGQ6WmNjcg4jYJumyTqWXG2Al
WK/8UrpgWPUAhQUjvbE6v8rCjGbyCSgR21B6UcEF9zfIHZor344rJeVhl0cdwZkrNOFesoHfzVUD
HSNaEUJyvc/rTX8tSyPYENGFugCgrqSYwBqyggxMX3nuR+2+txPJ8ck095bNRD+0wyT6dchlps9v
BLXwx+sS1sl0WrLmF0Jl6wX3gGDh4GIZUTqDX4YdXoinSsBRo6ipp+LMGIPRludDZfTaA3+b7SjD
0Jm50QqcrHMOrQPX2ZeYx8tqrefPilWc9e7R4ngWJBqINpXZnG7kwTCELPhu1hkRg5qW0Qcc37wK
rczSErKz56keREjF/3IIwOfXkWlYowFMiQethVXi/04xS0kpJJ7r+NmXYOVvpLG8kPUpvesZqdJM
Nr8XrtiW9OfbaA9AP1Gtm/Fx/5W5GaLffq1jF04eczE+IBr4SF2WyHLAxJdUSHSrJfVPZwdZxVZQ
TwW+mXo3nCRYL1mcNV45rWmtq7ks3Rpr4AkzsEvT1KV88bV0Kpvqg8z6OBwkWFYQsdlpm8xCkQ91
WEiVYcP5DcVo8OP3IrumBU7Nsn4Ftb8SWkVXugI9L6rrynWoUgUk9qoJaZTVPjX2LAK35dW0bqvL
GRD5MRkQRv+lih+ZWUhqFQjW/KKcClvjziZGBkCFCQM0Twbmi5lb/SsaeyzrP8aKPxDG6rPeUEO1
8bJKeU//Tk4AuylZTAsltkPri7EMr1LpDizMvY1hyaxcKmGEXCGB6JePzOjFr1cA6BLDZGoNsjbD
uxZS/Demzt9FOJJW7A5GPTpV0MEu9Zvbv+axo647GEFfwSeZRt0Bg56Q0zWuO7IIY7PD4KuQ+TIU
5Mtcc4FHlZICpViVDkJTn7MX/PdCL5ui6JEn3rOJMf7dD6msziaIJIK59WErTPrg8CFiNDnwx+sT
GGR9ztpAaL9KBlOoP1jMS+2ponreqAoZfaX0N1g3ebFSutfy9CaCdpINK47gREo7qWQ6f2f7ZaJp
zKstcVN2DSszVB/u/jZDQmTIt3Z9uAYdAGp9L+2H5WSLov5I5pNYLVN+fv0UT7a+kN7Q5GGPnl++
cO+81TqksDO9zqlnBCw9E4DjNdmsx8yAyq6c0NlkQ0AvNc5B1PEpRwLTjvXOk9hsZzoJilSweZ1b
15aNmaxv2nMBVh5n+f1WiphxNV4i2dDoMA1LR/GyajBdku55G8dOuxRU3TuzOQ22mVIXQILoNDK8
HBHWbLajfkjvRQdqWDF/eG0YLiNMjDut7UwZH2F4sljeDlNMHgHfePo3b9fjZ9XlbSdXHwi8zBuB
fQ5GY0oNAepGZHHtKcnPsAbxozzETEt9QsicocF42ctve50feOj0sViUkrKdof8jTcnomBk58LAP
Mu4V7SSy9833ZdsFdy5OevIYtr3THP88HR+/PIedwcqFRpE7BVixmmwagPn9fhd2xU0NQZgNSEER
ETxNNXI27NK49wVCxz5fVS6WjSXdNnj9XJA0Ln/XxkUPaCOVaVVVH12TyloWr+l/eMSQ2sjZ0pQj
qrzplwqKMIMVff317p/q7K1/Ic6DbyNqoIU5Q5XUWnq/19Pp6tYi25sFL8/WhQGKOuDDdTiaVjlt
PeY3h3uc5i0+HLX3IgDOEChFMCWsxDiJuNYMlArIwGx/kLha57NJ7Dn+nsBFpUBcfWwKw/wvS3Br
atk5//ItNnTwZEVDVyDH27KiOn4Z4zsNsQXJpg1EBrlkAwcSwTLHVIsTm+QZCH57YI/xYkoXEBgm
dpwF+wn9pEqdWPfKrKj6j9aUBoClB/aqTgykH7Qyn2upqaDHLkJZ49ybSkRv8YP16tNOkM8cjNCX
J6YqmD8BNoXQSYOXzVAx7hluwLR65e3RFfXj15HoKg9kuzNqEfpBj2a+LRBYELu4hXR+LO2N+mQv
HjzIJe7HADLkaAaZ4KXgRuNgV23abc3TlSn+ao70tagrjy+XrJPFBPpUVftL+EkCaKnmPrnsQyu/
GOyFBX8ARHOPJo84xwg655jdPhrwXYcFnBM1MsgTs/ml34xQoALwowRVkS4YcXxZ+eQSeZg66/yF
28eQgNq9MCOMDKSVBUmP1gUESNrjngol2ITWY36UOlXpfgnfIA4At9LuedOx9oemZgOCI+eFMdnc
guMX9XiMS6mEX9Hxrojm1Z12SX2hgzvjYvfHDnaHCTXfeoFNcrT5CdoIZPaOQra5zgzgFAz1SbVh
p4Lm6yabAQVZ11YNWpYrOEIxfV/16ujA2D18bDjqL1+heLUEHnj/Ck20KhIM7mHw0S5n1Z0E+wew
eaTJx1VXnpj52YOjyCEILeqX9foruiOEPYeAthk9DKjWtRy/nbYTEhjNdcvAaq2hlDiusULYdDT5
LYhpaNKqlrSaq7SIIO5R5wOmcHIS8TVXhMUs7Z5DS34eqdflhu0gM4/yrTMR6o16kdiJLX7J+BxY
M3YYM8ltyIZV3wzLg4Iq+SPMGgXKMshUXb+YWirQDgfl+n3PxEjb/NviCv3Cx4BNf2RSwn/+qA2u
BmddpDm0ZPoKs4CeTPymfnyD5s3MZ0m3yLxQvZjdygFDirsWztVFj6lDid/1dYsPRYsFRcJBld+1
XIt+AExKsQwcZx+lHR5W5pvEyKg0nAfHKIZbbtPZFbfuxFoq5x3QjQUUxXjA5tb8K3/npKE0cmNb
yjTGqYydN3X4nPt0NvzKmWJTmOdrO0f6xion2uWos1VRJg7S5wBT4c+VbZS9GXx021Sb6nBNY3gl
+97JvSvLn/L4s+T4cziA8g201Tz3DslHQoJb+pLzvrkKrke2potNsW54q9dO8piegNYmnuwGg08P
zL23BBiE+S9mfixKfbZe2wj63f4oNTP/RHcZTD4Ip1yd8FRWfdKYA2neaoAuX77smB114moLDJzX
1UaVn+nFQpLOzRbeROL4cBz5DPdCikGxdYcONQdXJJ2alMIPM6/sbgCW4vDlUYNDOUa1gVLhZiRW
ASW/KzA29cD9e8VI6NTJ9uFvS3XdkRiVEp2jRtY9nE5Da3o6XodWOvD4UERPa4U6jhtImQ3/C+6V
DNAkotNwPri2GuD1YSekgBnndHZZtKvJMJCX68z6Eb8YK/1lvTGGXj75s+PkD4sSNeTVMd7ZTPrT
chlUbdunu9Yj2tdybOQ2rBYtnGgwNxcKSGWitIRv0X3vf+P42OC/m+kVGyKwuOMAhVO6H424LOqw
f0HBfs+In4OnUeJBjCZtwCmPJY2PesHRhF6+vvnuJxyPPR5+8U8LM6A85X/BAnwPaoukhGuug0aI
ySwXY3ZqF6DC+RuPIuDASRJYVcStP+cekHwowg/GF4hlqmAyBd6EgMex2cBoWiCDV9q7XQoMt76V
5L3ePdCkoEidTP4AP/D0uMCwXh1iJQVhwBp7+W9TGIMxwBPUO31KqYx8r9FMrwzRYKHVcHtDYVj1
2cvIgZ/7J3qfMdi5jFCPGlvHNE5seWXbo8as5qh0Gzda3U72IJwD6oHSOC9ay1nE/SOnVOhgMlKN
mCV2i7uFFP6JUZnvoVVI+KSxgbc1EyCA/l37b0D0Iw1gaSibo6ELc8h0k3/2ys8pjB5VKHSj7wA/
p23uThcLxtoZ7wri4wBwB/4kQtmlAxXA3FzPuKuNIQZTR5Kj1zxTTnDslTKd9PvPeTQen+xretja
5xazGGX+TNc86ydGXd6ZZ8YI6Jyf9fauS7OcOQqPf4ZSAW6acFieMq4OnVxy7bJ3VAmbKCaA6dUR
bfAO67PWZAAGEffLaUMKKPW7dk05uuWPdL/uVQd5VOwCG+m03L4H7RUR3C/f7Vov7zjQE6ZdVgtb
enOVAecQUgebytg0MasI0l8lZp1WWlmRPkdibREZ/36YWuNpTXhQwQIVk6potK+Jn2ez+1SWTTMC
ZlAlDjeX4gV4WmvS9zoOsFSeUEj0IqkDP31RDtFmEcwX6sXMD1bS3BUuwplCEJhZBrd0LOwli2TN
0o051XIfYkjuYTxeXhDKpxtjGbAy4gfetRDZPOJX7eFYC89WRLdSpXlZxcz9ypSpzMiAlVHC9DNr
dnrd8nhkh12i5TL1iAddWM4ahFb6i79VoSg2FAC+sFuhAeFXle2Q3JR/oZwyvlbk6b3ju4wxI6nA
nyJ45NWUbwbvFcRnr59riKI/ZfM1JxDhDKnexg2MXim822NokRT8JE1vE7Ujz940DuRi2a84zYz0
9E7M8oICYwqaxri61g1OzEN3muNhijN4Z9/AJuES8895MgfZdsna8E1jCZo2dI8dBBd5oDftVZk7
+VzwlH3JyydCR77piiL/zqWIUPZ3a0TufKbKbau+ZT5WVj5Kq/1o1hKjiMiDpVPidij54FkbPSt2
O8yry5EbHDf+7XvNFx9N0UqUuZbyIJRjcQdOgbAsew7Xj41c/8PJqzT1uZC74qDHp/Bl2zQOqr1v
gQ/kQMhdp0udYwkibyYWLOJW3EyEr4/InDU9xyhUOI7NZw4GmQiv0h1Di2dNs7vHYK2HF4bbzpFP
yGXIU6ZFHiT6t1bBq/wz1dxNqdqTd956CL8kc2cnskmTwROJLD4r4eTsolOLT/r6l6HVGQ6w9L5g
Sz7tNuS8lx50s37tYvFXkty+XjOZQA9hcVSTG45aZrNgWoFnCKcEppek7XT/UwviA2zC2nWllnOH
6wjrpV9cUPQSxa6I1CXJtolzNoELnjUXX89xmNNb3Y6am+2hxrsZA/KQVwZ+cBZCGHwRgk4XO20r
i7KpXDgRxbg0+KD+aR0eLft4BxqET7/Zwh9T2WRojjfSWjJf8ac2vLu8PI87GR8c0QYsfGF7Gsw1
npqQLM8AMKKi5gvSWB/jTEVPrZnRJGv2oKQmkWU/XTzjzpfvqe9RWkh6PUv+cDe1yegP47tf1ZuL
61q1njLvore2xc212K7W0ZVDPjIh7/yikjm2vcDAh6a3kDYLiRn8oEzgyWSE8EbS2QR/whI4a232
jsWQHiehw/va3t5fYAEGzvW8pvZ1u5KNjGr3K5c4FqeISHOjz4nMl7lw+EBcVn6jDcLj1RZO2t5r
mpnJiX6uVBPlRyAouyFQGNqsyGtDEt/4wpRysqknNH4+hnWHgNlRzG8KpXVOPXfhEYv350dGYZ7p
r6eN+l+hoJDWnwnFCWl5Ee/1R5EHyv/WhTr3Etk97GCXT84+S660ri8pZk294VqBjBGz1ek8o85R
QpFggUNqy0CMKw+bpb0i9u/VRfjCPV0EmSYwNk2TVU/hAaMp2RmZYWathxZRav3J1Lt3G6moPhqm
9xSWPMBxNNOXyTF78uBqT8cDIiWFu+R9xjK71T3JZ3je/d1Agy+swrEJ0fNu7i+ApNjIQySgZ1B6
IZCHUwGTsLMqfvEPRJwTs5pDc7duneh3/ikE1dCAW6Qv7fOyeQZ0emBBY8zOIMbSvG9y9x17OfHs
2wIzebQDwpRwDNtiKjE0y13hOhTO27y8VXkC3cJHoQ4J6zZ9XORqVxYGK/fI/336Y/0HvoTprMzX
RotAfeYlDbwl1ZQbdegsSQqMHeDieFXSqGEQf5bU6mbx6zSw1x7BtmgT3X6vUDe7VjtESZik49DQ
9O3PPu+7v95QWuqtrvb/B09pzl9GYjvYiItTTe0B6G5esvkYrRK5pYAUeK/dK8GQwxszXPMdjdL/
kbLMrmpd46qXWDnBfPi0Bvps2Vyx3ZOs/178C5sslVWuBMAlP0hk+4DqlhOdub6j1/Ax1qaDFoXi
0l4s03G5lnm8Cu+YjD6PvB9kC7iX1TwPaOgSXymIAlpJTX2w/LDJvMuCJbCNTm1g334LecRhiBoa
v0+CQFeCCCRnMFMl6pBOY7mHt2DWDCTHT96Qs93rKCnv1i0qRtMLDnKN1+vdCY8u0tzUJZcGCYp4
X8d+KPwSp2YKi3Sjp3GFT5KKraZ/YKB00Z0vaLYrmYksZHRzCsZc6LliCeStA6Aeg7dzcwhDWl8g
PisRAaHgsiLhwpjwpX2h3twQ0lAETh9rMUhgPeYQ1kHJIiWgaPKR+Ad1+O7OQMShX7QFK34/SmYQ
S25XCQXRTmJ3ldbXs79ZETsVIq8GKQkOhXItIx8dSUKOexOmKzz3v7M1kO3azuwA1X1AMWd8LNLK
3O/ZX/JduMbVxiIIA57rlnhdrXT9VPMX6wQrNF4/Z//XauMbUkFrQpI0VRZ4xGHY/Qa8Lups5C+0
at1KZNF4PHkWGHIA+ZX+FikwcLOHOhqBmWLHnZ2d/BhVSAPvajYRdmZTTifzp71loiifAuiEHV7C
2OAxyx/ZcAq/Nk2DdcKk6EL3iMed7Ft3UcNzI//BO7gocvJAZejUYk4O0ubm+e113P439w3q/evT
N4kRhMZ1AbGncmMk+qd5VmqreTpPIaNhfUi2j2wMQFPHHRPYJnAwi2YS8HL6d3GOamJ8Z9AaIY9Z
sGPOsvqCif+wNgU4nL+RoSkt7D8IEladjNPsa3auFJKVkq1mGid2iEWbAyEYd5cWY7X43TRhn3dF
tXYiaUppR4RGLFkgBkHmxNsmB/WxQuiAmfwn0hotcWtcyazMJHJTVBquMo2XyKqFIrRzTmEOEgwA
31r2R4LzCzPI3GWG7MEHmpQwIJ8MJ9ERLsLHQu5XxZ9VmZ5T7JRLdKe/v7s+huFk/9uhNSczddDY
Eyndr1D1UDB8rbnZiWAAP/yE+f0p2IUXAzqHqcC9979UL1z6qerXgelt2m7DCmR9ilfKJ/71xQU3
azAquf67J5KR8Ku9dvX/F+8Mp31ftIvrpf5lDBlePy9LM5wuAQd/GK97UKo8L7+y1fNsHMZSZoSg
sJ6heSEG5aOJJuwNYRXf2sE+dwDNhOHChZZSdc8iXWDW3MIaN4Xrfgx2pZDV3gS9W1YkKo3tBLJq
uaVARwsVpK5zu/fBmNBn9D6OPvkmyh89Yy+qoGSsH9vaorgLlPbe+2uL7oyqxE3HpAxdqrruCheD
Acq0c+f2a3eKC5Iv6N3Q9JmROtmwwZHSLiTREEknpZFbw5ztLg71hchfDnVrjHlfGZQqYTxkIiTS
QBL2ZFGdQsvBvBWo1CUwzq2nc/OdHMk4fK9oDLX2I+vvLt6OsubvQG1jPEcfQDOhCaP8LnFRN1UM
XuJTC220uhmkU71L3KYIn/Ypo3wb/C+8Un2vPBJI5x6FktcACvK55z6HqhS5Gf5LJNW2NN5tCy82
VpjtYez7KX0QZ7epF+Un6KErPPdiE88A9pSV4YZmA1aO3ELFrkWmOvbWX9auSvgzFHV4maS/Ayvv
2s4/3Z/28atk7oFN0YzHcUt5YlrUfyqN9zjvH2Rd2sEvA18QIy7NCn9UK7aM2FFckl/K1xIthiKm
Esj3infv2k94sBEGvfaZg23VhhtpjuVPPqj6AelPo7wLBMAoTA0j3QPZIV6P7wCQKKdl63oBWMUI
w5KkA9YOUEu2j103yXqTcCBHtqX0RdpI4hSuePKdtXh88kibTUJJv97m7PEqeLo4s0LdvgnmNBou
6Gnt7+kejmb7lOAHWliE4v7PSeGt5C45Xj/3fU9iLZPwLt6mxY8rQF33FDcVIXa98OQ6xuusPI3s
sflWU/6Tu7BTL8hWDO3RkoBLh+9rDzu9w8A81Xp1pIW9joN2LT3UjpVJ+TcXXutcslWXHiivs14W
DGra37yVY3u4sr2AErgfeuf8p0tRaaEc76/ffEXfGs9oa0EFPaMfYcM8PMrYKDGrJ3xCu9ru6XuT
8br96vB2Q+eH82vEOK1b/cdmUmJLEDI5uwqftDUOcVKcp6NgUzkx1RgAUS3OZPJyDfchPawZpACd
QaPLLep94/YM77m+msWspHPn4/lXpmjjKc9xFVe0qTv8LV91V+E4WwBKjeERBVoo/xnT6oLxM2UX
zrhrJ6QdF2KPZ5rOY9kC3mo6YpYFE1Fmxw7VfMkWtFNRy4yJr6QHsGBqCM9TPsyNj6pnXWjNlR1V
vEEwSlsqBAD1Oo8AHc2Mx4ltXUrpo3ZmYqJHStXmnokK1+2xZIc0aWImOVZJ//QV65s3Ur+6Ib8z
gDGTQdy45AF3NRyGpe754AUgCAKrtsbRLPVEqSDLxGiQe2RJWn+YvCgcumK5M7gPVDzIh/JhpOtF
YKnkLDFOZuDLvO/i4N7OiR19ITmYwIZXurDgdSkUgjRMH914VKjFvl9Q+jhnl7qsLYo7P9JCJSZI
LPouKQvEVn8UQ7/65CqDDl0n9z6Dm2dlA483D/HDosEedbNW/d37cob1AYPn2LOTwXkb08/MTHee
tuBlAvGAV85IdabAw+IEXguWszoqO3v1F4Vkey4Hnx+tqUxZQ18dGQgbnQE0ImrAd60A7tVhzuQR
EPraabd7O5mLVyFedCij/7H3zp/8B+6rTSyA8IRULNl9yT7baZGMJgvIDpxm5E0NxTyfLDHiJEWG
LdMy3mOrO0vMAR5369iBItMouIEZ5YNDSe6Uq14O9lBwSDXah7Qtfsa6yAixY2Nez7qg3I43soVr
1VZ08JRxeP9+TkwqZNEVspEhRHHvAATIsu5fyy+OSQB+aVzTZ+tsYoYDF9SWtc4bdSeoH4ESoeF/
3ovreUXdEMpESJdkWnfZ5h4lxOdXsck7UIFy/UXxkyOiSzAiapuqySYPcCD1w0HeJ2G0AmVgNNEj
pv1aehPD9ply81oKviOZsIZjRSzD8Zof1ZdpQtAH8zzLBGl/EorMsyuX17qzSuwhtAWUKEbmtji0
ZJIfis7cWPxNYrQTznjLrAokQfJnMhsOT6JP+9xfdznl1dGuOBjMQCzAg1OtMAsMJ+CsY01+N2qu
w5H9AWJ2+WvSQbgxZaFlE3AsUM93G/P3bOduKWEQCxzw4Giq+xk8ORsojhpES/nCRM/FC6PaXL5H
+YtFKF22WXyEFu4NNmnbGXd/eu0xJIuD6i7Z8Aav+VtX/lq0tr7/dOt+Q67Dl9g30qwq4fY5F/lL
KQr0TJgbxvVMetbeksiV8TVUJt+SnaLyjZ8eyTznSx/2dowjmscrjx1L/7rVNAo51C5otIU++LqK
99/uRa/B6gHYL83+1VJQs7HukIk9IyJ0mVe5ZsESNCFpQ9HGrmGC4GgmqUlF6flFQS9kl/RNzrel
FIjrFFlWea+hE8sIxT88i3dhlVhbnPvtNA4YDa8NitTdetLv4R1i0RlsrlV13U8ugQ6A7oT2/4Q3
rlBHe7xH2TvHprgGvsGsGd7uv9zL3en6IClAYVH+/wH53ljkNH4J7eFAxfDYM6F8JgFQ8dyfKJNZ
42mr1Z+4pUjftF0hsSsDgb19zrjqSJrA6lTKFdY+7/PDsgYkXTRpM99g4dLcrk3g6sImM+ghwjXO
dDDN1lIQQiA7glEmnFtzMKdqJfx7uTvs2Jd9Eh5U5Hk3BWM4gP81rY5sOYMeC/4cJTRyrqMKNTam
JLiaIArk5alSZFILqE62hzsi+sIVhPeF+79GavqypwlAUPTdz/TXWrluZocFs/v/dsHN3JOnAEIq
mswkQYt+01nFNB7CHozVkLoedw2uAkbuGDe3WyfYDGM10GhuQKhdfxAKohT8Kv4k2efqPpYHtEep
m7UCgtJ02fMQxzvyU+mtyR0wxqKxQgbTXdiHnvkw6GHC6a4bH/z91z9zPqBunfWgW1OOwM7ekHoh
bzUapTvIpVfeP6xFSspxu1ceQTROJgqM9JMS7NFbbgpTfp9z3RvtUVuWKHVtLvhCYU53HqIjussd
08d2lqbK6q14q51jkIudXqFysCado8Jk3nqvO0Y0UPR7tb4DzMDxeJGbumOS0mS82Cb7dfB5oJZh
Q1oKfYmTTY9SY40KdkFeJJ97Esn37vsL9xJVf2RtTw5eiAyu05UM2f8oyD++LpxMbsgmdI5zpqrt
ER0raGCdx6NdYbYufWmomxSfym+s4IU936ecTfKhwhLLrX/PyGXKGRb5ZKdfKCDKDV1Dx+c3D9OV
GKMK6/48R91TAOw+NCett8hnZM/cVw8HYF7MvlCswWTSSdpM0EU/5nsh3gXHJ5QrytUdHAGA5bHj
RhqymErYQGDg7XyNabOPUHbORQ5kK0QW4hgM1mxwvo14MlAmGbl11A0vgnyd1Xu2m3mJPcSU3uRo
t3MPLJbnMleCGtJwar7qDU73Q58bRHn0WA0lTrC5omdU6dQiA2HkmJu1uAPNtt4ctRGX/z3p5GWJ
WPIq6Nlo5dcHbSXUZrrt5GROcxfSRPnWaAG5gfDq95d9GSpWbHYg/mhXL5wBXlcFOJCOyIbq58gH
VSxjzauE2htwF7xErGB2t3PFgWP5xtdvJoU+RVb/HBVcs5ww4feGvyUreAzdY9vvVPuVZKI8oJ+S
oH2jYm00q4lAaFI0LkDqYTuUIpy2B9Et27S1VznLDUV4aMF26xkRC0JUyaHQ1QFS4aOEGKqVu2jT
qNIXtCp/LtKYCm69tT/wUQ31nFE4sQMVWkuZ8pXEtX6xKs1ajsl+FVVvrCOTKflw6gJJ9ZWGO5oc
KtOzE3Sq6ni/3kHCH1JfWQRtprisWwld8hNjLLmbnIig+1NsN47coI7bY9nnR57G2hoAUdpa81OB
EfI/KkeZF24zlffjO6YcoOFXGKT7L5ST426PoceDr0b54nU0MG4xYKHyKpIVzDARdXVD7ViTFjPl
4zyo/L3Z0aFPpDZKrc0VpOqDBKKeT+LRi0SbtIB5IjKFm7xUwzuQuvQYqThuGK0eYiX36lgpX+bT
Z6fLR1k5LR7ujUMJPvnwrMYD8ZpronbCZp9gyeGHijpzjAy8ihMCOy3FtK6sHHoWgU+C04wa5hKc
opAHxtKl4lDWfXqWVZm14Hq1l4jtZRvRB1K5kAuIdxNwDGcQ/QOiCrzzyNc568iVvn8HyAt1/hat
xp0pkbFCcYDAMvELHg7c7N33pG28QLDjls6V/d5RriU0mGA3jYWCOKixMj4xmoDBiWDRTP0pSMe0
lzQZtyhgYecXR3YC5eVjY3nEKD6l99lD7LzUIkhgoR2kqXF7NCuAxI5EyZbMm6B6rZPbOL1364ru
qWs2UrpPPrx7JepcONP+8ixz3iVEYWvsk2lcvanaTkpE22qNMuBu63k5/+PEjxtcxB8V0G8f0hWr
n+QouYzCePha6lilRFAJA9kHEIU0hDL4sszd0eflxoI53aH/EJ56xsHy2YTwRRycfZBxT595aZhK
e6jtMwnMkGQxiH6unkcj5uk4fW30aj7ey72ObrVqXr+GKGF38cCFB8v33Uh/ezjFXX4Qmb5N7SjH
KR1UpS29/kGUyTzL93ORSfTWmmSTPv6UZpM+iJ37ZiuaDdNN/mV00UrSISZzhm+7oi7rFPWxZzox
Qc7GV8qHKiJ+2Cr6FqbVKaCVtLBVfBVxjnH3iq6At7dsUiZ05ChA0i1n+Yy0vtpD1FoDgzeW6DYj
xxqCxYC9qdIEGvsARyULRjK722a3dTmPFStHJ/bQ5tFXlhgd7CJ743SZLn4xy1+VdX5/nCkPc0Vj
P2yAhLWfvWY75xf7fxyHzVNIV4EwDOowxgL45K2p3pbSVBefmGxTjaxg8ZHxPxTTc4Gxxl6hSVyd
qjEwU1g5XyDV1k6huWxsuKz9d8DayTZPpn6VLjZxHN9b3BenCrN/zuA9MJYLEoYv0+4tMuh6kX7Z
slGfyBze0GMAjotmB6iHrKu/IHePXTgYu8LQSNTIB030WTMAhGOpUcGw//+rVeJokeeDZIO3quLU
a76FLD223dR6ZsqIHX2brwWQIIHpkJS5A9FbFxv4+jRb7oWiwXAvNwWnvWIlBRDikQ0z7G+3mNxy
ehQ6/ghu1zS1Az2SZoNsTgRzwCAidokYDJA8pLOE61eAIb950tRZ3Bgk0g9/VIhLk2p/AjiS/4/i
iS+QJDrILcgERzd0tkuu/IA4L4wmCwYklw/DcCLZmAdXuooUuwcn8jWR0kV+7cVQIguKNYa4vIh0
zhliPyO1S/vxuZGta3NxVPqllVqaecV9QXETlMl0UAvTuE+xKg2XDmBP9lWlCH3upP2buR3c0XT+
GljwBorj1O+Q1UlMmuY3snhtyVSnvZTYdv0UmsEpnVIN+Rt7rPkuZeclsi3AK9qKFaEtnNgn8V2y
I2s1qs4vQghyJ5LwDaOmIF+Vkla5WRtXRmG3alQ45imNV6xV5ZBXZCkbVI22TGyBetp6tAaFJ3n/
rNvstC5i6pLAwVoX8s1n3OZokk2u4A/XRL80I7GM+86OhickD4cVIqakiOfEMPGZaEZUMhiPfdDm
1o7yvDfnt7kOr9/Bw2PXHeAsKqY468jVpmlBbZBtfqNbrTkUcDKyEhgHb1LJYhemGU0KqOaWRoVO
P1wwBy745f+9fsGF1jjbnzjxeKQX22BSrbnkHdstNTU53byWFmWHocpybbdtmhqbk6s9oa+GY2q1
ieGKkiG2cEzfRWdGlHhKzefF1J67WAMQedQnC630fiqtxBIveaQyHw7jlLFYtRU/5R5lzZ9T8OC/
uZOAc21QNA6aKb8pxu1q0iwMFCyh+aSSY+JF3zhktsbP0BC/UKRhS/utTJB6A9bcE+Zxdy9dzLEE
2gzw/DuqCduWkS7HBSfrzYH53005oV3zDATbpoioLoT53rTD9bLfxC8bQhrtVOW5o63nxoKY5EDY
iPymsG3T7r+62yHyvSipfljYT8+bv2Q1Xul3V3ITp/O62AdJxRg1Z/+3uTYsCQX40NcQy0E/R1IV
u7MT7phfyJiNboznK7VOCZrCzgn0Uduz0AkwO4rFie1JnM+j0vanwYdmRxQQBTOv/itO5e1fBbCn
4xOWaNxSiqQ0WRkUAzwf0Dw2lY47dnlk5SXWZmQKX44Vyl17eCKEsf1v6jzd7BFpgGGYMa3V3AM7
lJyVLqYEVlFX/FsTkIOIhKp4aoryyimLh8rrpI9uJMKHjRtdIQ4Lyw7ftbVDzmJPBKi6vL1GBtyF
Quo7akK6bofVCf5CxIPm2J13hDKkhUz+2AI1lgLLNCMGm9UBEZIRihLA56pWSQYsF7zVB63kgypp
jQVmDrZ1Y7i5jqQxKRZ3dKUcAt5Zypqt7fUn8lCp1qrIS81NzYw9CpgPn4Hbdojrw1LV91PT6fxj
s8arNOl7/GbcbCUtKocKpvJeBShu9i0CLGH9WZaXokunLYF66L1ryX4hqMkXfJyf7aLxvqzPgFkP
+jMJr/C8nqM6HFGroCk8HuCkWvG0vbrDPvmYa6nDRnUdC6WXtUDjIbsDXOKRBuZ3JMXubJcl8w4E
cZmypAD1LxZjWG9vqgW8tqiGmEcHmdL6UV6wYBk9/hXS+dUGbu87KecEtFJ7UlGFvv+EXUSgmSps
UuOFSlt5nN3Z8Cynb5tiXPtsIDbmOEBbNnYkFETgoGijpEyI15hsYDYPOH9STK0XL0Z1GTrG2ztu
Lms621VXHo35dbnmHaSk9FdaKZmDdL3OocTnIw7neJLo+sTSKqLpU5+D/ZuysqynFdH66WpgjXCU
uBndTgvxAUGuLieUfreLgXAowPFM2RCAF4PN0alU8Z5vknBo9plvX9PJ+KV7Klrif1Fp13LtBYdX
FBDZiTWyTtEAa6k3hXE1JlDcZhEdhTb+8ZL+Xxep/f0rwV5mPxW+GtQ7J6cLj7GyahtotBWEp9Hj
hshX4enB06awPP/zwePQnYCQpP/95BFihL3RqUoefmSewTfKZtfl2utv6F/RHkW7wxSd6nbsuqsv
zByDh3lQyc1tAM/KOdmLwXrqh/ZbdLRHzno7GHkPFdbskEhzat2B/roI/6or5FnzaDX68LvwUDVF
VJx/qXJOIsumTHPLY+2/sz2z024fWKFoKpeE1ZeLv6z1J0lLLBEfQazVLszDlHQBnk6UwePxjO/v
V6ozs8i17MPtMAM++/132G7LdiQ3SoPNIdIvIAVgwiMP9ex2SC3cvU2tm+DXkLs7ReITtwR3jh2P
X0Qq2mSHq4nlt12xirV34m41YUHFDHOY9XOPfBTKdAyMbaiWu32e8M4+dfDDwYF/IZ/NCyujusxt
3jfrIxr3/9DHCaDLpGjFeNq6kPGioV8DTkrHc0Z88GhjhLTCMKwjowNredA6DLe9X81kg/6b3J3N
u6Hs6W5ImYbG2Wt1QtfLHwlzUT+eFPHbZHPSCs24OYKENZ9dTOrkrOAjGP5/46n8M+fs8OVjsNB4
+o4vIhAJIDX89I9aEqywCrW5TDcWBQfrEiM96ySwXNQd17YPXisDARzJcXhA2ID8Jf0hZLuxGtgG
3jKnnHtZwH9fZnuGo3gjK0+mFtXa29D1OuV8XeFSPfB8y/pvEvwHIDilQP5d0yDR2TmD3o3lYzVB
Wl4tKsD2GAp3EYqtK+OsvMao6KboTK2ElMd3CsnaZszO3fShoe7a37CyuO6OMYMnGl22dPSUfbJ+
GGpdyNuyiCtp01y8cM1HZYf0uDYc43MYJQO2dyGq8kHlMB7texGWAOxf0H/juUCBqomj74/WlaIb
pvfI8FMyIxcvHp0ivFFmLrxLwdtTiAGT3qsVNlUA7FnqqYW4vE6tldtZKAsFORPZ9hdo7caJpMqu
neOlIILsKt60QZGuk6HsLgO7X+RI2/a/9VDTfeXFmh5p+jR49G3rgnuVurcIQDj5a6DMPyWi28GX
1lEQgxCnAFUYdZQJ8bOQnAad/2tkdonBp5yB/bMMd1ZaQSXKWJJWQ/BEPkCP+SUIbJSfj3LgQJ2i
/+bMYDTCkJUDaWTJN7KeQieUME1WaNqXXAxpzElEa955J4BczwIolhScm5GjoffOCCGrSgOICUW/
RR5P0i8yP7my6C57vvJ1oFxGimQ5bAnHrrrwHMaMTz8KrSzrs/+Xkx8I699utQLZIq7uECuDMwAu
R2CIkvA0I6fYwdc4qT6TMI0Sa55BZCj26AxW4JbStG+h8sang2R+8pRgT6PaUx3VBr6gPYC9rf3f
Qv2gAP4DwzBIW4ikKNHXu26DtPe7tJBV37WydKv9dJW27zQrNZODfXZEsiY8yTktIL48obm95Dsp
tZywm2Fiu6SSlOiwvNGi0oD1F+zLwkdPVDPV9e394li9CXieWGiTph+ravDRVlSzqovhcmUX6u77
+yLr0dBFqGl9tZF+jJjNAMg+/zUfjIaN55jgoKGNQdgFaQEYOZ4dQ8Gsj2/RANA8zBkvAE3mFlJw
ZZ7rqWLGvUVH1MdKNey6C7eoAPPNgGO31zY5e1jz/oVchCUP07c5eScZSvyXpoAqdWcltqAIWPxL
Jhnviax7S5SRekcMaLrliRk+8/P16Vv2y/ki4hTgDARFs2BpoGV0KPKT5GYpoAw3uFZvsWm9GiSR
i2FGSuNPdDKy7wsItcMvm71vssWzyK8cd1nmsNd4wO145+FgYz9mEx0jeZcX1DxTWgBT9Hri2A6i
jtvNDkgoHQXD68SbuXTUEXM1hD94HLFdvWRPBWdeOvfWvbwz0KYrsjl9Gi2/qG2nEt3gF1caECIG
1sxDG3EA/qP7241YE1KBBEeSOwDQXdKUEXFDqK3M1gVXnZDalGf6UJRgNfe+klzehlbayChXf9fV
Z84oFC5DgPgW1EwHgydpBr8IM9/3OymNybE/BHg5jwjVefHi3tb0PKyqUZFP0AgSonY97vKwbdeR
rUpwMPWR6pDrKXp5O2/xW2M5y6vzip541CjYVdBgRuDmtlLPqgl3ChRlwCehtGfOmEMotmdYr/EW
sxcpBCXJLG6FxEYqcO/6POaBaiHEno+xH2aWW7s9ynghAQw3x5mjgBqYINNLER8bhQCPX/i6h3Re
EoIQny/2MQsg4M/CYEbfBwYilyCyn5yESXyFqsrfhRZrsP9ZCSgAPESA0eCRZRknc9Q/rs+khewn
6Yuei2KthsirHXZLcda9+9/BSeRb9ODw5OPfms3R+wT6/tlR55hH/KwcBr0uG2ysJ+jdulOE6oUm
d4ngU/hFbGnb9ev6IGxyxptIxYe5D9+F+EQrhZWNFY+i3jX67DOyPSpbuR+anHc8o6AId8/bv0P4
k6+GFMfMhw7woErlNQAmiHfk8Omb+9VLhHYOnt21Ddxs/baTJnZLZF33anyj6OM6l/IJBOfHdCs5
SR0Xg9srDYUfOf7voK3fo6sY6cBKSidj7leAX0KCpAstJxanSPMn8TPCI875Me/gfJmk8V8+N6PT
T/sWv9sgyLcbQCgzYTv+9oMXVx/id1Vq76e6xQD2azs4B49IlnfwT8C1xBSzOwqjN8ti4NA4O1DW
4m+G+4gky/Wc0trOuzK6xQBJtQKV9tijysvyCQCwySMaNv04wdw6aKzquio8A4DwivkedIBgwqaq
N1OfdviKcM0Rd3yOYsdGLmiXPhulZcQKFo6vMhgcn8egJl6Dnr/ZbEuo+O/mzbJt/hzGqTDXMS+2
KkrxGk5L174hcAIEade2Gq8xvQDhFVXlKOIt5t37xHHbXALE//v4VCUUDFpERWH5y0UXVA8FSt/z
NBgGI0HDVOB2QxvKb/vBPyifgGt+upT79TOyBjMeixyiwxsflDWtYrgVHKR00T0ydB8QJCt8NTRU
caN0rnipWJUuQNShJjxoXWUDuY2hpD/E2Yf8QwCrQXbfaTprTV14JrJWvmk2BPQBrMslykEDHdCt
qI9ZAleCD/CkcHJn61LXEa88cRd1fYvyNBsHtS5r4qH4jIzDmDTRs1W7KlLE6k5ogt2bXsG48mBS
fbQGuFBywyETE1gwL6+HPXPiP9rN08zXqYfjwNHhvbm2Fy1YN9PgwT/qpLzSRYFfsGeeVd30aw5S
awIJ6GCeU2vESUTGtfInJ68/7JB14dYTEgNN9sAjdmCh45Yol4MnH0bC1T9fKc9/oKU6fjj+fk1e
nBBzeCxup82Oourn6ceR1L0M7540wIvMEe0zx7WZmpvFygKusJuPPYZ8PRwpFxSUXYZLexT5/ikx
KrJNrIEYPrmk2ub2c/Qu2bc9UL6lU1CzsroWiel0ZIR3EuCzJOQ1p++pXLkHY9/QtkSvFPf0tdp4
o3ebWwbDDjAmMsQTLLfg/BdCLL6P9XpItw9wx3ddl4QnmV7YbbjRvGf13ObWf3GPhTpFEvqlPGiQ
Nb9lHT2LKRB8dT/l6yFTWyIqedKIJL8/LVxjWOambzQENMxeB9e6eohP1Lzde865LsF8DqxNgb3A
83bkTqJoElQ6C26AKHIJUqPdamlp+QV7HFCT9QcY0/ccO6wkMf6b1SuYAqW3UFEKaz2EyygFR+nG
4VP0blJ3k7rRMXZK0EVHnqiRHyZADeHrXhwZBkZgU/wNnYyE4act7xbec0/kFmIAAN5OA5OITbsz
QVb8RUVBxTuQxPDvSaNyrNVgdhAV2ZV8cQXvAmEJJOqpIG6ZJgMMVFo/JamW2oQPEnprbBVD8OI3
XzHn6HfVho7gIxr5BT2JBvcZ9YkQy43SNqUwyl8PKo+Bre9EjSUWhZIvTGdKrvZZNTc+Fi4FAIQc
RAmo1ySdG4w5i+QsL8rvxU5ZFF8yj/4uMo7YfCU9HE2EUPIrRQOkbETNwYyef4fWEFAcWySqpypq
P4iK0HBjcrDNnpy0Tw5J1hueZa0j7S4ZkxlHOhkVzXujvMZD/mTqjh5tjiszSlLmQIXtu9I+8kVc
4gqOIveGeLUOLA5ZIoVfoXSH+MvDSTi5u9A+lqUHG9QxfEG+061GRtJHZ2K8r63+VzhuOoMhrJIb
KMesJxiHdJ4mF8blZjTGnRTWIvmAFf19bKSbZmdj+4jTgokkWXgnRm75t5UkIE9nZHND2o51gAm1
jGbpzIc6j+o81TdZu8VgOwAf7JZtw5OMZ884g9S3PC/+HkfaSNGufze1FP4X/OEbaY7T8rSq6eNf
upvUgLx2hemyXeMQBHtoUkctkgNj8ONlNLvJnFcAzaNiyGaNtKXRvVPn5hAhNBzRcdnlHfB2edIl
TU/o9PCfybMqtUMlT8ydF18ZN1/gCpe3LMn0YSsGwKCjzEfUjDdlWinFpbhOEJnHKXDkzZdo2l6/
acoc1soPzm7iTew8c3Ax8qOPt3Nnh1lE3aU54s3uN8Z0lhCN4OssQZxnKD21S+J2FiWFdv2Rs52f
fUqVZSx6ehka632zqUIw40OQKFsLLCJ+N9OM5jIKnShV4RTnUZWIV9wqOPDRywmDdyXPxLFJvFFH
VDBE3I7Zk4449OQ+lXZ1K2NOvV85JHDvc1FktdHRU26lIjQCkmQ0jHThCt/BABZwUCJgGBnJ2B+f
zgFzPGD6mqN6BNLbBfOppCBCMnJmrapHWD7/11eh43lZus6kTlTCB2uATvYwsGgb7rP3eyV0idSu
hrMPDnq14pQcA9rhcYuSvuyH3cDGf/T9nq+wKcpbz50CvyvGYDVpl0DYxFw7jm0+MTU0daQR1bNv
7eKFoy7umnsYA99LGNochfpvaPazcuSfuqVlh4bGhhWBsmpCh1skI+tEHTfzag6wBo4YkIulQIPA
R9V+SVpvuf7feI4di6H7vkDp8kaShoZdhL7zNfUUVPDkKJz16Z/C+j//E2LxErXTEDf6SascsSF4
t2gPTRK+CSBMNZB5JJvpHrneTGwOsa+8C2RbO29crVmlZzUG3ApJ+BWimi7vhHlJl7EeLFaW6Adq
2B6jhac6WVebQ2zdxZ4/+3h9LdYZhTFsJuKv4vuGRs6IFMJ1fhLjpeG40HmZ3ML/cIdbGF+AXRq8
6F+ciwXNmFdBcF1y6szMm6i5nG5ShmWGMGzt3A6cmnbjTMcy/jxeBTBvzhrhdP3GL+pHMc0mFrQs
H5aRzqDFq/iQSi/Z+3k9zPjemevp7isrEavP/YvXDWghHBs4Ei/hwsNcLN5OGIp+v2JmI6oJtKL7
UtNU2vR49s3StFCjN7CBXQLisJumgMwCvkZaiHLnppnp4EflVS5GBuXACcrHy5OzRKs3VV8KTNw8
Z++kbRVjnWOjPGHQf8L2/RpELapIC/1jTDUqeP301JqCWIskGigip2e7AgsSgY0blPRGRba7YiyD
s2ac8vpQOWxRoSYF/44opq7L7KnXrVZRl/E7Y2195vizaJl2yaRo1FJCPsAFAz6I9oaR3DegVmVf
4J2rv8UQ/8c28Ope4QHQ3m/Y3LzO2CXTnn4duHsrlxGzQaSSwm9M+7XPBK6cji1v+H/39SJw1Eet
0zdzstFo0ajVxhj3OmlSJ4XdJ1OAPM4OtzBdDCuurXthz8fIwWcaeIWQwk9xtEjT22hri0scBMwt
FyzMfnd42LkIoF7uOfWChhZRGJHgjkqydnXvAhHMPZ3bCcD6kZvZIQq9AwP/h36xxAwjXp8q9d1r
qX5pHhPj4Gwe/lWK5cw1S0dXbasib+/66TK4goRjM98Q82VcUK6pfu2iOeUZvLSLqsYM5npVitGE
cp+s8mE4GAjeCr9AMoeAwrRVB92dP/kJp+MNpsP26pAH+zaJqGsly6v3BEF20oo52g7xKWnxBgQ0
EGdSC0fZaUg0KCM/5dyhhQsCe3AYPX5o6fL+LCQZ1EgsYp1mcfCFDfeOjh5vWkvrLvSSjmdCSR3O
3uPXfYQ6bEjKfFLm5jYq3ZzWGbAyFHS9fKz3ZlAJzMRt42nKwaFquECj8TtHjBd+ptUnfcBLSnRW
ntc3d/An0frJeIcUFSms1C0jd8IzFef+hUO7fCpxQ6ACxtcDh3VpID9xJWRfV9IEZy4hLDq7+fW1
Bz6vmXOsbhpQQxd15QkauUy4c3lZeq9dtclqIjL7S6wHnLiZ7MRjLugkf/gwtUPP0Z3CLNnaDdK5
sVjKlUkwXLHdZ62K+v/MLrU2DpfMDvLV9QmZzHlUdPTL/Mb1FiviyVwdsQEymxepWbN8AB6jQDoL
Qh9gC1uVw1rOTn3BjI7xO5wCKMXCj+uCUZt8TNIepO/kz9YQGY0ScFrWzesk4xssm4XygPjPT8Et
ddIfPkht2o2dNSyfY8VE3vh6DcUNYUZ3p5jJ1wqV/Pk7159uQLzRp89ceMQ+g48DCnSy0yP5c0fM
UvBkYwyikUsLW85rPosHF0KEEJM5d9SOjt5PX74GmpVC6hkl8SpGkIKPmRmMiDCFx+XlHmj9dxXe
d1+aYuAeHiTZyLBSVfRI7/lJSqx5AFtC5D/KXrfUODN2VXL8/zqaHPsQtpC2mJHcXiwH9fUJK1lK
C7h7cJFcigAgJttqp06RHpyYeRJXVy23RAddHWrdLKYMp+lkr/I9VT1jff5ID71rdnLYCcOokye9
0PueqsCkPNF7J7QkdMzyC49hcddiiMpBvfYOt1dm1ddQdtN1b+rVLJxqpC5fAeMKepgQxMpmjn9I
/SlCiFYzRoOL8hWmPbYiW6ecH4DkAxPuBXTJtD4Da3w0Deadtib8vv9NgPuyuunrifUD1CPmwHa2
8jgYmu58N+lKOA6W8df+Y2yOI9nTJZsJWOU8aUGHfc7Tj5h+yGjZQPNoPWBVmElwAWS+5Z2z6DRz
yLMWoAGcrr/Zv8wr3vXeJSt+cm5B++sjakdG67FkAm+I+uK7eoQs9uNAcxH0Cm9dPcdZ9ByEnfD2
2pTUbqq9Norvc4xQNk7SR0MBI8LlAoaiUGpblll03UJethGTugsVUQJ1G2rAeOG72Smv9CFU52RS
O+K09UlhoAqJjpRxFt7qXhk8yp13It89uZojIpg9+0tOnfIgZ3XA9jmeSKQ32ZJlwej8tysqUT6W
3FYKnVnLBMz6kdbsk/3WGOvmq5evj1+JYFtIt0zKCbWBtSxXFC/942NLRpMrSUwIW/NJLvJPGSp+
wRNM4jzWuB43MGlI3wRV6TtwVpBp8pNVFyb7pbtVAXIWhpedZt79BnD0hfeTubJZnF+8s4HIVFgb
J1gADIWwK6DJCvMvlBWtBisBCxVHNGeSqtKmR4yomqGzscSRk+AqktrcpfPKnIsjC3+EHSxwOsRM
MDdqP3CkJXI6rXX/iGojV+IHqOWBlCK9hnnkkRIYqxKIHn5uf0pgqYw2sDPSWxS7fMJc1bqr4y32
1xO7d4Ct1HnEbx5tCruqTrdOHs3aaNB8nAePUIp6oRU3cr6Xx9f+m5BSX0lg047Ysq3I67pzjGmS
V9J6S2DL4Fp6qcp8wvRbjQPGlEUQdszPmPtC9x2DcEoRXkaKW1I7dlsDnntK92WTEUXVqclJXNdE
fM0seyWBzrIq8lJ//OUSgJ7sUuXy3eskg+3Fi62TG586GT7qjDQlPEer1x4TrEGGwCEzl9++kWdC
F6ppk5OMdFRREUFntwRGxAo1YMwfZGPsui2aVkdcqD1G46ZespB+9txMvlRvwGHZRC2YhiuVO+tR
IqH7zGOpBYGA5h7wYvybXCH/B29FNrmUYkaBOSj2MBR/OQCPT0M3tLZNyvrCRCixSORT0SFwBDb6
Kjs2PVpw425PzvPSM7n7PZJteRy2E9w+anigBLSF6xS0y1TjVLhTdtLCoAoS10v52D6rgg5SlIIi
wNI/RUzwyqBqQiqmNpBIDfTSE0tTPzxlyujDRfWEmkJA0c/zkr2yRnOngAUmNJlo6HEYA+x6lGwt
QyDCFpS/qcaZWSf0kT+oWOT1d38hZRl9m9/od3m0UotMY/PI16vglvtgRuhSoktnYEa7rTmoJRc6
yO89VPPAUEkWri49ytTVQIXOUoclNmCob2WfXL3ZMP/hxBF9yaQ+gLp4h0oxp3Z+LlLhw8IBj2qx
X10yFlmbkhWZrQ6fr3opUSjDEFdgRzNQVRWJ4I+E8b2u6apwcwjEY14VtTCQjuccbHxhaetE0eLn
T9qyCfFgFbJbpsYsU9UDoayMhQj5TZIlNqm58ubSJSuOua7V/f+XzG4t7faUvXIQzqLTdXU7a92V
dQZsz5cvI8hlz+5g742J+V3uAZIO60F1NaNc5YFRLWw92A+uykKiPH7zbwx5fuyshUVsHzsMHEqL
0ZMW6Ju2JTpXS4a1KddUP6cGFVZJQ3omyYUoHZtkn85y014jJP4SJchY+o7qEQBjg3AmhjC6gIaw
/PvmkkU4kkNtM6tvb0jVpo0LYHY138//0UJLAef854tK90RnlkBMpStjal3WBH+O4I6m7MZPUgmo
jajtO63aw2gAVckNiJ9vwdy2EYMGVDsSvYOmNBQd9BtvKT0oHkDCV3L/BxAtpn17j/bc312D86KY
0XDn6oUGGcekN+9xY/1tgWTUaQjb37yNWsBBWAxXoPpMqdRFjaBql7NW4aS8obBhxFQ6+e5XhZ/2
OvSEbY7Bq295ZkDDS3Kg+UlchNFpx6PfkIGjKgTym7hzwBOUS4dZhoRVoqF7y/iCiTXx7/VjE/6A
MhCH42LNMCWVqNCL7kCc5d/OLL3/g3lSocL1e5eP4rlPKSBQkd/VUPrHfVQqGF0on16nA2Bxmxs4
+q8jEn9kRD0oZPeJirzWJ0ylDXIzd05DPMhbmIYIlmPkFgT5XAKq1VEPLhsXddwGquHHkEpK8l/g
mCq11KXDusM2QX4rjZOZE8t0B9MtylFESvlvBFNIhpKsaJAirjO2vX03wz1YnQjQO2jC7OurpDZK
AsyrfYIMRkYTnulPAt2t8GfQK+JiOeWpL+CeDNdMhUnMFRC3NWUpuYG+QF2PiH/NBobDVXTAQLOv
Z1hX3QLWKXTh2uDIohNvnG8pQSt7VXsnd+BHOL3Ugk3NvTJK6yPypu8HaXBJUPkuyvzOiKShJush
QK2nL6LsiQQXL2M2WrHwTP7oH7Rsheh3ikbeZwqxMV5FtGAe1woZqskoc4aZ8+M2KIQOQ1o6uVYM
OaD3GvBXouWf1JqXeUQkrF/FmaYClQTtYwsQpDKzd89gH0Wgt+jhF7/uD9cr4n04BqxlXisL40Mx
ggNxNKaoJXPB3bUSURVesU0UPcrVaM5GRmVmjMA4tn0rFlkwER30SurUJhVAOx4p/4dbesvN8hZ1
580J3Zya0pMT+0zD5EFhJEbbCzWo4ismYHICsG0yB/wNYGDnJVUqWdiUiVIOlD+aXBY2ls+u3A+H
jgCsl8DN8Vfbl+4zXjSMEd0ErxM3EVeLVPtGyta3J7gbxN86SAooOiCCLj5Bp5MY33lUlW6J+Wpc
7uNQNtUIDyPDN8eXa15/NyZ4RXF971eDIPwl/NRScP/GS4IpelPW7V6qmeQe6rsEW+ExN/tk3G4+
DKPpFAX95gclwIReoURIXjxVMjyo0UzaJ9xS9ZaTOlLRidYU6nbckrrPIi6IVW38RllMhe48yhvT
hUL57LG8vdHH8eKGPDE/IKmPQM7yQHtoGJqIcLA3ZwBLetxTCPGPHH6x+fN3BpHvpAkXM2mIufBr
weiDDuSlvIXRrzVjJam3Vc3NbmMFqr04GC/X9OaGTA3fWnbwM7gEhL9rBYB0EAsgzExO4p9Nq3cX
v7TIwLW2YeJ+VmD+TEdvXc6GsBGiFjvlLoAcF70Zc4pgqARCtPdqI5CwOoQqLUdM8o5oQdDtqnqS
H9PqinNjLSAS4xm98FOzrn8vlUw1TBHtmdz3z4JjHe20OPoAWNh+In67LQrezH5qukPMPqmrpaVQ
lTq09/B4h4pfOMDi9tb2U8uYNcunY/xBpnYruKARbcto7CR9oiRUr2ZFXjZIrIHgRJvElfYujzxU
r5K7wH4eiIQIsz50N2TlASAZQKsvVuKJLBRFP2HM47k4o6ZQkiYw9P/0ElkuTOdxDGWiHE6BQbXY
n31xYli9AtHH2Guz81NGjDMGQXX9RHJkGINtxy8toy9dS8tJo4U8hhjRyQy8VC5vRaH4WW4I9KIC
vooktwQNCo+qTh5m66dT6defC1Y8DYfnnosbzf6aj17Tc0hDfVanM0Tsd4M1fY6b7jDs0VkssjTn
0WKeFCZx5atHfVhUjJxjKFfQCHB0UMbzPG2YO0bzi+Sq5I39NXjaN1pMfmxObffqNS/R9dNxQxOI
h3CezcP4gTSUdC2bfG80U/h2ZUlDRKxKwocZlTPwm3u2HzrZJj0GD+uZr68c/XhiIceZxdzHWFpx
bdVGCDvjHLbDDvBpZiRYby1eKzb+DTw/jgUq243JqFEbijHvZ8ZirXI3mX9IE4ucMwWgwaTE8ynj
98d3sXeRonhdyrYedAw5UEIrfaUJGoIzIMBvaInnZKSIjmy/GFpHAHdoWGYrLoV5T5ekHoPCVglw
ekVd//nxuZY2uNH4cB4vbL7gg1tuxBTAONPOo3+0pTreCbmKTLA2arr9m7XUItv6d+jRgAu7e2MU
P3lfTaocfq2qjFcg+DbgALZCEpcz9yMEolTDQO88i5mdh+5mDgAPm2p98TzG62DUjrdAYSw3HaGg
396GOPOfBrJf/SNVtH3lNX3P1yGUAazi6DeKdPFbj+b88YSNVbU87V5/KP9C8/yozCSDUQnTxdRW
Ny5rOyMrOld5v8j73KhWhrPAuuc7Iqf5RQaQfDdycCYlUQJJwr2HuR3jQZm0NrteSaZTqXYg1i5+
OD0cH7OyO2wntvofDzPrFDU59qe7LbanZg46RB9IP9TFAYd7tYkLLFRp1EcmQae1BrA5Y+wgtWtf
T8E1VYBXKpIqVX1luR349FIRbPDMcNI9fXtstfAa7rNwa6x7aDvgVGhiwmB/t2QRzAu+4zmUW7X1
WbIHtwCV4pjPguGvoBbUeyg4Jn8NeRPZJVFKgBA0iaHX7+OTLAB0wgtNhpz6ygGkOUv+FyS7bEqs
kL7K05BjUdazLwa7tqofwwnCff4e3Qpz5p3A0eFX+Hi3vykaxxfy1Pq0c6RXkc0SXZrKhW8DA0AD
HeoJxuOTxCUsqm+6KUFCiIa3d5e3jq5yQ7uFXuo9RdS5kToMdOd8Xh+3yyX3WMXgeSaC9W8mW1fp
/z4xKJ16OuFeL6LvxB0wwBbZ2GfMy7dM0omfuQMASJ3xSojypcexhKDTgyqEJE2BMktwcaApyd0A
kAVO8t5dkdGCGDWH1K41dDyFK48SlvUeuMZuTZVNbajA0gAwH8x1Q1iebf9Bw39Osjb44k0zS59j
ZSdo2P0gcf8hYmpZU4J56bDEf8OantTs9LnYuyQBbkqMx7B1rU2QWMrvWzkDvXgngK8buFf75kH6
g9k3yEgIWqlJy+wQugNTNXqvY7xsIexQTcmdI2Q/3UnZUx6s9fHWewY5dR2sOQZidP36mC+2eTq2
du5ap8xPFk+GFNjiD7QPV0IkuSMK1PmvJmnpTxVq3zG66l7cxWUu3K7ppST35c4GGzA9W2R6xCl+
dBsYP9Dk+Hd/WaNA3O0HyvW9k9YAOsHI5Si2ktIP+FOQ1V8GdTZBfWxhJPy92tQcnxwat0LLOx1v
BiqyCKk504DAsLNy9VT/iQRNIH8YcXtyGv+izFtJGRaKz4VsWRlAHlEIkeJEeHeD5+s28+jcVHwZ
JjijooaftpTRIvOIbtz5U3xbD2Hnt5PCJJ+W7c/G/ZHbV2PX4NK5UFF7PWzo+1JlUfZthwpcrfsd
qFThvDSCO+plLGTvmTQNeeIRpCAmTA+j4bd0+WwnL96aGc5d6WHuotwUuhD03lsvwtSBk1G/QHVW
/HiS2rRcNvYmjuFFU4QU+skiKxNS74TWmccqvDRDeByyLP/od+YQOhICaGdkNhyF2MWOteHuFUXz
Rh9sek+emPOh0ipEHOChuTLcMfm6nrut76sgp2CXz0dFUYlkG4ehwaO3lrtnk7rJtD5/3h8KW/Z8
RvkCV7h60Ge6qLVZdiFRNERt/XgvQIf0Eqkol9Xa6ez9ezlziHYI/RiMkiR2ZcnKEML8yJ3NMFgs
tc7VCDElqcUNiSm9lL5mVS1tB6NsGwSjIPI85Ite/ErrQ5yVSLAPIk7stiDW0smn0E1ow2lQ863M
wSK2Jyb+wW9g+cqJB9W5aSWRCRGfcpKdKf3klVMIkEyw3vbKjvxnIUxQ7NF/VYxQnSGI9bIfQFrj
8wtVoVI226bi8uCltOBEBsu9t8TxFR3TT2CcNqiYG9sHOl1q0uwl/eiMvHXn8n3f/ZfOxhZ/iNSc
7CxLQOMvX3iU2ECfcurhnktm3I4GkzfPLLBCb5OQTsW0EI8NvuVFX/X/OUOs/owWSTeNkKLFvCiN
yB/hf2DF9TYycSxJUI8Hmgyw+Z4MFlIvIyHHuVwp5eBibmFBdKr08JVUjjTRkatCXqE8HdF+P4NX
5sYyWYJkYnPF7/TL5Z+Jwnu1okmMuAJXKo/KCk2KK2HKLCKCvFoShTOWZJOX+ztXO7SYua9oWB8h
dfjSc4hQZPqcMXI2rU6FypJjy5u4IhYfoKLiAOa+BibNBe/dqPMBG4ZgnUq4gOQac3I2by5f7WfK
rLTkSdAjc0RacizctGzxTTz1VYXfWU5DnCG5o+etQ0XCtQrRpDIm3OetNLlUZt0P1QxvlCW9KHM8
BgHk3ZmiiKU1gwXMCn0DICoxlEBzFZQkfKw3kyDSpFPuZNrjR1+93OYXMsQCYbcxvhZn0ZTMnzLn
FqowS/n7/uptYMvyA0SX6xfzYr+RU6r3dlc7CH9AiYSmtBNNO33nbC5G755ZlpTvGt+od+zHsX03
Orgw54/DNGe5QkV4hxhKLd12jHMyj2hOKDq+nnya/CPkmRjfGU95uLKmQAezC44pBLzKrRpPQUuD
wypQg5hXNXDvI6UvlqsF+MmrEGhyYA+QEA/mwAGLH+pO0sLMYa+3VmxKBHM6T/M3Ajp8pG+PN3Bt
7/YbbsF4X4wFRlTRPxVlt84w1Poq+DBowT0CUdhXytDu4f75c1HMb8UCtNQgYR+SKDh0GxpqznRq
zDxpX8LbNTWCFCazohzqzK1y8DPuextRVPcK2TU90KNSYk7v1H7IhDx7qRnoZibXpNWZPkXJa1U+
SB2aF3qD4tC5jX3991Q618ImecrYhUxXNd9XAQySKxCa9HZyvEINzMmR4T3yl192CbiSZ0DG1DNU
3+zex9RgmbQdzGnsURc/lTPWIV9lpj3jYDGDfjCAiwy7kd4BdhYq7j4LKXF+3eKaD8aXSihJk7cP
vmacc9Z2QXRgcXPdE875bFNtjC0jKaJITXu9M5LKb36sxgjl/K3blb06iE8TfsmY9WuzHH7Si2HP
5UB4sgn1DDMVtyEWmt8KHVQ+wKfwZ0BejUx5oY49B5Gp0IJ3H73VKDz9UBKW70u3mCNJL1Rmgjkc
OBScQHVFeaIEcgVpRjw6KCSweIOEDJyuAHkOxz7pQ0t6WpEB35vEdkxRNingZGIe0XroLivz1PbT
7/vFibMLB1zLOphvfGGULQypDbl8M2TVvBF/G7PLJcSj7qjTTe3037GvbP34EaU3ffbAIPxAiU0F
8SVttZ6+5jL2QfENM3QCbW56ntPc4X6QEHqYDjj7cV5LB/xMm53vN6G7vhgM3bbRtG9PImOIRbbm
tsgHV5RZtNScrDZI2/KUYSTX6wzar1ObxjbPaPhYQu3M2E/4tvXVpv5BXIC+SPdxibHYHOI7rD9q
NRthCOUIWY1U8R0ewRFpnZANFZdvsKm2HhJQHNShUTVh7EjHXfeJ57GpldQk/D967dzV9MVLzdXS
jI9m43idkeCNXTdFCR+RzXe9fwR9DaIbtXxMKuc1igIgn0a1sbOPt+7k/l8rmvexNIcUeMIcCoYF
fl26Y8kQc97Y+qmJOV1En/NHBuy1tVilwEeIyJ9ZFfchUfl7HuZuviPK3sZvWwy0OZnsvnmZHZ3x
UW2RCFwK37/n3StFNg44xP33AHsJBX3rDai+aSXvOQ2rGkKOGM7AsOjtIrTyxiMG88hKd5cMXXS+
qumEyRpIBcixkEpPj0DrnxLOh1OskjQIuwQJGVOqWcrO6bPvipk1fx8lJfbMC2fYwoJUPiN7vG2Y
MfxiSQz2OyhFzcPfknWH1MyMrB0yQ61Gz3GKJ2mESPZjFcBh8o2amAqqX09u33d2jUR3iAftw0L3
pvIKtRb5ZTO6aodMmYPYFsmE215jkPJLJrngzPAGg9MTv7HIm+Oe289UO82cEyut5crwE3Nw5RJQ
tSIoONBlplzZ/o92l7GEBR1YqtUsxjD24r3E3fR/wDqmWV5L5eUU3vRgnwmtwcqtWnX4BCk//KXQ
i++LEHLyFMat/4PIMBsVLHBsF8+tA3RN2RTxdGs7nqGQIIoOYhSQfIIh6DheJkvj2Re8XF40pgyI
HojRvuwFMqp82SrKBUW1abdO4mSJCFathN/SAEx9Fdug2qO8AMYMZd0D/IxuZvhnIoAh9eazZY/a
759C5tq7D/0VXkhms5fkcUqJOomnOFR9yrR9TdYCOeB7pZ/AAe2DhfgS6NSuKq08mh0t0uNn+36Q
i1aeABnAarSRY0c9rDiO0rqA7G0MLhjmWz4m3LhgoZJOO0COVSjpJVzr1mvU15PDbDiSLQF9Z4bf
7No9qR6lGgciQTX6PzP3+lM8JgBvvpUmMm/JyRko48eu68FBPyqeSe6t6EXmCfXCYq+vOjctvqRo
sDWEzBYY5Z6bs4uzaGvFX+qQg4miPS9f5cFbRBUGNkNVl+U2EeLz/lYO9HmZ1YzXRwcg+XgATt3l
iusXGzP00VRIfrGgIsqT/82er638oOc0hVOBQQj/OplNnqX1uBRJxoYjNl54XulEf6J80gNxZcLC
4yjOj6vrU1WQfCIoARCHq4WHB9bNe5wXk/zY5qQbdjGlSClCR1feGCuhtOblm9C+RXkSPChUz5vD
cY0JYdYlewsv/yzG0fssvsAlpFSiZluOyOzTqoE/3zlGbNuoMJQytg7+lWc8vUnn1n9v1icSYL0+
tX9//SegXjx7+ZU302v31P4UPPapJWfcVMdnWoxPrbXXvW1FxtqHu3NiPtH77E7v5yXVFY6bKNcB
y/xMgxRH0n3O2tA6NdZ8Fvu9eJ2EbHyf7+VlcYOnjmoe7ESc/SGh2oLSVHf/q/a4ZqYTgS2E2nih
r5HZAQWcXKjf4xPkWRyqV9y3yE88mmj7nJbRc+u26jgrTVlpAV8vwgRhFLS7jlYuDMT1gpsygj5R
DH7MSQLUKe77pb2CaXAcmfZ2I4ZMdMQdEcNvHIAsKdP9xYRDF15LWEq0lLkI4iXH97jP54puHtRi
SFgtapoYe+L33wysfPFc8QNyoGnD2VGdCHFB01/u/jK28pbH3F/OLwrorxSYaWjlUsWQGGTRg2G8
RK/Ykr4Zg2HPNIw1D2ghlF9YN15nHahAwg6eaBc54mbnwhahQm6C3ABx+GayN3FgOZU18a33xN7L
YbkJ8rppe1BL0AWPbU65WaY+kmpvtL+3UwTxwB7ipcAYg66qLK47Qxj8klcuCpJ71vsastaR157i
Z8YdnbvIdlqMVGZ3jixVL9fBkUv7zJM0GXKpCHrM5+xJvQtJBQCUczd5b6v8vZA/VrdLPm3dXgxC
h4RhUefZJAHXXlIMwN56XTNZy+lX34lFAvafRNZKkUm27iHH+CNWxB/qAHCYbR580eQVOQQ/JC0y
vzN4dHXtI7ITJcY97suHMqV3zNx0dWuvJFIfvqI03N4tVgYopidTna6j+rv4NFoyeKHeTQgH1gaq
TxtxTPSa7pA/ILDPJX6T+viXcNG9iCJcJo+v4zK+XmXw9G3+qAVe0I6NHb41FDOdzyyxuufnwzQ1
2bYVwRdw+ZejUyyLR6C8inhVXGnZJ4Q3ZQWhecnUyjy6ileQGLYkzpXdTMVZYb20+sN/7lTa3yXw
JHJOQozxKCgrWiyrQexr6GXPbVOrlejYSdxIT7O3OqUSeHDUuSpWPrUqpNzzwmIdi71GjYhjeQMk
tp1dO3AKCYTCKNr2jD51c0CtNZL72FfOjbZiR6RtEGCNVinuMR1bHPKtjDrlpTqCnVCVUCjWWWWq
Mx6cttiIiFIoIsL2O4bRlztXLoZe/x0rSRZPly0bMcmq/RTQZ93IfDPrJfve+VxIzhtOW2Zeu5cD
8zsdm/gEW4tuvWHH74m4pnuUTt5no7mc1pj2/ZCg92LRhp5ttTXxQcXpS5X+9yqBSu15txi5Uq5s
T2WDr92MbmAY/09UBRb5ihQrnmLB9z76fC2yC3+HOVZA1B9qNPRHJz+D1zqr2B+UTP0VLinIKdB6
01U06gtSpq2c/Co94e5CmlDPQHsL/JmpvRb6qAhx1yc2+5rwU4hwZ3D7hOP3kpgO+aSWbBMZrIZ6
PVvKUTfMBLrqSHvWVipsa4hFyxcj77hI4Yllry4xvy7PSFTb5lHE0a5lfuCl/6ohkG77U8RdCxjR
Z8q4ir+ZIlzlsURsHWSfVGP1D1UvtZIm7qNT3RylflNH9YZn1YVpqsORT9kn0xsV1DxoRgucB1e6
x9mBsDW7PiwDJUPzwYDzOKI7uS0sqHG39lNhjbBaIMvQQqjK0MlKL8WxdaSKsntTc2d7zZ6McAeZ
ioaXs+4qOd2Vi+prz2LN/5uCQC8+BQbKc12WJTO55ahth7Ic0dcrT9GzFcZ9N/IcIkdYj00u3tiD
xAu+MJwkBwTbHWKnSW49a46bYvvXLOZQwQMCg4NLkZPBnumU1ORQToUgOjKDhs1qlH05yNtG/uR1
Ev8JU8AgO9WE5oxfSt1UrITYKZdhk7RzisiSt0EuA2GHldBVGOibxjb4C694Xnw5usZP0MfdEZwl
bATVyCpwCn8iAjvJI4KsKbORA9FMW5DkGR+l47MD17QE5a7fARoBJLKibvz8hwH6O9q/HJFGTkDh
OG9J9cpvwSnw+8hxuOR4rYzK5XmkDQ9QT/Qek3tiSHneLgZ/tEUTT2JsSL6uXJo/Lh4ygpaODofU
KIrFlZGL+PZ++3lvmjUL29rpf/xZIFCbU5791IF34Ulk7gmgD5TY3I2EywZqG1Zp48P4TRzbeBBe
F9/GyFYzQZhh8RBmSlLvLM3amwkjgBP8vbR8kqy8QmGf0SuwSciAuyTxSm+wc8nWHPMejnU3DH58
zI3+iB0tPoCadn2O5hrlmv6igWQI1O5CEAKbBfJidKU+/Z2yB2gl+qe9qFcs7VyAzlCWHTNv4Jhv
Hg2M8Rd+hNyvlgU0Sog/nLe2FOA63ONUYLr2VxpTLt+3gKYGhXFBo0v+M0lBQIk3er+qda9IuSvh
pcxooxLJB+n0f2Krk/LLGY0rdMiggtdOwlinrKUi4W9cTzeynSBuCnkc7RE6Px0xAaUgsQsHdXF2
0VS0pqeE5uQ+ciO/cWofN8C77fDEQtA1kqGI2ivmvQlfYOsjUwHLLJD5D1Ml2SdnF24TWWYqgey/
+y9889J6SfYXZQg65XOFJNLTrZCxmArS7Qi2h/YOFZRiWmGtDWMUxLbrx9k8ZzuTN1MslM07LJV0
DMNGRS8Yl57u9CzR4nW8ZshpbhN7I4yir+93ZVV1yAJwucdalHwRZcozvmQH3RswsnD4NmODAFec
EcqcuXUcvog1fl+zXsiZ8N0gtobocEvsDCyOn3KpnSMvKzLWFyilRdIT/WdJrbZnU9nRnJk7UbIr
qiMVv2ojBXsxkYJ6d9Zg3wq/yJsHu90EvnCwg6CVuP924GW0Sqz9XNW3PGomY0LVvJAh9LYjqGlT
16lILq1E/nWNE1FF7YdsOnBviD7ODU0hkJN0lh/sSO8t/x9CCNFJA3ZWBrJjrGr0CxmsArIvXeT+
+CXTMT9aGGxl/PEH3/Jfq/bH3DbNRzTA2gMyy0MbhN5Peika4CaxmcNG0oaaRo6e6Jfd+U8OXi5e
+LKH/oG8/Ug7WWfKCP/oNrg5j8pjwzRjObJG6Fxq9wBWG4Vtb22J4Q+Gn0tvKotnI01umH7DOWPu
H8Uovsmiz4FA1X3X6Gofgc2gSbQOHa81i5pwnNIkP97otNbTDN2FHusHamSgURCtwtXOG2Pb6bTp
fOSn/SYLAsTjqivyXbgTmZdDt/+J48avpN8mpmWdQjIfhXe0bu+IvmwXkpotuWDSgEppJLzJkn7A
l9Hx7pmyAucU9tlVsTRub3upLGRAFZ+dqWewD7Bnutm1VDPGKJxA3c64FhPM/Sbugz4vKWAkSE32
a6Uw5/8MCGv10EpG7fRJw/h3id0iop0+vHnE2xrbsSfPtOexqhohNpMOqBVkcJYejaSAC2Hw3fET
+z/buQmtoghWUBswZrEw/TdoEA2bRENs5IN3KP99NIt8X9OFM0DOsdytMJF6+/XO0B2MhMOqpOJ9
VKTIGO83UwRVzzLtuXyhRwVrt7vEUIUll8r5xWoBJx2ad1+nIh49P9dnaF8QgVHU5shG8rYgFrSe
mj01qvQoVs+J8Y+iq1Uf1ptmTl7dO3qHOFgfeOoFW88r+tfkRMDluU93MpHDJR70b8yY7qpYKhNb
14A6rLT35kRJTe2kumZCbIRLA75nKPV7XuNyXaI1j0OHqW/PBRo/w1QW7kL0QC2drq8mcqvEqCX/
kDO83kYziaSSz6sr7Y3x2h+Seb/pGvuV0acMufvIiCiUUmo5Lg5bF4YZrdffO53fFFiZy6v+fqoX
0jFind76SuzXkmFxaktsPB2Eb1hfGwHKjzs7q3aolBDrY7uQHQAqO73xg5IqFMlu4LSA2WQshS3d
ndmjgLpLCBhemu3LANpman3bripq4a7oiW3U8UVKdS7bpNJvghzBvZRhzPigW08GnWVPx1MnGa4L
MRt937roJY8y55bTr5jRnEB765a2wCkNA5mmAHqH12euPCGXIVFsu/Ex+TSjcbNSJovyPEaKugxp
7RYrY1pkF0ootdOkEjBTT/viaDLe5UF5DOCg6aPHi4I8riKCkdEcpiuNqDNr5ZwW/GSGyzJWQPh6
tjEk6RRvr0UcNBAp7SRBf6bEZdI8NoUza55KAepbCP4tmtuvAERUTjP5H+DdqYe/EzN9LprvAHkJ
7dJGUtYvtNnR3B/paMiFKsaA4b37xJfJl8WUon5kk05VbE9d2cw7jau004Qio3hei3ipxMeMHgQ2
5FhalRfSkrX5BjcZtheUSZckdoy5MSSWz0dyluYYv/mIGJdOABguK7z3AidCDiMa4gSdbokj0Y1F
oWTLGM++zePon1KuYhs3DuoLzO5m0MyqJwk8+vc4EQifUA+1OqiI5gITzesZErcAI9mtr9IlLOrh
+uhjF0X7uCbkOTLRl31s1tRT/UVltVAAoOt3tAJ1GoOcHzQVMWUyxsfA4cXApeQ91nSk008X+tEA
UTjwsxi8NhTPc/SRNPCy6uhy6oJCJX9KZLMUZbf6FOY5Nh8DNW9RqPCpldKcU46CYzSzF/0AY9ag
8CdDT21xdAMspH61l+XoOG0nIdTkTjPHd2tTgX5ew9ehkbZL8Ac+K6gLGmAxMZ0M/N9tVHMDe59p
2b3g+lPNnfg0sUot7ieaaLyBWz8IH1OEtU+MgTUy+06HQnvBg5wKunbSgDUlq4E2YaiVUhpFPgTF
XQC7sYxYE/ubtSr47gPZ+M2WwydogCZ+ZKfM3Gkhl7Cuo6GZ3e51rigfHan5W/ceoPu/iSGEaqVa
a/j5jy5Yw6LcpM0Yxplsq9L7jkxJ+ynv2cLOz2IAhX4/SDIP4Mqp8ubvm1J3ZD43Hi0IfFzmOGTk
1AtwE5krSNMwcMTjHiQJOEKsrGyIFHqnodgidqxv9b467vfoz2aaNn75nnVz/Az/hBseC7GAXmLa
vEn4zjNMGFd16s9mNpAcu3Ubv4kI6gkIvyeBCsZMmrkOy2y8S7WIWZUETv/x2BMZ6zN5w4GN5yO5
p9UObeHh4qz+/q0ej7YkHgYxoFIyUWc3t3d6rAkowZDozWCwO81YKpsE8xwuPdVY0Sp1/sCZ1qxL
q5BZZA09wUw6jQlWQf9hl7cdlE/Hdrsic96GJxQ8PkbU98cEn2VKgA2pcvf7s60u5xhZvoKLHfAF
RCUjN/IU/ZM36ejhzHrUamG/G3OgfZGLCqE2MRL+ICq6/sTWJj/7XAX0O6JYwlqBLDuS1v0ouzML
CjuMB00JVH3URbphuedOua5cEBGmCnirT9TNBNSlRs+JUGWPWlJFVXxuPRuLgUkvVHN3I1FDI1Xr
Cs5QVInmejTJJPnyN2HDsqbqnRJtcMmsp/7g+fVDuZt4OucrgZ0htbQId48oaiMt4NkEQR3D8xxK
/+G9hdiGwZYkocTiXwl6pG6W0G8d2GpvKQuXfynCn54IznoPUXGk4dSkdV4F5no3C6Xy0ian3f5u
6DdF5Ss9HJJpeWwOuxOYlkd6pRn9SZsmcnTbMLGbgdXyBGS16f+8uZ2pP+HO3iaxHzUgKu0L658o
Zofo1pXCDxMjBdjvRdmOs6n3YVlQYFz0BGaJzKspuYteRnLGCcYaI4AX1E2qzTPajdOjDGromv3K
LJTsJo8G72GNqBKIPJlm96uw7/ysCMop3NazWSJbxJc+AJdlArFiODOJjgxGYSNoAu3Mbh0ewlxD
S+13JGQJ8HTjQBjzW3mkQDoW2TaemCKxOJLUnaszOJsqCSRPadURlay8M0LhcXZAxIHLl1dPslmS
phjVUx0calvi3E3p9EfRF8z2LhC8R1Ff0QheEwRzpWW2hAnRtCaE1jamH+oA8XMNf0z9KR898Qkm
8pOrxpKTvcnZU+8wOnQkUY8ljxxTSIOGonbov1AC0DQeo0bNXOSrj3jdvKEmC58VSb11xZNrQyKV
4ORs/E9iTLNTD+7YRJuGvu/+dtkP4/o6vUodqaVwvVKLlFgxrBJswyLC2JQQQoBGfvUoKyBUUWsU
6S32eGfxp/QhHllqynM0dAB/qw1NeZnxrQpgAMy0up01QUJSCkl3vv3hFC+hh4ZF9WyqLQRwdqpD
c2knC9DK9Tv9BjCF5ugCGuoEH9GHO0Z0lgZoaotex0WOjfz2GOMCOnhbvtQbmQfZMnAQ9Lt/AdJW
W13RATynsg14xj1WPLFPOfZryK0/J6rnjOz2uQwrYi8FfWkziGijcADEGecRGFgG+uJieAoIC1YM
J7KfnjEminvQJjkYYwJMg71ayLtyBddKvhuNWWZxeNmusiJXp8oUx8j0KjbIa9PWHzYVjnnzHE1L
NfCYDXAdrxmEa0KP6akEhxobx7p/HVFYSL9VX+iSSIW7mkb4JB6QAKNeKzpho7MudOyfm5T3sNhC
1qBdQmzc+Wis3IVxsAvWaMcDlpik7VmzBB1U7bF40XTvNMNcFGLPMjwgfmyt7vz0nKtitXUa9AeV
iuywwp81Mp+Ht7233buDDRtFzsgupb/Os0XVErCOThb71XjXT34ANpn/3MkpLq4qn5FANhzukapn
O2fF88cTPrx2AUCaHw8Z4GpYSdst/txUDKin4d+bL26iuyqPfVL9dmO4LHzXq0pIOxRD5PXjyKAE
zb4ta/OkW6jVvYDP0694n9kzJzCc6fiUOqfPxk4XMa+LVg+IShfgExUxHPs3Gaqq/6yURvRcV1C8
8IEv/7x6OHzssrN+eTra3MmhR7W/bAjRnKMiA1exhpgIJ8e98Tq8oUHGcu4x/uPRYpdqrbvr8Szm
hl+Oe2rtMpFshKqFZLDbmNWSYRnd+1dzZ0GN+QnFXV0zkEYO0fQtOYOcSyQFwXSfdJLMdy6sXYMu
/bCmKJzZhFExY9ogSY4G2UJBjnbN/1AXCn0DkP/tyGwC5F6+WZaIUDSZpw8iVTdWajbgadJ5pIHs
kgZQj5rcU/XQ3OU7W03kuumRlNBHgu9XEwm6ZT+wYLTqp/8w09NLe1EQB2ozow7wxZLOv91e1v8e
EdQXCUHliFWNxekGMstDA6EyrDArXJWNZSfkOZChYZDN5FsST5grhzG8R/mxh8DlQygfxih+GH9/
WTDt+3hES4sj2tw2pTvwgDPrD1mchkSeYzbg1C49ximB2VADdUIS+0rifG4GGzypZh4dmYACU3Ym
Fcw9fCDRBJ/OWJsbrZ4T4p2p4cbt8Erj/rA2WyKTs2tdibWxn2Sh06P1KY4Fr9HtP2U3Iny5UOBl
dT2Ee+SEJX0gDiBOMskIpVLJv0T/5gpIVDqURK3X30SQbwt+I2Ke8bzf07IsZHTUwVuF4vvhrn9g
e0R5kYcG5gTOEOxNb4srOL4cWHYw4gZ0yaSxzGN1FL999L0euZ0nkH+5x0Qp05Tw3csCXqn4AbXv
Z4ClJDi+RBqLg2xtd1vNhn8D1lXrLuz3MBYj21gpH4oJzJNz8oPnzCzAaOBECCcKv3RfP8lJeKjI
ypnwm+NhGLBKhr04Rf8ccaOIpHeI3jOZJR3dF0ywu+VMrhBfRWMKhtIxWqgg6Wn00fg3N1D3ygm5
phCYn76EpIhI5KBpL7tn/Bmxp5rGemJ1D05/bMILLuQRaScJ44DfjKh8vGJufq2CQb7bbtqVcrrO
UuXH8mlSSWXSNqUVlbHZ/g8UZ1go3ywQWpbh1NyhreRb/hGh36l31+2I+IYHT5JH8f8g2Ry08tIt
yOGlgh/qa0fvQXkVfOTEZ1ffwpkSRsQ7EgPpFnD2JYMcB+/njLqtW4RJVK2SJLiCy/Q0CWyeuba+
rWzEfjgIBj1rP3yPxf5cDCwUHc8vlXIs29wEmUrv/XE1KMw332mb1kP6kG81J5cp+egUWT2ZmJnT
5TJVdanmxQAn3SVSlxC6hRs7Qf5vaPcsRkfrP3MAOn4vkUCCKMju87/lZy8qDPZVa7LlEd4NCNjJ
lsRt3FsyyWhHCoUS9XOSf11CEH0y0ZXpvb2oTJpwr5eDVayTRu1nFTfmWtvqnjJgH0eJEgdiU2x+
mu0ZLqpKr8L9jYS5hKKEU/OkAuigfg936kRGDQxxSs/bYBMhVJHy6ZkxqQgnjW4mJ/FpI62zxG/q
9Rg0kEI75nizjAuCHWkDJdunHcTYvq+iLZfqNsCs20gVsdpm6pLY1jBZ7VIyL/ojQgA3RA2EwTNP
PjK1suzy+cUvUWkVkFUNyXJcqBHY0IRnpHKVIQEfHgBu0ez2qQj3R7d932AzJTLwP3b4V2HkE0QP
N0JE3LKQaUPcHHQXpi2I7w5NUcDlq23gLU/oARxxf3c5hBkrHcrvEPj6pZNnXJ8Zdz6G5Q8HJX1A
rJGTb9BBqhGyQb6koiajOhIH1MWtLn6BE9lGmeexiOR4Xt9NUBHli3k3qxt/x9BdcZyalJByjiup
Ho5guupOSSATiedwqBeDMjIizue9iVpyANZ1EWQWGBHukNk0CDTNNUKGPOzERAGLO21O+p9KXnfC
Qi3Fk+gVgMqGhmhRJhixaCbwQyE7ZQKXvcwyhAhkWImmpjx8BANBtT/wfj4YzaYqY5E/Cj1maEOv
xNlM5fOl7VIRylNDk06N7EU26SbyUJsVKqJ1GPH4hUhulHqztAheiWNtqzdz1Q9em602ripM5a/l
Xe4igVyg63pRTpVzwR5HOHZ0A46g80DykCVbQ7YwMV9jXaBDPhkfaLd8hIXsSEN6YZJW3i9qk6JQ
JlTgld6YK8xjOMwEjgocFMjFlukStDaqM2FKYLTZejodmrp4VDpS5MaPsCAQcUsRYdXnGEf3DDjf
O7rD/VRjwSXOlUjwdmkWcaLigADgzCXEY8ohBjy5aWTbqE/OlVNrKf0xORoFmFcMhuuHLXXW+FK6
n/6L/jTc6D3hFP/3/t6ufNL2mBiH8piVcppuBw3l8FW+NGj138D1QPA5Uswvxyyw85vd/JwTSggT
nikB0Y9G4/xlzqahSVTXlBUEnu3Iv70i5mTtuEBB7krpRsLOVPHX5g1CRUd+gcWKdlOEpFSGWIrD
ZJU+A5/+SbgC+dki690wqkKzUYnbtkyKmPr6QplisjYAmljNhKC2SdWZYn/ynzNDpCISnlV63XvN
NrSNMrJekaXysvjyE/UuAh1xOt33GNjPA/VuduyeS7VOB9hlAtXQDGAegL2Q3onC/o6Vd2BE0/bM
LrmziwwcM1QaY/B2EfOuR6d9GewAXpZXDfpRnfgcDvDcXFwYn2n+Ekonz5yIkRJB4lO67VkQp+0Y
w6wD3VQ5QwJZ12yUS7Dgln/8KCmqnKRBzvJ1/fQrrbiTh1sXomWZBI1nZMziaR+7zZOgy9kz87XQ
fZiZlEw000yALGO2R+4Jm3oKvkO/VfrimChsdIaT/Lt+ngON/8tK66uyHLK3/DRb3H+3yBPkLFhp
sX5AGONaa9YsnYf376bDP/sfgfYru4EVQtvBfD1JctQ5ibiXB9gurU3W6LCmyUANluOxnMIteUII
XvbNTHq9a/goqQXkBLHfzO1is8oC6RFBRxujgnqFJ+meBlGjFr8SvtLPxIBYwxcLVGxjJizUXVNA
sZ79LHLJSrBKxxFz8DxVECGbdxo4vRD40xNUGKfLOXhk2yQ03cSG+84ElHWRAuEm6MCjKKzEbmOj
fRjpqQ/zszig9zQHGqfjrUnesnFaXxCR5I7+irFjqewLgsN1a9fbxdJq2eRkYK+fqX4d++ZQYPWp
mVrsA1r/XUUbtSHfLbW6UiICMGUmf5OvKELyGw9G7U/5eW5hLh+sqMg2bdfjvnFe/n6M0icCkWJh
TZimsUPawinbAcWvCad7DspudyOp7/tKtZpbmyqnq9hASTx0QlBEkikaDDGXqPO5Pa3PbQLAyhsZ
Wsy2s4UbQdhx21TISkAi9lOLdXp2j0iNPBBCcNDjzH6y9tZJXDSLFq7hCKo8zunqhHqmNcJmvdr8
ewvET5OlyZrc1D9vVhuU/bQ0uquJCQpzh8ifjiWRjr+8610uNTsY/Fc1G3NgIOEg2Ercb0Sr6cY+
AWu/K6BjHd36ZhBoK1vktT+md02DLmIcylLzFLtTUYnwSCAsag5/rg4ZUUfS+h3Wb4R0jNQxR243
/UuAKiA6s8TlTandXeDJ6zmBGucXfKX6oOOFzzPmJLf4Ln8eI/cUxN6WOv5QASjLF3H2mWNfCcrV
F4lqgPaFnGbjnWy5UdjstwtPsV/wnsM3Nij2DmsLiVF4KAjFkEHWH4gBM43e4SIjSN+y1cSuHsqm
huP1lkNP6AOAdI5bvGwgtbOZ1zncrQm0ntuaAcaleJFDjixzxZs4qgW7LYXYaY23amZLW0Wh4xCM
iCsk+DxGtVoVLkbCh2o8vUPtwv4EIMt0FoP1jQjFaewPD5EmRMStuoOJ6WWHuOEuDXyE/OcHwiF4
zKU22IY/SyUarpYqR9YstBpKJYlM1xrBDRCu1c2wPUm3DxhefLJ/g3mkmsS5raLcBt3vx7ksPacY
4cHsLwpC5erA3Bw8k25u9WNGO0yc/JkIOEwMv1qK8A3J1ChaYZzdKQcRhFrbLjzzNLugb+9iiJC9
k3gRAFniDzBlCHacenr3eaUjYqFIBm50rp2kBLA0yydYgIyqW4ZUPzWw07hogvQ+edzDpHXH/Zyw
du147UsmjSpoVpB5e/uJSZo7a6wk4/604DTf2SKfp7oW7a9fHWt+Hs4VuVojdozXoxFKkfWVhNAW
OYMQGLTPzq1iBDfuXi+RXh1Ad2MQNBqS6Bgj9yzEtCJ1dxa65A6b5ZMaDxId/+FYjKHUVRNir/Iz
PD73dswwMqHNj7Ge56KBjh6owCTpL2Pyg0SvCw12ihzVvJaJHWoAZDKslzzo8/uN9pGc2SlDyKok
Zg/zynIk47c6jVQXJSWnURku0Gd4JYRAvi3d09s2a15Ju+/PBKNGcJCJirvURAy7SFGNrS4aX83E
Gj/mgE1T9cjUOmPHVOXYZCmjrL4VsTtQ8/vF3bKS5Ou2sDDmZ1T913ugkc6j9L4sVpVkmjeyUSPx
jUi5Gpha31q+snoeJHiWmEzrN+4+0Uv1RN2+AKQnvy8E2vZYCEYaEnZhVccqqfrp3AH0p72dQoAJ
wPcsNPfFl6v7DsBBltrAYxd+qjfiHZfjRaTnrgaFaEkxLYSR4QiKtSgZ9FVfMqHoRP2grOB58NtS
AXf0HjgooIHPUaIuR1bgfB4kIOSUCnZQjyjGv807eQAJgvHgvg+CjUfBqUkCb13T9LOvYZ1w+l29
uG3S/54NxBOc9Ozcnjh3dO1yvy9mh8MuRtjXEuZ0RqyOu5rgtOe7QPls9lpaljeeuowxM5uf17O+
xbQwbbuJPeO3ZtxJU9bBiDfYhzOqLFbC7najtnLKCBgAyNaAI55jE0ZBIKjcf+Y3u63WHIJZGMW8
PN1q/f0RADCKt17MXea3ClGkDJIKGq+0qdOaUuwIwc9YuDBLBTrn/gqFMHx4z51MUNuf5DawbFo4
9EeyLaPR/TZrlTQ0Cdw/eAJwHFtYEotYlNazbUrCZXqrXksYoJPtRFvCE3ItX+ykH2lYmbtvfpoB
FBHBz0xYzMoghuroHeCVAyD8vumvFjUGkDIxjMa7cZaZjqNmpwGEmzjLFmJKqp699B8tSOQzL5NK
7KY6f4P7ONhaw1x7y80o5BuQ38GuX4HvGuw2jjxzDdbUZ+stRjnb6sS3wc68CzgoQqHm0bSQUjH1
qiy0W1WJRGzzfmlnMfFWlkXbDFQclCkxe+apfFznwcd6GiPRmHNS9QfmAd6o5Yx3zhSA5Ynb2Oih
T2I8QIHwseqnmDk+2d5Pa+vTHDOa3BMl5mFMvPQPOA/mjMUthowe4dPl6C5T+YTl8exKmY0fUisY
z3tX1XFLKGt2/pDkJOXguNlpUcOPmnvH9suROjE8J0FzGzmuOScMbeajGmh3N2mUyl/H3Gh5C0tV
Dxwx2B2qtjUQgEWcXYxi9aqbC1VG+e2UOhYUQg7yHCfK+2gl84QNxpBAfLi/R7JlNkJtI2/arbom
L7Je06FvCxvp4EvIGk2N6+ZJGX0wRdqhY8UB0gL1DX7aiG7zEFpEiBAtWg5nSSe6tD4VoQW4ni9T
WHCbTZrPUv8TV3pmJGzjoAeKml3Dq0tBObzYAFAVFu4s9oBJjWt0jqXJY5thTiwXE9a7NiC5G764
BA7jy+71BFBSuJ6c6BGu+ZyqohqpFAGVGo6+PbBGFGBX5bX0VNkKUo5qKayu0wiSytSyKo7Ow05h
nCkEiaVA+cVWXKAgxgXR9BWyPuGKQtunakirHqtc1hz/t9yUXjU/FfRmhvCc7EwxeQ+N7lb6+RPB
r7ATrHxIoIK1xYZYDnPh9ngITOn1e/iJVUUXv64bCOnMya912cyJJ3Bg3a5zLiwksguGRagO+5nT
RrQTLF7BIv5qmd0WZszUxTaIAl4I+eQX3VSusmP8EIanIG72zflfXYnv2pa7Rqvp3aIkb6duH5/C
xG2xDFAViDK8vU3V+EqJ46fz4uXyagZtw9Ak3A/6SYh+hISdcFPwriVOAnMtiKTYNitGDuaAFdTe
+k3Po/OyEmbVZntk4k4GBV3Rq/I+prDuDeSknc8hBc5w9P0sIuEYRyD8qscQesRU3wIP12EOsYEi
SCrYnLnOikyOTvtfb9Z5XBKp3aUNnP3qe5Z4PtPiWxipVmbSP1qM/npJrgxJIWYbra5q41QelSip
Tn+pabGY1fb47Ssyr6nElPwiv6IAixqZkfXWj9Jl2DENO8JLJdCv0t9x9Pq0QTNAmBwoFMyLPQTJ
Nq3ToIDCx36rmIWY9D4+SVoBkcukC1yz0a+Rrk0nG28zIdRLkkAeaGIlQhhfas4WmYxhRx/WF8il
f+ZbjpnzS0HtkzM/dM+waJ+GU2Wf5JuBZAkMMamBHx5hmV3MfkK3d37b392GEa4JEM3WyKHQkjN2
JRVgelTenwN0LwXHR8/8rvj5Vq7gUKSoKAwvsOH7Y7eM20nmTJk3KNIrrralvnJF++sHNzgBdWtG
ljtqBjQN7XvuIG2pBelGPe2PixpGE28EJEXZewDQifZ3hYW7aToe3CBElZ3d3VWV0uE3jtdjvqv/
5JoiORgt51/Dc4ZYonDpG4zTZtFosZ4alYrsYQNAFppkMquE6P4ZBs0nG++0BtFcw0pZzi5wkwOH
Kd1VmX23u5plGMjxLFm+ERujuWoa5QICqiWmkx5g73kABpTbjAtkCLR61MuF3tBiErCjvNXeT6m9
Kv2PGDoROojaHmFrY92xdvoQaGinYoguR2z0kleNmlemumQprH+TndCjyrGLAdfbHEY60PBDoKQ8
tgPdtdLqD15jw0eZgkurr2WEzR5gjobtDSikf9cEmskkeOOwSlzTVXgoYgWPkQUoTEy0OCVfx5Tq
LmG788lRUccajnxOiHixfGfHe5ZkWnD7TKy26QMF6K9NO2QqKgpvbMz/6FSjMgJsBa9WnbNbFFFr
SZJzygU2fYzP3tgDCY17BcsvUGYdIMTLwUD24HtApXynUtq5iJP2ap3ZQIBvaVvipb+R9bt6Os9N
NsIsp7ZM/HmSC5CNbwNpDVZe7/acy8gwgobxT/H5A5mMuhjcGWlkUvbqBff9Z8STqOllhLOoak6v
sHJWzhduIs0rfh27v5YLKkVkRDmz6UlL4O1m0CJKNZ+q5Iliq0OjdLf4QMPSnKaznH/0mGm76ihk
FWz5x8LSvcl+JL5862hQIMZy7ZDp2FQyIXaJd2W/3WAniSJtEWJmcXIHqJETe0kWtLXjvf3Od3rN
6ythkcUVzuNS5D9AQaWTdz0bHEwK8ctue7jpG6Pz2nYVCdr27Jj/oQRH8SRiETmJP3x2WzyU10Kn
wcsPx1dTogYzxlckSKPdB97Bo+2AcOL2L22R6f6uSFczAZLbB0r/fR1TqtkcAWXyFwWGG4eme4c/
aU+obF+KeAm8nub84vtidaNME76siG2XxsH2IS+tkwRVSGST0db+8QRJMmfpURJECiAgsZNzD4wX
qnbvnRS1Ws++50lXF2rnELxvSq+89am2gzZRyyS4mMUnPAoMgr5hWVlaH3rf3eRDs78w6+ZGnejT
ls19YfvWQ0hd157vSMlSdA8vRsDtI6NUHO15PmYtPlNzy7rg31B+zYIrP5d9qq0jdkc2WdMzSl2T
wSRX6BfLyd4MXq4LpQcLEqyyuQ1Kz94xFvHKhLCAXamAIiB7CgYZFgbGOQAA0iQS5KEsbRChdmHt
J4A1/G0CDWaimlcoACtO/j2y4y1rx3VpyN5VmRQL1p0lDSeVtUphQ59z49HSxwqF3rYzS1/l9RjC
xWO0qYLolvPr+l2SOKHlRK3LlimL7l6bLeI+RLvG7SPnVA9iKb/smKp6fT+SCIKaeuTo2PlNGMIf
Hcp5mLSLGaL466D971cL7clrxUHTIAWjiKCwdx2sV6HZ6+WnbxovyRDfCW4OTGLym9KbqgssdF3K
22HqmpMBNhh5Ei9X98Ps5fRO4fo8yFGFdZE6hTBflaJcubHH97dnv93gRFwb10+/JcYt//kKNWBX
GFfxugdtj69GyuvRR4o6A441JWZa7GGLsSVzuwp25iaIZtXh1NefAn8HI9YWXS9GAsJqmeju5S6P
3SLLJDheTjCbazuP1wy4GL1srdHEgWDoAWWW8Fmx4x5Tym8psXDSKXQ7nzT1qhe3UrlQOURQ9l9W
kVioQAqSf4T2EkRb7pa6bGGzKxQrv5LmW6BzmPUHDExcRcle1GVctsGBUcMbWEb3221iW3wNPuYw
0pGR7pr4SBcRL/+3D9W7gfn+vyTwEjaX86SJ+ZqC6NQEU7oX5jBgEho9Y8AqO0mzypf1ZnQNjm6/
l/uDxx2f1wu1b9SIs3d6ZmWCmS842X7DNRrTjjVmY8AJ1nWiv6fGF9P4Y7nPFq8N/vguctalHgr2
9/KoyuS3PiBvzfS2kwcHL8thnH0/qtpTjFE/qQP7DKEP9zUHog7ZSqjnnlsZVQlmBzTLrYVqQy3R
NGBdNgapJvDFpw3D3AcumLTl4Zj2fZeRRmsuy+X8WShIRHUc8OKjiq4LmCOpu/zic5JNA1c8ekJB
GvaYhIJ2KD3JnYy6r6RoGjDqTb3orhqhqhWNc+2BiO3feEUgW36k40h+eXeOUc5L3X+YJgT2N3xI
QNjzDNHsu5G0y2UY6aShV9Wgo0KzQIIp2D4wfzu9eYQn3BTxKTJnMVTfg4GFt9H0roZ/3K68UAE3
J6DSBZXanJPcw58tjAifLapKV6ca92g1gR9svrCOzLDmZyOs1xGJlLq27FGxWLGOaNz8O3zOC/wV
YH0axZSPmhpS44jVoEyniM327G+VDDh+8g3QQkuRtqo3cFSBb/n3nnxiV5wWCCxnj2TEAm7HCWYp
LaWsxLTHqySEMGDVjPb2DpfFa6bwwSVVhpX4cE7slkolCTFB3VUgO7MeMsDauWWMLgNTq0Uf4c+r
0Dnyj7HsCRMwr29veKqDXo2vx3Q8D/r9SsXq41nz09ZDuQeYIpaBr5tTH9GYK/7goGuTzKG4Pj2t
79QphHcKvp5xWy4z9u5oEDARY8hsZ2DiGE4O/292cq5RLOp8cYDX0Wj6oI8GyFgcnR3mRNDdkx+t
d27HB0Q06WErPuOuGKhz/ujUiM3UITJRVjWjwdpxwVBCJ/60aQX77xalv/mgXD1XMDpVCnPMC2Jp
SfcnYRUV9O/5oixjOvA8zZqkDq4r5GTUdl0V507WoX78lNrE319kXZqZSmi2xuBX4H0Cq/0yfd0+
wdR6l0QK2oJGNdpIzPmKk1RLZQ+bzAzbuVjLwhCI5maZqUKfwtZjChI74t/0dL0HQptfBU6/AC/a
9Fc6LkrbZWPGyCENxhPmxyDeN2lNOIizb9t4DUoXfFsxLW8MjFU3DOcroV96z6XJkrAem0nB6xHp
TIG4z2d3oDReyiXQj+C/WVhCF+vFUb05U6REhR4RIjgjh4ZEFHEoY5tw8domI/yG77jdW2JAfXZy
2GGL/1MUxy/8diwev/Q2ZeGxRjit1pcOQ5xZZksvEhYrchnFlOFC7zQMfgVqDt8XGJn1bAwsY/lZ
gvxUeXho15wmg7+tKjD5qYoSTVnOFphEEYbpW2Ttdb4kwoxQQF5haY0M/L2h6y7171dHuH8M5bR9
xjs/yI6soCwC45Gtc7CLFcnHR4FXcM2d8B/7cvlgNuREaWiC+Wm+gdzK+cGZgnL9zZqwyZWZXh6m
iB0yY/MsGOYaq7NXK7Q3h/pX/l3wzgdg+JZqxe3ZLRMipPoZ6KZVxw0OxcpcEVaCyP5cSKQvg9AD
+dB3v9+FRrXaMCfOfGuCRpWKzjzfvzC0D8C+30ixa69edp4z6jpfWez3Ygn0hKmCzWWZfp+Mq/UA
k0I5X1yieJicWuQcCedfxTfEl+6T0KxZHIwZ3IJvSQnc2R7G0IOLhecQ2EyBaCcjdxUzpEw66BKm
5Hnt33lImMdB5i6pdFcWfUecEPlaLPn0xKxvxSBrYru7Rs1VxX7HVYgMm9RIkDI1RgkU3/CWxUkq
9NgwiVrrlUvahpQ2QMnxEsF5h+daZRu+49R5VD5Knnd1RUld4nlYNoSuoKga32CTgJsiBHuq20Va
QEhxJ2G7HQXbdS0IqKM/sEtOvqx8El7mMNDsdyZzVlgHMa4MqnWlgmP6p9NaYvHEiHBmCn9RSXO2
OVz1dCw2cDp+pbo3FeTnZM33ERWcwZsEQQQZBG2q0RtjgTgyj+pkjdnDYVIJdOoDMp8NGTD0dXYh
fPD2LVVTrmG5waXPZhEfD/H5qKd85tcOb23itRsMQIdW+mcrKtZFoyDBSSV7d9naU6znoGoTJCuG
x2dw8rNPhKitfIEbF5mYiIwLK612JsQfMpPO7OU55L2z4kXa8WQzzW+DsCeINHTxZo6EBAl9IOJF
4OA28wmbqIQrfa2pOErsgpYeOjRHmBH/j2VNfR3dT751LQR2E3gm/g77cK6fkkJGoJb6r9L/qAXn
xhySkD75XIbQlkFx1mrqPK2ftbxCu0/5SLinIArA0g4dIATw3GySrdVa+jNNDG9FG8v6EO71nDKn
ErFk5JrLhMLLA339PVgNgwMxuvifkrvLYtfpBGHok4Xrk19+DcKGiQ4spz1eTpkUuEhYt8iLZCeh
6HszwUHVAvUbY8tfSZDtgSEUEa/A4mqWLBJM36bUK+PCy4Te+hCgIRFDp0uE4nH8Qesq1Oy41Ai7
GZ9vujGUGCzPLt3DkibGy+gqIthdkWhtd9dZ2OzRLBE89bfDQQITUWGpam6+15yfrvjPk8VjUdQY
CUAMmRI3Qoh62yQnbVbNpftUBn3Kb3BzQ+eTtF7uSqkL7F86/EHWuL0lHHzhljqxKOXfiVkuMM91
D54+sfzfoOuh4oslYp8mOXPeQP++d81B5HsrAVYsWqaFkkDRHUoMOlFk309F/uThe5mRwGxR7WHO
dj3gvhf5oP+SAKy0D6780znMtbNBrlWxWj6WZw0hcIfze225PSaK7U9SLTjgLLT5DYsrDzk3RsqL
DdqCOiCQbuFWylsnKuCLYzovbSrvYh1AW53QXVIKoGNUd2QKC7ijaQOgpp1Vhf9Rr4MTolCrp2Cs
jKscxvWY4+I7FYtlXxK8Kd48Xy7nhCtc4W/aiNQ2fLy+CQN7U7Qyq0Vc7WdZFb2W4/MR1CKHm6tG
RNLz9/MBELNkQughKmTDyYN9FYkyrEfL1Wu3zxTP8m2j70uwHTcM+a8TWOfaPQzQrC2BSkb78eFY
UH1yLAma1kZ0pmMZmrPuA+5sT6jpgA19YilnZfT/hj4KrvZCefQDIYGGmIniIodvvFifHDwsvGkq
fiE3j5a2PRn7xZaT733gqANDYoIlRSK0NBA6JbYIxY77WUduYDyc3222kIkP/smiPDBdRFT11wA5
JuvZVMszrTmj5V4CZMIwKs/ojarfOlHpyOyQzb/fzhRTBDNAyryjuH9U799pgAPdrHzKoKn+Do3g
okANndIMrWmqPLmvC1RnJ4qI+TImlnliSc/DEwwiFWYsnqVi2Ng6uxzO5OFt35HzNHwgHVNIvlp/
M88z6/Gy4VUQyjxRbxn6ob/HhFRxWLMOPrItjGG538MqMnQZ2zBBfCQPU53Xmi6xx+55xYCDtpAG
u4RD/kaLNUHRhJpaJaCh3v8JU7h/YrqdzZ8QTcj0Z8tFbXRXadXN579+Ni5jfIhq8ErBSQJ/D1Ae
DQvjyElTnfv2+XEH42JJk+bortiTMj2ypdiZsU1gItogNFT2j1dSUOSqi75DH5KR8j18dZOf++Z6
7EY3UmisWgt4soKq47+4tsAfpp+PSicBeN3M+hSQNn2BAUlN484BiA51h+7VmYRilBlCkyaFyLET
BodSTVmD7KptxZ7QKgmZpRMwRckzpsAXH6LK9OYR0rYx2mDrLFqXokR3PNqTs20k+1GGvlT3QvyL
cOh4QDrukdBBXzqh0UjJA48LJifxJhKWQY+TUpGR2h0ZgjIfpqvn4VveJdYRcFjX/8sjxKX0MUyB
/YeW4DMTGM0hL31jkamhyDkPai86L7Tr0vO6MwGDtFh4PyJKpAIL2E7LsDliE/I+yGIL+67yDdcT
ch7UyeAGJpi0ickrvXXOGPRtLIV6ZvE3yEDnSYcqsp36duFPhMxgwHuhc9ks1aTkeKi8p2Kf6O//
QxMlqwuc/7MTCQcXHoGJ3Z9wKh3dr/tsTHTUJZRrnnWjzBQ2YDcpd1LHcy9bproDqvQH5FcZpywO
zusTUa8BvdjmCU7QqzgQVjM5hB6CaPNp/IhcOwqqc38P1UDNtHKaHluqLqbjVxxPXAHTuoxpnaNV
SgtcU9pyBEACQZGRH5g2GxbopWad535SKwCwd0adhhFrMBE3XPn0TUb11Zb0e4g+XyVdyKSqEBp+
rrO33xZNxfQO99BGjTVOckhDk9LuuN6Pu+Rd3BcMzKvqN3v8vRaccCklRvRiboQMnKSMfcA79hh/
5zfwgEFmyJ95OziIzGeToh4LITxxxNNOKdZwLG/ejOoYyaMihi8crr1UynTTUDlZ/dXS7sD6ICIw
GeQYeK80CQvtFc22QobbDqx5O6josV7Q34dacCmcGpc/UT0Ky6FPl5QsyVoCOdI6rAa2SrZmMTdt
s9hM66d6Mb+IlnVnmhqc+frj8s4Mg1F1mKf+J9o9QlY5ZUsJf4RMgwaaxSu/5+P5mJZ9eoHKXW7u
yhG/YYcEykm8i8GxZk7fJFJTzUiqdVExoBTBKDsA8DqGzq1dN4PmgG2fsJjQYZr6/To+yRqtZ/QS
wXL/hk9fA9Svkks/VSQGIVF1mzmSqMOt7TwPHvRYxMSqEnlrKvJW/u5yEIPlZ8V0+3SX4+MPOJYt
7C0aNqkAu5XTgH+Bsc+Y0uSWuGTGM5Jm124KCKFK70HaMg3UTedxHdhkhu9PuJZFF8PDoemjGFzY
Jcg52Tde3vzf/movu5YNSNRkNwTqf50xNEjDX0feZIfPB82fA18u5CPIcnPfdTsqT+Hz0FvN1cjc
u7OLGIBt2+3+qxgw0vBexNLOU+gwX9DAty2HRTxEhikRA1TQV20p/PkWPL5gXK9F4dMFWd+uK3no
Be2a3sF/CVuJP30+qbf1xUjvsm4Z3uKyKTc1PbcNqDaXorSTPaZzB8ki8TGjOJpBxpRdAUKZk3/q
7/a6a7bnKtumZvJaGADLsABQG5vgcuDmjQLrWGjRAC9HzUUWJaNMWIWMl4fRVA3CH/P41S60gwfF
pB0ACtV3VzeF0EcN+EGzepzu4Apwc9jsWqdSPcEBHnQYiq4M+seyapO+A2xQ057FOnFGbwNduEqj
4yuwEB0eJdopJqsfb3NBhNjLKTxzOC4v8icKHQ81ljQJmLqlr2GdNqPEm2P0zOFsf+87W710v742
I3fBfAtlRDorrH7itFVOxv2weXQsOtQ3b5dve21HhK1L0x7EA8A5vMYeROJVqfify3jSCjpSERWi
qwLcUpFB8tuWkOhT7hIbFMqEUTQSTLr/KnV12OiIH4+21elUGVB3XCTKSSmaCeuPURWAeZw+eFAG
mSduhowld4u7+qHOgxSgDzDKmiIwCDRxkRnDhAuzEQ+cR7MhcSovVnZksoiqaKXFCZz80tFYRA+f
INAxFljlJVsO1pUDEPWi9M/vp+g31Ii+arJC/+7xwYpuQozNCc06Qpl0pOqTSt2CZ4S9JNCwuO1j
+GNmfJhLfz9Ob8uvKGVTFeIoXMX1sXMaKTsQ7O/vTIqyIWpSEAVS4Wfy8BFgo5pBWM0bbIrRFh36
W1TTiLeEIL3LXJYDz2+YRfgTKlPikPn0PfG3FnNr12KAD1OoqdsC2wGX9BB0+/6odcXQO426mnK/
C+dOJsFKW2/WtzweGUf9dClOIdqKcJTXSceceU/pd68FlaocTkvzVA9JVwh88mRKNKg/044yCysz
Bm8exEBgupuGynPyOmMyO9kqz4emJaVai8fpl8Qe/yjCRVK53CCs5qab7L78rmOyjYIqDdEltN+8
JRKBOenUThwGutGF0xEkQdu+CiDJ6Ep9rJij+BN1gZwieJ9HQ+N6r+pdhD/mnwIRWe0dLv4zdBS9
RwXviYhOlJOy7XuSpUVy0SAyiEIfZ1CglfDbKqLP9/UPlsKpF0niZT4/u8T9jrdGQ0/txyr4H3Gg
qcZPWMzT0HE8OPz9DHVH0FmblUgjBSq3y/rDsSbB8J1Tzc3MdUAWneLUFZUOOIHOC/3rEN/3dcGH
4BPBWrhcXDe7vyhSS0+zMxYeOTWmcj6FDPVKotei/4r2joVJsF3vMuQ7GecMOxZPn09lzJtl5uM1
2pRd+l9edxaibVDKbfB3bnCbX38/ic65qcfXsXnVdCyjdUHrKgz86o1/3UIAAhiVhkGPNfl8dSCv
TbvibtqAIUbQXp5Se0TQ7ieaQZq9fkzajhoNhHJ5hvlkVOuPmBDZ/fxLgBMO6wIKcd2LlXdT+mYO
URZUqgzNGb3wmG+Dze2KCoze1EsDcIrEZVQnW55K1ZuJPNoUhMTabFjEwzjAY7tDvdyc0i6S4jad
Y3zhY/2k3keYa3wPCnoAcm2GDADO08H805zoSjiJOCbcbsqbH/zLAcQbxjRccY4q62/tcK+9q7+b
cpv6lNGPDTfrB64xLGPUvucT635FMSpKLzBFhbdGc84k4GDEpaHylJrJlTSbAHfuLllNxL6lQtsN
04pYGLYlg1LZ90eE/KGh1OMMCwsEPQivq1ymsvv5p8+Sb7k7heCz6moOsHpqSOGzWAjO5ioKWk4P
Iphy3Lvpt+2Cyp62vHU0yB3gfCd9dIJQu9IFZjVDrW4xbPw1HceYg6gvSOHl7FRqCaYaYkIfOpF1
jV/wrkCpEkQTIwsCSQZZPE77O5wamZExobLhKmN8xjK9V6e3dAs68UCC45wCnDc9quKAE8jICJRA
SSASxT6QwdzMMVjdghRucLcdkRTsepxyy4ydokgPqOQZAxf4EOGZl29hwk5IkE9LsTQsxtOftVdA
3cFwazUPBmZZkN81l+iC6ljb/UKoSDBHgWztz0Lriu9fwwBpgCXfGBN+TFpBgWAwHl3n8jWFLZx7
X3AhoKsWvhLVV7F2Ss7fvWmqBKlg3420l9Rh7E6Cwgn2oNh7UX9kKvBWKQnxxQOn8uxwTaThvZJ8
HJZG1mk8OKoyK0akNuZTPfXh0mJHrXXNTtMCYWaV8UYM5P4QB2FlQw1dSvqCBQPM6s+r9AvlQEzO
8B2uudvDYzGxa37MRVhNJWK9pCRXAorfD0rPkL11BLzSf2L+qIiyHk1S9oSECtlp/HJyxWBnjsZC
qQKz/IgrbH93b5v5h3w0Wc0qtf27vuIIr4cCqyYG1WmUPP96Ap6MuA1nr3oU4gaFWY/JN5vaZXSF
aA0wYEcBizEmhJoPusvHtwfBm6S2orr4Ffl0OqAD0oGwkD1yd9aRpMNLlvOyTwNjx3IcjVSEvMa0
mh5jNpDEPdJ8Xwmqu2NSRol69FOt+p+J71zzmUN3da7Zypbr8ygtkuLwPy/sX0vWN0Eo0btn5LIy
7xpiubPu/F+Xu+j9q3wriEYAflMs6d1Qz7q0dvUCCZG7cSVAWd+4J2E0BSkSO+5fN7dOBn576xcF
7MKsxwG7JqvJbGkNi3/5QE623NBVNQJQIclsDyYyze86Y2hRcadCaO0zsIb5Wil648ducGk/Rq++
PcBzQ0ABMWJnntiIwH5xy4jeNvyg3jDM18eeI5xL1H8tIVUZn/gHZ3CJqBZ6+NuAv2cF04PA5B/6
gjBmnEPCdVYCuyMCEWSyov3XeMSRyuE6M/2ryHzpoMFEhC1iZyya+NOYQBMjQhrfZQ9/+AeYqGoV
+Ted3ojpBqpLso7w83YccwzaL4IyfPzM+bze+DNt+hrjx/w4Yl39TrEUVcOvADAsgcvUZsQXkcE7
GBFmsnkYkQS2SSKMxXkdu0ykN8N5vq6k7rfFDwTJ5JeYgf/85o1R4YvB80v/C6YjGfrc2xSmKpBj
AdNKVafgBsEuZc3PqJx4C5Ygcjfs5ujQLBmpDy12rHXa5p0jlG/+UYOKpnaG4kmsg4mC0hYSHjRH
yQiN+0yGACOLTI7J7gBmpa3Q7SZOwzZ0T/nFpxh2XylguEkCCV5+uJfxnOzp/XTUBnDy4LhazjVH
ZWnzXIhxM0tJHJBrLzTMWp+PhP9/EpW70EHrZBpBbn4juAXc7ByMsqm6AMNCapUawkaBaDB59zUG
Bre9fMp76s0n3x/MwASV5U+LZUk1umbgGQBHHLcEkpZ5zt8PzVZAAK+yfhtHMioTkwOWHBVNiB5w
ohCrgZhTOYQG+FtUI4bSh1EF+C1Mnw0CVIZUbZqnE2CIZCXGvBqDAJ7QcQW33NuHgKo7IFaFpRta
gP19wl9rhcIuqnxG+BfR4YxAwyy78ICT92OxGGTjNtQ8DfMNEvUnxFDMUAi8C/TF47TpqL4Zl6MC
maapSWj2JT6sz5BiYX/qTBUF2yURTD8HFVqvNVBxUQkC+GWYKx3yyNi79OsRfuz93T64r3yKv0Pj
dt+Eq6/nKyQRzvGd5C05AR32pEPipohoU2NMqx/SFKS6UziK0QIKARNkiohtNhqAG/qd2aZ3K2B1
i+5agVTyr/MUaXTSxZ1cITLcZ62ad1EKbce3pJfK87Y8wiH4pp9lopk5EE07riXnqmH3yvYcri9u
EN/xx71nTRpZ70OrmAB+SsKQxH/Q819RMWL3yxLpJ01id2m0cULwik9ziSFxuMOZhV5xW/xWXFBI
Tq5cUQZHdR4xnGlU2jnFIh2+G93PWE+GqAaHsF80B04JLXk5vR+bC2ysxncMeotz3DmjvMmx/SZJ
7Oc8sPVynAgN102EIOpTZYgFe30i4v2BFR4H70XAzxCOZkjBjUem8LTf6I+jqvMW8lAdB1V5jiK9
MKvKkz56tShXpAjh3rqvjNDgsFUtQE9FAIvy6Kh+87FmT+Io/LOOj4W4idh5UxnoaUhBi6AZZHjJ
bQf8Hbx/I9iC3TSJUyaTcOCUbcKK7pipkZdDYGd4tDG68LnWEl2ga9zomNPMCMklaQpkWn6eNGJY
z7gR3dLQi4nKd92/UtZvheZYv8hOgSZ9Rtt/GGnc0t6FA3WuE/BAYKtohXGWfTG+TmULZy5Wav2l
8Xd/byjpyzHqcz/+uEce703DAPpGHgrw+o/kT+spT88fOJyWYCp4iAZwNxHo4gBZsfX69NQAz3tP
+9sUIBHyBsa9yEfgC7uHD24HuNJPubiXYw2xcdmJvDMY1QgTAhKFTa3PgpAMSzGigpCYP97lU6K0
1fCEaLd6dBP+SrRx01jit30/47NRwzHsTxQYQspFes4j+gLcTwMS8WSlmUW5N999JQigIgdVlWNT
HjW+bvHQCjvHYF8O0fEPRw9EkNh85zmaXvwucXxmt3xhlmfHNfHXSTz08TtGSlgRoW2a584ac71v
SNzcd4QN8vGeDEzumLxnolrmxN65YVm6CTJj5iYsF2gXST3wwwV+2M5BSIbGwUKouU89mqaWJWAT
kkB07tlvg3c6urjao1S21BI/+DS3fYJPBxBMXPBR/gpO1oIbvUYc01lYcmns/9wIwWr3uCBOAjw9
eI+lFtT2wTuM0pWZkZ+svcY6BpLipaVgmKjgnC2EH67EaKHK3BFLWcOaC0rrv9pkz78prH2BbiCz
9BHn+iq9y54AHQB1JSqkr1zpT+TVkeFrLqqxtRr/j/INwUPWFEq4Ox3bj79BlW1uQvoaZixi+ysf
YQCCu4XZPQXtIeEOayrq/fOc/OBN355hnBnZDEQerbnxacS07BMjlCv0YWHqmiZpBQ2EO5qWs42Q
OMczcOfdn1bXB0LGzlhZmX+pjqoSMK+c+hJGbJtM026NrOcQiHBhkv14A2buO3qJarc3SR5Y+PsW
d/+g5MDIJTeWCOaX6HM34u+FkOXpC100EH7NR3oFNXZwxuFK3ih2dpbbS4ZiiMWvmqAeZ/KZkknp
g1eWbe4Fj+KNE605TytV8PgJbc/1kYXdj8+L7dKvZs6hqBSWpKVCpQOvaLF5LRZBQm5yMOaNcLU7
7D6eRh36a7NgqsN3UUOXWCcIgU+ZsCwkMz1d4XKJ3bmwobaSuX+Acy7CDL4p54mPow3R5HF8Qwvf
/iuCMQs/4KifybYuxaMnVcpmhNKlh2jfwJpcB80TPxQL2J6bZKS1ZVPPXMUN6EVg6FwyCgKlQoD4
d00rzVzHGmnOLLLR2Y3kvEEiQwAHKLaurzQriuCdhF5Ow2kzDqBo8vnVRZV1gx1whpBXjXAE07xQ
9qpU7H81BkV6Cvin2wHiFHpBmTSiWQRgzWWMxLrtzDlm8IsQrLYlTEzvaTC3j41hzgC5ZzdI89Nl
n0GZHSXxQFD6RyzlUr13YYprujROu+AlUx/l89SIuFRjV+jZYNCZB+Wi92BbxOLS9wPuFBnU7/po
BdXVwFIR7JaIfvELAT+tb6QIZtG89jhJPVUtV/Akzkn8EvnXyAl6TTMx78IxkFPNSIUmgIU8mRsD
T/qe3LRaWlzAffxhCGaCHXPDP0ao8W9qHKc6aDKxFUCEKV9/W1bfSck68DVLLWF07jm9mNf16Rbt
E3IQcyAAwxbP3k8WC3u1jsuMDAhFwin+AvO8DJYYrXVX77vKE8+Nob1YnzYqkg8OqrfAcppQ+nga
Lii/eranM0XQ/rS6irYepMzAfqiJ4Liwj7ete6PbZoKWQmXy6PEd7/ZUJkrunQAD18SX0ZI1cSqm
ugfluZ7pJTnEhL6yxortZjZ38kwzfHDc9RE88pl58P8Kq7LnicL3rKd3VfUkKYWHtNBWUVR1GwPW
LiCO/DQdiaXXWD65Qu6RoyiaJtXaHEGPsoecw3ZXr47XTLZVSRhnIt7FYmaGF5MiQk53wwUIcS0C
rqe5AasYniMk+DNATt63hHbPnUHCfhJS4Rb9EDcvy1TxChpoAKTY53vDdFPMGIVF+H3ePr/+pzxz
nrwPtD2/z29HrC2EIGSI0QYU2C3twhUozUWthG9pzMwn+1b3i9qGAvy5c4CTH81lPXX99OIbsGd3
odsi8ZSd7bttKFY9Y7Of24az+ih1kYwdSmDZGyMlRvoYvWfoFwhsE78lKfTfCPJkmnk+U97SMl8m
0+dukswbEIZQv6gY4qpJJcvJoUFQW0R2xKJtLDX7LS9lUfIxAqKnlxVuGbGJjaR+hJGjhgYKnkqA
JKXoBSOkoUidg83piIrtCEifzJ8T8i9yngoV9On3DA0GS27idLtgncxXMhdMrnFYyHDaoIM4goA5
wXJXw5ohCvHvjcZ4WfNjNzAFjIuTUkmAMEh5Do+lXKaXeeSlIFMqPDVU0eetifRgp3KRLTt7O82F
FaEKF/oue7cBmCXjJpf/ImQUIHCqIRAYYsRfLTcRv+zZxtdTbQo7PZjYoZLsR605i2BWIPTbSv3f
uXu1fjlEfPChaKhtQJKE5bz20fqccD9zFRPvUvb7O4u7Ybm9EzaQEmCtAbCIcgN4paVpRAPPBA/X
2LoqoiS5OgVV6d2Hn7tSPv+Bx//TgvNqziuvgwyGkslq0uny+zUqt8YYhfIoPU9eNYa7tV4U6o6z
Sz0h3oYn746NgudkVtbhFIjXQUDGmjwYFoaCoS3g5NxieKzZuZdw20QRoynWMof6YhIsLUlBnALF
uQR7ydZi6Z5y9UowRg4olv1tS0YEE+2kVmszDxGHn1Xe3e4H3RYc472rA41bfD1qRiEWTVMJDpC+
JgEAX9WHXT7mSqAc7XkgNQd2Kc/9NsGD4TFC40E8hvH7ApHjPWlNbiWHR5mn4fCBjyATZaJo2/38
UctB3me3m2FChveGPOkHwdplHzDt7VUH6vA+51cK+Mteq1WZNKoqCJH8W0ARihbzuJaD7G5AgJQw
0z9/LT+fKw5R6irNK3ZR1a+aEhpb1Dcub7V7AbY0DAG/igkQ1CU6HzjzjVpTFYMjxoDJwpd2fHbV
UROeCA1EFzvy2BxmJRhc7r5nGAe5mYIhL8CgNjE/DRYk65njgKKjo4pHUasx3KIGjKCrLm3J4gWx
awNWVU9RExcs34oZap9ObDvaYSBdHsRqh1HtHYzhRbB1Pf6WNxFKmfL0jNAF3OT9OhI/+dL/iOuc
4CoPO/vHD9jqLP82mkPVml8Hljuz3vPz8dL+L5vzhwaj6bmPvU5JMGYyQhRuz+O1MPijn/4vZ88Q
ai066iS/JrQ95NIUWL0n4iKmeziOdM3EdaK9s0tZobmUtnnbMUswd74e6l1Qu5McOhEeIvPegJFf
sWY3CmgK84g7BT87VIJSBC8jTgtBRpjAIJKwGsteuVTY4+iz/ljitjHH2+7Pyap7HTvAyGdDibnN
IZLvJWX7O9x4L/7FpiU+7m3gY8Q8UH97HSnT6iItrDf7Qnl0fN6K1rDHfCrErMF6eKHRug3nRuQ0
KT8MaWTjElzMuBAbzYeqZM/LU7k0sgPAvYt/WSrMqGWy1hWe9mPQ3R8tgulL1yvLwrbM3BxaEr0M
I2uMVz1iZBexzJphNtxPIDszL3AwHIZ2JH285Y1+LDl77m85tIgT91mOC0DfsU2lKLcTeHZkHB9S
lFwYs+BL6Uf0BPFp/9IYZ80pni1BXBZODHGjN33NoX0f20aZCFXSoa1CmldBjyHv4WRC4r0Ohnls
McGyomyD0bMAh+Yi6ZTaBRQ9MTS4eIyLrhTi9a6QQPQVlVQxS7NJLxPrRsZDEpUaJz32jBWmOWJs
KOLAj/AtVkMEdCJgU8h7x0GPhO9zEzS9fc9uhVjg3QVUbvyoKMxM0NTC23O1SyY/kJ2BVuzYQ14g
78APF7cswWHz5MYef9UGlrmB3yXEC+14IeOEwzSIJO9vJHVmal0oxZQ35T63CHvPPPxH/BJbemwM
e6IsBmMcf1cWJuctQ3ns5MaUc1OSlY3rOvybUzeResSOG12Kig5CZqPWx9EdYUtD2u+EmwvMGhsC
5FFzmmYDopJxfasIfTgfIeTWKt/lOi2gvrP+LOKXQV1WbZlTqR6NUceNN+513avt8z/UiHw7defX
xEFJgaLDlBEWjsvsSMU8J26KC5bUr+v8BaLIeYgu2j6IudfV6gFnop5aHzc5aIfBeBJjiXgJd4Uq
jc/u8IIOcXUEvssWdSJQMQYHbJ4z4Q1rpgkjZqKYFHCCe76jpzhqu2tiKxPGy+q27c2EXC8waMlP
ugP3hgW2KwITE6O3M6Z57dGkVryX7tNKBsum0kY/T/TKU6r9Bb9IAcsbsYClcnh6fIhL2HQWY+u5
kYgeEZ1JwCldJaEiCFqN3Wm7RmlQ9j2oIbDyTen9NIBYxe0XHs40NAbT7fH0wcxCwzu7jGkBb3t9
SKQxt3Fq4C4Pihzoi4gQ6MpsKk5lyv0Ho7/zk9CtVY4aXwWg0RyOMZLfNay8zAU4oGl4NIUwh0Z+
P9GcdoVRA2k91L6Zuf5cmv/V5bGMHfYPSd1aWdrY3+4uSdkLiGpWLGniWZ8+/x13vsuuwhmYymBy
BPOpjX0ggVaDEgGVztIQnioa2w3P2HRfTYkQIUfurRsRiyPD4qeRlENUX4HqFP+1LvgzKaSrBdQZ
03UfwPTA2ZpjCb4TuFLN03xQQvtu0q/xT5+0zOO43M2U3epmCcpfY5Hkulw+xzx5y50KiZw4qLHg
I1cNcxO8YBpUx2B1r1cm/THnILselkfXE+hnv678XodLI6CQY6a+b4w8KitZ7vHKdWxBh1nNZaxN
WNAjn8ddSyD68r3IKnTC+8Zmgqj+P6HaTJxJQrbRF9/eZAm/5PpaDhlqI+c4V40iX+9EmjVp1VoT
ABMg5HoaLFmiqX2xo/S00p3TQAWp6qeGMpo5eISTBdPeGT8DaFORfne4dljPIdSD0CaOCYZABdWp
8dHXx3LOguQAXUA+q9Se8q3+Kixtohsyilg9+JRKzgJjCeo7NBEgByOpeFiIFCiv/KttID6P/zl2
4cIZAkw8agFJQbmhqqctExskQQwc3vVqUoMSHNRBUCrM329wHveGSjYtWHZWaD0hDxHiqcSXLSRx
wlMXk2exrIl6r1Id3XoC4kyTHGui1RvDL0JerhKli+y27YfjmVEMk+xHvjbLZJZFi39+YboZWbYp
xfxwL8C8oXKm3L4t1Iblm/TD2UNmeIQzNwyIop9JTNwMK7gqQSxPhweRiHYAmOXNe+TtGFd+9FDf
fQ5ZHK4z8tzVcCYN+r2WSsRLE8WtBtQpnZAXC/35AvbZdrqD56re3VqjmgAa5xGE/52jNICs6XTz
znu77/b5NdMrNkQCM61lM8JOtnu/ImFdQCJzUxq5UNv8gvz31V4jJemZKdq2PXwWR2fZV5SUh0UH
XtsRB/k5FCluj8rUTBpi9ZTbIbxQLmA+Em5kl95HKcd7HFD9eeXitWzCt58kNuMammvxl+jhgrxk
t+VnCPWDQdr0OV4xfzzMqBBBh8VY4j/PlBo6hwkBm0Ew8Ef3jIaJxwW7GfXqzALg4nYf6rrAXQOA
ShmprKV1D/hLwg9DdWYnIpv3djDndCVkjsV7A1S2qzcAAJJPOjF/zSyK0sfQmt3Wv2xlPcCDqw9L
QdkCyMef6sXXUxmWdhZkfdr8zHC3IftY1uKH0dVU5nXWBaeDUtjJ7PyuAGun2fcnLDP/iCdrmLsm
utLEmS8l75Br1NUofL1ss2kghKE7HfKUvOdRk0hzYETLARThjQv7yaqCFBo2B3MzcwpM+Jdl9brp
CuXRLIJrDd15M4EPim0mGhhj6l91MvTlpJHHUzo2/8k2oTsYrB0yKhqStmcAcA9w+kQXxN3n/HGk
isykOhrw4ES6vblA+G8Jklf8ZrvtlhTrStrlSLHMXyz/T7w5osNqWN0qoJg9Muix2vIwktDsBOmQ
GLEb2w+k7Gj/ffuTaMHVGe6uE4hofJSOItqDTMU9VuovnrS6kB47/b/YUN4gIQ1cKxCXDwC5AeSI
oh0V+Kdpmf9Zgf8KJAP1clBgosVLDinhYFVlPkQyz4/j3YLGcK2qWlvW7h5eMKbZl+GHps1aNWhC
vunW0nNQaL32IpCjt9uqvBEEg+pR5AWJn6M0Vao9QNack6T1nuwApLkqWMexcWxLsBk7edCMcDRp
x6rjtEVrNTPBkGoKg3jY5F021UPLUOmiYPN4L1YYdIY+aFKec+r4r9NUD02tcz/Ct1z0lGgW3zga
m3t3vvOUciI5H/ayK9uo4NY3GvH6JJPzPaF5AHF1qDDhbqPPJzh+B3xGoggQtCgqHZlPGwOKUput
fFOxGQMiMSLHlmeF2yJF+TkSXxQO8p8WF7C3lk7KnyJCuEXWjJIBLD0psGBLvyh8XZ5gFZFGa1Rp
9D9t5AkgbnDtqeTfVOgWI1Rme+jO1PRp7SaOql7avG4P2UcGjEFGcCWjoTla456PZqzVONu+OPLQ
zCfhrI6JvsrBuWSivP/2q2OFqKDqpnHURiA/g1qtd6NCGBJo0VNORqzvxoM5NRNzyxSY4kz6JxP7
Delzrs08WSQaYcOTnNs1tKX37vqMFpOWwEfKS4rSJ5V4ftg3II3ajCk8gfC6/QvOgTl5VEILl2nB
WS253PClxJzmfqgzqWOgB+iXQPnipPH5NPU7ofhx2e4mwWRlW9QonAFmqwv6414ftp7ffm1pWG7v
wZifuT5iC+X/X/68ZHV3RBltxVWasOg+t13SVmhKazsUi2Pn/raggFVaWh/GQlhutNy1K5uIcFeI
76p9Ngp6jUAmK7eN52wW0KGn6eMMeAifqWk59YIIzXGCnU0HIc4qmAycg+RrXW4MwZfdGgZ3QxLl
1Aqwcb4z/sdiKzmJFVEknJAn61IQpyrvxoT0hHl0QJPEkgsjpRlnwYaO7na2miubxi2UgKA74H6Q
ycRilEABQUkM7BLPbiEh3PSEaG5+zNNphLp21YPvIj4qZVQd1rJJrWgewl5KoyGUCSjXQwGRQGbE
yUckmSpBaR+U8SPPZEewPAH0Zgd0BqT1RldK45uBqmQyne0+oo0XvHOgPS7oPEGZDWnfwiOSrflP
59493JYCBbXWiUIZtkO2DIf2lps7na2+B8ifJR9VdPQZt8v/LoLyhj/hanws1FWY0wMvjPXnYKBz
lg1jFBiL+H8Y5xzSNmzZG4mICGbzg9sAFveH5lrdmBBfP2fpIAjEtDLvw13iDN1RZWhsexSgEsyB
c+eTv1f6xSxjcwbo8Rr7Wz5LqHutHeMqdZf88AXq4iSPuD050mc54LpId7pCXSV77NPL9eeElyRy
nRDji2VjKjHI8xdrXud8QEuUF3IDonyT+yu13y07suC8oGxE/mazWwkNlozmZqdsxDqcDqtZvD1h
voPb13QS2fsqPT9Mx5bmy1o+QNhSsrTwC3jE7ICfW+xt7uvoD1ZdBxstbWRFDHzZip6D6BTwRhHg
h1O0w+udDBPpFtVS3VL/QMStXMBCPWeAvQ+q1ahJi5FPOUxfvh2bbhqkh47VlY9J/BkJTeP0CgAh
axI8CzD4zhjdp/5tGrK7X2FgWe5BD0vxxPs4MgCflGlFyonhZFlydL09jis/aAMFVHQqaUQysnE3
WuXuBP6b6NadJ9yQhso9NqEiN5LBBEgLF4cq3gRiQO4CMmFPxqbGLUGzEZozY+pf7zzeDgK1SCUW
nCYGWnAKzNn/qxEeBtta8MLaTYxrxMYsUl4Gw5Ah7uCNOlqxcKQ7f/KtQaQRbPDhwDOGiF6BH0Ge
QfUQzIKrbgR//ndwgQ9yjCxvCn7BXUCuCxgrZZ0EXrYbnZJynnrhEo2DKKeFqPW//TVGzIiAlBLw
SEid+yT59IAMmT0GNJLwU4Syyk1sOthpOxFQYkbNAahDAwld+xh9/Dy3sCW2sOsJW4HFG6FNMUlc
f5scXVi9NYifGm9kFxNNf0g+i8ZC7hQF02wwkp6ZMPibtiqIeVOMuobIGCcp3r8cJiIbsA7r7YBz
IkHcwH8NB7mLOmkXwllNOf68QcElinsjPyE0Ta7HKkoyZ5PU921SGkjRDlKtdgjs+SdUAqOvSa7n
ESZSfUne5y5qXbLbaBCqw8aowTHNbzaip9kz338+0Wtq2XDZaNKfIjl+DESwjkA4kiz03UQW6r2p
uQTMeoOWrBz9DJD1K8N1PN6N67PCJvBYFZNJTuI21/uZAm+ABwHhGDp5Y/gKaxQ11XsCkx5dUTEV
Vg+U2+l2w4TsiR2Oqq9MDf6o05alf2Injfq8JYawEaK2gDyqLu2LQt0OkBq9owbw7cfMaepOVp2n
3Gzf5bZ2aB8QbHe6tuoIJVT5ELbewDjsAqqB8+RBqzDuRReyTxTNK4nYi6gR2ezikbhxyJfeH/ir
g8CI7eaZjoRl+049PmwLPARoPmCpBe+r09EldzwblqAAGKv5pBrK3fOCOSDl1bj6zLcefn76ZbBU
h3cMXllMxe3oVppG/zygMf9nq6l4LbvrCz4nnTJDEGs261d6U6mvZwEKlcTeBpYe2foUGOBRndKR
qlKi32iJXudUYrALss3PPnmQr81Ibf0Pj9eFwOtb8/HUVc9z4Tpr5kQgY+Q6+u8RaS58yQZQM0zl
6OO/6jF9XARz4gaSnIM1LbF6AJgO4Z8fnhKozsUFd4LSh/Chs3iep75Gttutx03r+Mdo9Qoe5tMN
jqxlupLkMf81izWmBhbFLK5vNtMO2VQrDnKvsJGJbIXavlpDhLjSY3DKdS5+lRWFKrobXd6DoFnL
h3eh3MY37zDhnaIlRg1iztas3WkO1A0rEoyKrixDkM7OuPIVXJHfXMuLBWUDCtvbWsv9mILcOR4E
meRfsxbXccrXa/eJl4Dg/xaPjKXAFbseKJIwki/dxu63UR+PdA1tKlwbiKD+aSsSFnXjjlCi06US
tIWaJ7SZw07t6cWfssfFvuTK31OBA6X5Vc6GNXDRUjtWqqNJtubnU67RCiccjdiPGHPVHY5ScEjM
Ig7aulYvmr1b+Ib+i91TsI/XjvT4FgynooIZfJezjk6S847ASgyyL12F4rgb9Jnm9dyF+kDw8sDr
K0gsSBiVPCudq82kl7Dn/VkzFSRBpdACvSdZrbmEFhB/F5BQtYle8CNBr3ijX7obWACgY/MUKhQM
P/xejUVTn+WeoOFTJ/M032L8aIDwJl9R80lrcEn19Dm3EebqHtBHLh9fF4wWaa62f+D/fduWTOve
00E2LjCNMqKdv4N3SEkgIDf4/abfBxEvYMGSndDsdmLOkHJ0hlWeBnbZLirHxRUPZvUgBz1oDqj3
6sd2Ne+RFpcw18b9W7D0ujc0i2eNz+AhOiA+9GWu2Yc2IwRhlEHE/gh9eaU3pGaRO6BNaPoE03RS
o+ClYMvKuQ6b0M72VEpB5wR+s+17cyxL0Qb0cTw1bUkqD0Hto9YixhYClVwNzbofEA+8ZURo2kxu
yzOo8qQaMBDvo5kW/l5Tad0fJ4vC9H2A+doWjF8yU9U4C3PgSVIPfe0Eg9eAOm5TwXJE4Awum6WM
1ZKLH55YjyjXPtTabqQaLOCLtl2rHdQDa0vy/Fo6rOsHGv5pQo+JNDf0hmT1LSPXy4xzqMd2/LnY
tytbjcy+czXZBRKLQLbp/gRC0aUif8Fvo+zjLd+RSUrstGHuSGSgZFmXUvYrP5H0iEsN2X0hNPqv
B+p1HOzsswL60Ycuzdn+feEGt5ejwru26Lzm2OXP+PlPmuCfXoEHJvqu977SoPhvTcO5cUNcgNOo
vf57wWT9PP422eajhXKTO+n5xwvVK/5qtRIpXixyB09T5VbVTiLzeUS2sweH/8hBk6o+KAg1RztN
Pqb/HrBDpl20axkQYJhqxux5r0wvyRkqHuQQKOP+StVZ3j1H0FW1blPLTF07tZSJypysd5Tja0Z8
BRlOlwDDrEbWwjJbz+eqCY62CMIcmjQ2VlGYJvvYGkBnY1QqHQin5b5iFR7uMZFRAWyE4NKv4CmD
K6U7S0DziyFQpS+wFzJCPhwZkg1k7BSX+Rco4+QbD1ouG9J9E4qRQej5QTJ5NGMvU4JwJlmXj2yn
1nbI0OILioC5AzVYyqsKVanF9cYXv2QcoE9H0fK7vk1euBAIeN8J4t4zBvwSvaIJtkFBNRwnkStU
kE1qGRzl7xmbv7gggl6WUje5/tgCyFvqs5MSIQpPsJZFJk2Jot63/CIxoNj2ms8IJGtqypkj83C4
kfb1WiH2SpPq1wG295MdcmymBO6ztbJigGpLy9mwBtuh/FqwbD25iYsy7O9jQVTNiHIbpifoCrfW
I9NBedfIwW6coRE/Vl9JKzJLx+Ak/3XG0lAPD6S60ojiYC3JSPxmp6qE76sAlCUAR34iE7ZCJHEt
i+Kb/5Y3pHAxLLRHLgXn5oYmAVCHrLj8Yvl0LJ8lQx2jCoojxgdlTp+QzxOf8hq2d4SmEmq3khbM
8yrw5nwYMw+jWKWGKu7PxGhZ//Aa5Vgj/N9AsjM30PY+sJgb0HUpV6bdJjJNeEHVgiBXUoAOcDyN
Crfndl0BCZVIqqbIM1hNBP4SzPcbKXB0lYdzkdH3KPkQZhnUYKzIypuw5nVC2sGa5+TRDAH1g827
tAWh+p3IaLRnh11/N/zWSmosNN1HkSd+FkdlepIybyNc5U2TW1bgSruUw9Vuady/HjkxW7KhTm3e
k4jeBER/58HumsSOJz6imSAwrErd7Kcru8qB/rbZpzrVvOIMpGinb4MFdk7w59//HbrdUUBviTJ+
K1XNddH+kxXIDmQGx8AYerFwgmNlXRjseWkOfS+F/6948+eqh58oCzof7Qt8C99G4Qkt1RNDJAqj
Ix2Kn7Cn7yqzI0nFW4xaQ9oS+79cN24Ua5gj/jFxNhhpxAN0wR1FWX+EL0KSvjLnSLE+qKQ2ayva
uKqo8+ZfM3t7hjEPH8pCzzE05d+7LIbcqYkfrWX8pOqVO2Vn4tYrA24+mEcQfygvkbLEdrf21YKy
vXyiNndfam0NevUMRu3XfxYgsUmO71cE1Vbh87pcZMQvjjsHUcRyX07r3hZt0PKK8zeienlbqqAY
2P56r9U+I2yYsTItdTDWXiPjfw7nPzmZmGxpJKUlG9W9yonyNP5dXzP3YQQXSbgpThIWuoxC6/LL
rJYMov0g/fwmuoehMdhYaP/hGO2VrfasQOBPvY9PPbmn7zOKqPQSiz9xHaUsiBCstF/ySIuzYbHq
tGf5MHGKdNMWiN0y3iuGPCDED1c/75KJl3B8SRqHpfdJZdkTkVBHo3zqXue1yhheoOCpzc5TWfsw
/qX7HrR1Lc5Go2Brjir4GzPuXsVOqAONuomNU1BBjROAwsIWLQ37gMArK+KsSV1DLF88C2lSuP9u
a3JTPDJQUuS/Gb1SqC1X0PKL0nT1kmjhqWkoYhWdkZAcbjDF/iPdiLAblPPG3Si8UNlxLFfjCCuN
LKBqv6+PaKptDqjOfIBquZPJvujIdyH8ddTXXEGX/yUp5cCGrIHWr0vwVbS+F3xuCObcyXuKJDGx
pVEvziMkV/DMPvarOdfcbgyL/qAtrM9TAbf5yJK1eFEtVPS+/lQN+4QiP07wc3ag1/+XfZ15JsjQ
Ev11SBtSMOnK91KYeWBrz8qcKE6M71evokljrfaF1Uj97ShwanXf3EZMusdPYL7xAaY6lIa9oU7H
QX0JbDpijoBKl7IZwmrRkWY6hA20UtbSRnZ0xAjYkbJ7p/I3s3DZ6doi9BVVj4spHAaOvnzot9f+
v3ytru8TzqGBlQkrZPyaXUQ3i0iUYIYER465pW3nhF+iO/RJbsK/jeNQmDsTnuBX37Q6ypBpds9+
nn71lrZl8gtUpLo69Ey99NbIn4CzDHb2/DBOSnT1LAC5p9epbfGViw2IaziNc28n0BF9yzODTsej
nmhTzhkKgBFnqFkco2dRQy9X86uD4+3RKfgrcGxJbVR+W7wvsBPqwEqP/Wfvham1s2UmB3f6qUk0
eeMgAKX6gNJ3O9qUd40egkGhaADhGpgihZAxBw1nTkR0PvK06qgVPaXx0hxXV6k9v22aNL+z7KXn
u5oSzoDVjju5J0UlCtORi+FSeEv8qqoNZQ7fmH5WvWWLPQKMGFlzzZF7Rb8wjEERK7m2Cj5IE5E+
SCTwSVlxt4+UTJ85cQHhZW0jD5wdwusLvOXZP25HlsqiCNV59QlaaLWQwo9cppxy07CSRQbQe4b4
CTjXOdwnPx4WRsvXStRnwSqr9ge5iK+hGP54pUSXmR9EZOjd8HIMcytSbZQTjdcM1bu7XBeuhLhT
MyLwNhJNscQPaXWkOPYdYaAQqid6AMObD4JPHNeIodcleGAlIN6CV5grk6Q12kBwHNpHAr5q2bdJ
29zFFzu2PkvCecMEJ2ufU0PleDOOtGALttDl41zIx4c5FRYAX5yT+4ZGBx4LxQCj1m6hpLXkAxeV
Fv4E4iKmdqImSair7RMJfHFipzcY1LP96wTffI4lRU3OjMnXKsR1/OEYfmZS4ItqJDvfe9Eush2C
pxbGK4nyQ4+s+5ercqeJLLUm8kuJtK19unE3e7juV45+Lslr9zYrXrN5RE2RIpO79qo1K5eKy9OZ
BcWiaauOgTa3Qcycji5Em2zqukbQSHa7s2Jn3edfUrqdg03QuQPyuJvzcayrpEaM4nbuGaiPqUfx
ocFeT74NwXx+w4YE7PdTzoeiiYsMjZM21aVVrLZcoKi/Mdzbk8/2nPHFqf1IA2z+j6qyfIvFQoMA
8oKcQ8T7rWcHIFvL2zD7kU8dPr/TgvfiZdvRrsgUWp8BmlF9DtHz+YPr+hWKoOpIjXoDqYjanA9x
lC67rJb+NcN3XRTtwOJNsAwafJnGt6zrcfdz8XQBEtODGKEgVaHyvBu2o6uXx4BU3N4PN9qb8jU/
d+ViUPiEA8PTcbvnfoSDQbdqKjfWj1ABr3CpLqTwpU8lUMtZlxNiBAgRtktCOFzrBubnKQxS6iKD
O6INeefp8w0rvADnodVdd5V3zKbKtbZ1slPCwJA9+xX21lIcsjaNJiz+z/N+Ug9IphDLsNIRq0oJ
K5jfF0OBJBALGUohnRDTbS+czPjXH/Vihk7ZzHfEhQLLBZPOInH0ds7PgLO9HdiFZwD+ZiOsTe5h
7PVibGipgsRl1pDhS6+KTwNg9aN+ziWZBiAqHTr3LFv84C14tpwtg+nLpNqxOdgsDIK2YL+9y5xc
gcFZxLIwdSdiNdPeyrQwdmsm2ZXriSuWzhPi6hhai1SckqjS/JBNnmVUkOgbwTuFDhXxUPqJxYty
E8eKz5NiXFNuYTqcmMsAvTGdN9crD0c+kb/yHYXS8NnOdurhhgnBm/z+Zi65PNYKSYKZ814mlFRg
kWNpvJbmERhUzCxmzaHazMpEtCBZR3QL4n5f74iv9BpTnB2EeSpMEZwV0A3a+n/B09KhDGy7dyAO
7hJbR8SPKcuvWxq2nSzWzwQifS16Be4kqk1uOQi+abAyoXjD/Nl/Gso9BC7u0zFbsL8rW9hN3eJt
AWbyNlDT4et9ry7Bxe96rOnshSt3PsafgjSHm5Qql34SxTVvAWXszZSDFikBhMNkkdz3k2IvNyyr
yYKTNXVYXHMQMYWzXUr7yd9wQbuBbCVoGGuuH540CsA8UxBa2lOwGveZIH8IZ0j0EFnEplRGXshy
1VrKlwsor2cUYDX635zV6wPcb557tVc+wNhsGt9voHKCvdMSKIDNzbjWgj2WzBM+Ncrki3jUniuC
iFeYrZKboCqfKzd134/4LTqaZSJht6FaEL/JcHZnD4PEyMK2p3t1bubK9WvzHuJp6M2GfPqlqaRM
yG6eN/FKkhW52zryHYSEmqny/ZXRWaQGCv1r1R4Yp2e7xem48GOMYG95JPWkKU1YRO/4VSyiE4+H
imF26SDW1R3pnXJdwgnYVwUnjQU4tTlX6ddIFVJTLBlNpAYKtVfZeAe0aA+f00Ok1Wbv1KZds2Lb
Pi1s9hShH514u07pcqMHoAZHe4hB4XdIkyT4/Z9ZSSAWWSZ6xE2UTKxMbiLTthClLw7c2iT0q/eb
syH0yKqk0igK53uiGONnIln4Ecrdi/TxLg6EFOnLRKizDShVDH9fe6WfYxxn7Snxaiphn1qiqtM4
4RzldHGiEzyi4thxH/mPagHmYNKKqIW1Jpxl9kuyzwlv8GZQDooiVO+dshn+gJTfQ/foF+cGg8zZ
Y5fnRu2gGRdUhXpZs7rUkqZX11jSdW1jz7sYJQLaJWmXW48WwMSL9xXoqrw+qeW7v8CULuJ+bKUP
FVoekBr0+hHKnBMcq4KgXN9eeZEmh9UKVFw2nTKdVGv0hUlQ4Cosu8Ixzjjq2+Jo7rTiCx2USTh/
EAvWKLIJwWr6lf2JkX8gHJBCIvAzcWSECdxE2y/lc51lX+s+2uah2C1pdTkIP+TSFDscyp8CGsvG
oyO063MazWIckEd1+Lcy++XAIuiYDCOm/gbvHgaIcM8Rey0YBjK3UXWWgfpVBqUCbYW9DSVde1b3
xX58+8SRL7QYGoGoakzkLjICD8uawr5c+Im7FfM/G7bnNeZE46gMAlLLycS5aeIyZRah6vzvO16h
6JyroDjDAq2nia49iakBPgeK9Q9IK1lIAZJbgRvJrRBfJDFOeZNjwn3Rcpt9GWzuGsG54qAMhLcd
YcPS6kRWy0xqtxeWPnUekO1vEJ3oxzpDKviYrrAwU+3Z485ffgzVrHgXIZMcXzp70cVpvZBNJYIb
q0JHXGzOBx/M0D1JblF6Pcj4QintsOS7k2ZEPWmJMF1/2NP5nmGydkonikcOwUF8Fm5hfhRNxTp+
YXvycGW6bNwYvZldIP/v9YhI/gTt1Qbqgw4mBbr0MK1n+aTaxHnYp5OukGkoWtdvLrQ3Y7h+4w+u
vuEZeGckcRkvb+GIj3Zjiivxhy3lPKu3eEizFNKdQ2dU/h16Qd30rcxBEcQjDZbsfQVqTP+42LHR
e/pEv5WMbVpL5amnZpsyAZILE9aJPuCzugQZjeWjAhXqUaLmicnybX01F+V6JhOidhv2mOHHJrfy
2pUpgfDgdTXBYEDj+BNE0IdgKoTeeQeZrIsVTPZsMLSlTgjse//1mInLD+kjsisZ7x8kgWuYf6M4
v1ZUPUot3Y6MH3iNjjofscGoTHsC9H9dHO+z8gLmdJcse/26iZfKzzQIfj2Ga9WmDN3P9ydLQBpN
qEr+DlJsaFVZf01OASUL3pK9LOzKw9R6I2N0h4Hd7vl7A/Cz+5pPMgMXQB2eH9yN6x/G4cBeS1Fa
7RZyboOPHNjFx8Fl9lvJ2DtlrJkC+4Y+9YdzHGf0TvVFygzwYVxf2oIpthrwkgc6RMWyNqkziUHI
k2ilIo91VlnC34CCA2zE3eCxxouh+G2ZYy5va1209Ems2zKFCYLpZ0mja+SmKkWH8dIsKQlIzVoN
nLwuxQs7+yxG6y7E7+XmZZLXz2ho7enE9CnXkae988RgQw/ayepNiOJtjjr+z46qAcpytz6OB/zs
xi6ODav1OZJTbSKybl0dYmMZk/l2axPHYS3soWPu9laHwDSBp5ixp6ySM6j1GBnnBlcORvA8OmkT
PoZ3qYoM4IZwtiwplrYAFJHyAPA6TXDgARPbNrywIP0dvILUz6cTE/El3XE385r9VfxgXyNoMKBQ
fKUUzO+ntEAcYOYZNh/b/8+zejAJhy4eamAo0HIBiDpUcTZ408C/uV4jt0o7CxL4qDqNGVPEvT/I
ZKzZ/cEkc46kejPHpHHM0x7Q2N5F3/eChmMQmsqq1VlEyjFo8oIq6mxqdMshjF4HfT/z8pwUwh1i
lOFnJcIGuS9ryzW6DeJWLgzPtBz+GAa23dQXtWZf299k0Xme7zHG6nE5qa5eP+D5dHDul0k27dvE
gIUD4kG3PAVA4gjHd6mzXYjf+7u6rwieuH4JgmiIDkXITHlODz6cxfmNzOxYFfCaXBOfbekPV4TT
7fYxFw87JPKkDg97RozoaNRXSVRIXEcw46Em5a36Y6uWDXWGo+Mo/on/T5MGyAGj964CPIlHK1eY
z5YHw1TtkoqTaLrZVWL2RsMRSSYS7VhVguaBN1PvAl4SG3FPADx50SdwSEWWOWGjffbLci8jEzVn
MmbHyK8LTnzXBjON3LmyrfNyRB49TVlrQ14cBFQainMpquIJNjtH8v8d1zQtEgcZakydZytqBTan
F1Zz7l0yWeKws3T0JM7dqm5g7fxIIwnO0JFIely6h6yuJG6onXiQPOCXF3l+fksPyto9WDMOKymT
EPQA2STo2x/cCYSa3neXyCebALgYcSwCugQP5abm/1tQNfqhRHmM43QLICLxuO4bL9rWSZXrRVwx
Var6fD9BKD77K2TMeKX/1roj6mbroL6ab5TySDN/xve9K0k4E7coCVHyhDk2PSmFk0KP+ERKcVPK
TfXCSkIW+dgOPf1ioOJcDE2zFYG8ALg7gq5yZQUgG4/Wyd5a2qm8h/ks1kBPRjFKXNftsfqhJDqI
VFQHhHTU1+JBQ1hZaAxhtW65jlXakmDPLC17B+7M6d8FlfgK1uT9/nCoa8ScCV9JnNcsyfMDsjN5
X074HswNwaVsITZnkoHYYvx9irZJRpc6WG//IysNdM8b1ZwPcDmCvWvkc6jetJuyzwRbM4fHe+Bw
w5Ctu9MZn6GCjDuo0sio2rDqguAkdH3k+Mqkk6KVTZSDVbzmkncSbcENtmjmTixTDZ/aZmS0yDHd
U1e4dNjdRZaavo+lW7P9lsWTMIIzVKu5mzF3FGn1ygd/so2ZKiMi5CUc9KoCaitZWyXfwASBQRgC
eyBEobNl3Q8YjFTP9RtH3awSDwgewMd0eGm0BLCfufqGoifsQnS9yiUwBs0D0GQfwnKsRqHEWVLT
mqBjUXQfUMeVmjLXT9B8tzP3QSoX4h03Pf3D+NYw1kZWTEPUSIJwkVANDDSE7MRVhMR61Q8JbHR/
2uzt1BJVPY4YuWa5RaZHkTRM2ph491pJd5Od+azTIZYXDgyjYszjdCb7X59fGfzxjsohsi/7ZjGv
nkvEWNWLuXSmJ065rddkKZLOGutQFo3lf5clwWS7oA+7m0VpVzed4V9m/7PaIwM8lF3sHKgvYyVr
uLvvTBAUDBBbZFwt+bf0NmyD4ys2spvzmisIjgM13Ej1Dk9OIDzib18IUVlXlZpB0Rrvqw6bssct
ZcTcGrRQVOAX2c1Lt4MDQefOaaizLGoL28pb4CI+NrtYagoBw1U0IZLwWffIhr4L0JNaQ2hu+SmM
OPqgOwCqnH3chfycOKCIE8OCB23MsQ9XmTl/KWOHk+zcST9B16gW5qK+PIXxS+5hcjFO681QoTFu
yT1aTYDO1NDGQ/KRLvzTN73qfqcm0O7Euj4D5kPKe0Nb8d5zQCctaA3yc1XCTgOi5T0KM8RoNS/J
u7H7UwgTLRbqSSvVvwURsMhr1k7qt/OVbsKpG+tNGLqa2Hua3jd3kF35uzB/Y0hvumTKt8bJAm8E
U/7ee49yGcAEsE6RGnj/Za/XhYVIPTeS4DqDm2o0r5mmjCuohYoC4LdewAGnVHafr3sDSLDjOXbd
iblnQmvm78nlHfliZ2wmuTOztsDM3D63dB+7Eb0zr1I4smOB17wohduGZe/fBEv3dhVwWgw9uG2e
QdW23C/OLox3PydmfJRykxxgCwLtG3Qy63j1vSwa0gmkat8gAh6qxjuy9zPOqTdLYz7n3NCUbYOt
NhGkhxZe8x72pAaORQUWt5OaPEk6Rg7RIeuEMG85yopI6cju/IK5ldX1J0P9zTNujvOa+tZyFtqa
DyObD+I4uMhBrY7EEIyTOqzI9VLh3RQYvROdlgjXerMe4zmYqCI+YmdtRTtZPEImg0awN5U6nIW5
cCBjuQLQ3oBsapDeyMHNcnx3j+psJpo/fT7y+xK7tSrYGBYH7ytqq/7eNTUolm1iHIFc+bkHZFkh
TyCjusTm3YSmvh24iOpuEWAFquRcz052gtB0pf2bFfOCFlejMj0YTkIvTfTwbZM5MCMIETUz0tX2
YLUEGUnDQe94e+j7ttOiTnlPIV2VoFQ2DnPjVvOh7k80r5KGpQ5fQIRo/MmZMB9LTrvRDIu8Nk3v
LRB6qL4YjUhvVFiVfUZVyPCDtJXIJ5lPpvyDQ2BSLylQ/Z8Xc3Uejztamue9Zk9O2DjaL/UU0tLR
nHHDd+63R0uCYcEB2rwrpdrPEPtf2XzPSBnjimDBqJ7tjgr2sRdoN4JcrWe2cYpjAdNAvLNuBKi+
L8FsZzF7MsUpjXh9uMazCgqNaut1TvQOajnkvoV+uW5Kp7qxEzltFJ9i1qKm2f9XPojsOO42qFmT
kijSs/OzwmcWpYNkhXKPWZAiwuD4hT37Xj0pmIZVyqtXFuqi6VUOPrgM1NnybrQYhrpsU/3Tq7QA
0ccbvbocidWhvo1+QYLuvXGuuiE6idlsB+s8Wl7V2cQafXxWMjrMNy45aG4t2lYGnKTguZzLC0Su
Efx2iVa3B5fgaODIgJ1otK51xpliooyvMtTWUEoAnpKFfQYlGaUCPlaKqLHWgoxibbsUB1IPcHae
s4Cn8K5raClG0qwzjiPOQr2RYf6D3HBcBeawAB7WCqmE77uu7s5gbx84duc9WqXAg96qD0GC0Vui
0AfNOH/RggI+QGw/9T/xC0/lhRaJ3ZZKWZV9Pa0YbqzU7BBuSQ2ypmdn2DIjDwsG/Wy7eeLMXEZ4
amo5359TLuRlXGafOTg/OaFoyD7s2OA6dJL6i94aoXV/ts/9edQiJhyJ4A4Prq3XMm7N648U99Tg
U/FBLM0i4FvufJn+1Dt5XZaXPDVRABFxNpiAoK+riMP4A+4xd7rmtbSlrVW/KtDLH4+guaUvA/Mr
20mAHvhhNCAVYf+jqpnrY1HGKbE3BvczH0XDdVJGCUt0rceha1jkgvGAzJuV+pmsJvpzr6Ck9atF
qICjXPWzjDFj0blqu6LjBLFwvluGmqQmSoVkFUNbqdxX3sAISeyJJA5ErZHcwTYiWicNxvqRDpTO
3WHzrnnujgsGGZJx65GFJQhXuVBHmOSdSjD3bOoSjeeh7015WRfCDEDqiMoMQQzGYVYQ1p/71YVc
mSY8otdK2vN0AjE2IeIip8v5yKJEAJyjAQ8xs2X5S/1ookgeIJ/eLXkS+BI3QDPjQof1jk/swJnS
pwIENnCJ4r7NzwXWXAMNgpLvi5P7c+9upBrE5E6kcM/9qlgAFBF4/QHpe3Z0DIkNT6p61hR8MKuO
ZMViDj0WGVlxAa6R6Pdz9bu0EzZHOPIKBak+Sp2WeDlwkuC05/FJ9GLChIWikPOI6PqX3kIcNh4e
pod/lx/BA+sS0a6vlT81Gpkjy8K6tM681epiqimgIqq9YBXh5/MjlwJ3mWJ6Ba7SiP9xn3ak73rc
DWUf5TVm67SqESsedM1KX+JDCSdeGsQxpiL9EuDGMeP2lq6btZ+00GwycF/FEoUCmUTScTftX+Mw
XdA7d3DNrC5+1Dx02XQQrvu7RbK9skGxbPHPjxe6ohakXnQcd+wXYXSPW/4VGsU7wIXBwKV12E8s
9oXWZRnM7ORR7s4lW8Rh624qhd9r8JH7IVPUIq24eSUUza6Wu4xFaAGDSRdq3a0QXqEND8JkuHjW
0JdsZXHQlavMvYDFqxsu9WvmeafvxkRIMhNVRnHsbjy4O0sDNUjpY50Brzorae2Zwagjnrg6wM5l
3CmGrsKzQX7WxTua1Bt7jRRx59n39YzTk/FHXD7klma8VIvqm2kBmJeEw79wrSfnZNlS0yFNEaxj
dxgTUKknwWgUBzZjahsvkT+hbtsVp+7uN0ci2dkb36fpEvWoofflnn1hbFiqTZJYIeM9nywIERN2
GBLjhBal9N3ExECoyiQgyBB5ExKr69fFtiJ26w9wB9TXBcxrh44RUWBIUW97F1KdgJ4wAGXHzfYS
IW9DSj4QFLjE65xQqLCnwTocNcCdXi6V/sJ8Q63DcDBuA15NhU6J2DFaWsACFoW6lAmmBbnDtW3j
S5rLZbyk2kYtmYPauxMOlEJcnByxTs84OT619ARXkpeBtdLSIfgDIazWpFqDuJ3yFg3BprB1zlkf
vv1RQEmhjJDkNauyZcbxDOJbFMGYIbBqbPun6VM493kornm/Z3HObJnrwkA3FrJWlTGaTLT2/bk+
MNhpIbGjLR1iyftEOajubWbmIAm4K5e6R89WpyzUDKt1wOKrWk69esBVieItDPUvTFt1QrM24RSL
tWpOpRzRl5lvpHgG4nIDRWUMsrxdSeAXbiCMRWtVZ8gba6PmjOdCXN4ODKjGHKzJXlXmWLNyVuXb
kmw8klBsv/evnJicpWKzy0h6Bp/1K2yALPfkBS2dRLgm9Gs37J+Tu9JOmdmj3WY3IM3GWIuFgwk2
iliG7ojCuqyjevz0MVauhtJnhL1kZCQxtZmaGWC86I3QT+LrUk0PD/74NE7K8ch1/tzvt3+fEntj
0hxKw0KA0pv3qpStSAx4Hva13QiFN/EapEUa1QBLKDBiqpJgGsdPu6IMdyDwfpznlyIrPuJGbDGK
dWVj3EpHTOiVXNqUkWvcGX1cL69mUk3UsJ99GaiG3PIiZYw55CNoLVBhMmG/PbIf66mxMjDlwpbj
WO9OwsQc6sjKTbT/dg4xD0A0pCAPyX3ZfCe098nwJ5yWTUHf+LRT8aQ71yDJbcu79QcmmyGpOik0
47JAFmPgsWtWjfpGt8g3SeJ63mo3xvhk7t8MQ+3Gg7gjK6ZCuSEB73F7jQfhL8BB+YqnrI3XYFnS
uEI5mlUALS2TOUA9bvgcLIotoMlXxgi1kwCi/J9dJ4JDbi07r9MOy9j5bXTpRVrAvgK3FuaeMfRj
WLatEiW7ZeX5Q4Pmy6TfJMuj/ofCrZ0Y+VjMkJ6G7/zSWQmF/9LG0bgeJml7iYKjBi+5ESXWQ+D5
LHCqIpiF3F1/UpQ9mVgiL63kBNy3b5IWomynUuBsz8RzZvryuS6+oED7pgbbrHpEN2BYHo/pj+uW
1q1s/k02e6qqdvDCHyPfxghKBkC0/i45hPSwwgu6kQoJ7J69KflWb8Iy845nkqwOoRysyP6J4DnW
qRmJ4Z/Iu03XVUOi3ECOZ3wpCGQZMPest3ogdl8Q/O1DL8AA3I7VeCW9adkPpG1Vm0SEWhuAHj72
W27/PDTGfuiTaWjssikMkdrAC1I2FayeMuXr6Q7lN93tujGj/y8GnVJv+Qf6/YgLAx/8WBmeV+a4
uFl2NvaHFu+rGp4fWhucFLkGPFH+pKgf3XDV8Z05FVE1PEmKl7BGbTgruDq06Nm/NKNjnzwVLNie
rx0kV3ahlF2HExXX57a42bvX/ututTVPzq4OLbeEV2vS4m/968E6/QhTQ+aMOY9Rex2z/hb0eZhu
QguT9pT9X0vBpAoIXQeft3xvfMkKXnLAELWGYAwwVFFzLnkjtnGqb/FQr0z90L9JDGYNch5vsCRd
3YJqARNXnhOWKI/xRrFYxQ5BGGProiG3IlbKkv0PlFe8c9b69xV1UkC9TrIldY0cItC4TCHBejsQ
dOvIM20dv/8XyFhaJx3EfVKR2UkaxT6uvEvkVbkVL+PNDYvsiRo+ss2P/BgF6zII2kgdoO/CSCGh
cadO/ZIbVzFX+lwyU5KKmigC4JFKisjMEnyxO4tBgPfxEA5zQLfxWwSf+1h+7N11hzJdxHciYqPY
pCC5nvS6J5aX83xIqh4XaTOHmkoy39HxbKxFjLruiVW22Dp5tx+XT4MRbEfpcEojYgHQxrtaNjA5
/kKY0a9o4pd8XEgco0CJntsRHjXCKgEtlWI/Tieai+DPbP27fjuUNoMtI878/E1HsR2xobiXR+Qo
QITpxrjFkaT457v7HKXXm31dDP7pkYEEF0tG2QI3mgDZnl7k3XLhVI5LizpfqNimXaQ7mkc2Z/7w
ByJ9LkRPjERZg5s+SSNgP2IabMKqyQ+m7Y1n/26vH4TqL8ZkrGoXVFlWub65Z+Zvw+EMOyL9s7Uv
u58b6ibLXf+lFwkPN6TF+MHgNY9qhgj9A5trCPPhyTxJnOYxVfosx3RbG9FDUE7O+mZFaNyNl1HM
YP+kBJEa2LkpIZ1xFfi5/KeEOvukrGLG76TSyt4O3Wohjytke2DyQ8envDzjqy6qrbg5opYE+6lR
KMdLe1il0WehfbetTWelmlzVAnTBa6TjITgvuUumwwEuFVwoGBcbQDoaTmm5C4kcCP8plNQgrHsl
9f+oQsFBN8I+5spFH7nqelQ2usRZHKhWjstaz3V7GGuyShw/Y+jBaFX32XEaiFrPpd/An7CGlJUl
CT/CseWKlcA8HQNjGsC6CY6nCzSjxArZ2bkNu52Bme7xiPyXf7d7nsRG4qg2PVkjINy9Aj6ZwCAN
ddw6Ur7oc3kdn2fiGjL6BkumOwkhU1rCiaG0KwM01Vb9XD66cdbLv3DtPjrAOrlZkFg+4WdpOZGP
HGzfGh7arChHCQUHyl6cj0Lq0AQq78XD8laaYTv5Cyz4dbPDnMxB8zr3gM3U3KuI7vLis0opydTg
GVwLPaQtxG9oLAuN2sXwrn0J4IWzigwc599TVqTvxbmUQDXGMAwM15H+CYA31gpUuQPkHwIffNsp
zXxOEGPWxqDMs728MuagtKSnrSzCe4WeRQF02SVF5UadE3Zo95wsTMLvgsGvKTYvdErVET2tlO5p
YFR/CoI2u9ph721fxNhme1eoc2PTxxC28jjS9hLRL8CmSVIusaiNIR0bSfhdjbzX+nAkH92aWsTK
geEiAdhhkFwQn+GrVNTDFVa6fkzgN21WySfBYvI23Dj2iST+AeR2uvUwqz1zFa/4hzScPoM5XQ+0
+D1yT6eqNz1Dmk3opwK4EmTwtqadAy2QK1fVXvru4rDqA+WkuZD65rcQ8cxWN/86F4dLPqVOdMOt
15Lmk+uZDLOWjnHzGMsGjxn6awXsMYJd1vGy6mZY9UJcakVE4A3WnR4SbTgfMRf7QGrY8QuZ7v/h
WzimtJ+JhPaHojgcGncQszvFoYmFfSy2az3LEXtjjEYYh+0a44B2J96RZhluacWvwNdPTKI7VZto
qAyRX8y0N+huhuf/P2YW1Mh+B0DwV29IWlSP23Y/mJDR0m2WyYx3ylLbs391ltnFW/WH+3a6vGIO
W+1DvqniUEaK7cHJHvHbl+vn5wXJBCcBuDEyEZPZAkXMZtNyKTETNchCGW4UJq1YeyJ3EPIE2U0/
zSZNMq2RXDruLZky5osQLENYYrv3kh3np0CszTOYjHgHCwhkGgiExz0RdoXmjg09FqmnuVvnT4+6
kMlsQ2G87Rb5gvIWHhaRWV8qG/mOa7v5h+gYbmaTduzx9g3/MAgCfQ9c9mbyDOkvHJ1b+zjshzjN
yB3CfKKYWQApd29ZHe9KW2Cdu8KO4WHlatjInzmxe0wWWNShjCbCl2uxyUQzKaT6EiemlBznkJtj
a9HJcacTuSEuZcIiA41Qz3NYh9q/9p5Uk1Jv3Zv4ny0FEMgChnDAlpOroRIcolr/srDy4JH5HCdK
PG33Ez0lVco1ygm73Zu0hiGLMYjm6JVh8ncEwR2IfDkqOHv2W2rmAaZq1fFeJR+KVUf+Ao3EryTx
kB72BW6OPq3ohDkJVMyWsXVST9c3hNixb9zbOHaazmldTYEUdPMjO5SDxrymWgjb1P8hn2PaUH2g
QVKxditG2Ux/NrdzGy+YejNC1izK+PnD7x1XC4q3Tsv+4Aswvr09W5HBP4wpVZ0IJpJMqQWIy1YR
BIGeh89LIsRrev/8teCI9AkX9AAulnDqkR33vvPy3Lho/WuNqHrEVCWMWqmUwXA//QtQGB6oYOI0
EDC08MXXLDY1nqt3bv0vG7WFDx8hbOXuKlB/TFpCxXYhUVwUcr2u3PBo4Me9oBIpw/0/FTYTyrGL
Bd2X1GjsTjwrKH0zDUJSZmC3WcSjiNypeAc/uPyvJv/4K8B07qEGKTd9qC2/Wq/mlvgfM5koubh8
j+pmHub44WJEhVuzatY5H2YFoaH54Qg7DOoh05FDp+4UxxbtosSi0ut0Ggju2sS/5O8OoJHO1Gj7
ml4fpTgdsePcgbjTRBQKG5U6c4jimzUNRn7HSjyLt+r9ZrJkT63TfzHTup1UvYWm5647yzJLZWyy
S+qeBY1rwnFcfkgwm2SDOE3bVV4PaMH0kktLp6zrhFvhnTI7upJUrRP0qD9ncwQsy6uMq+xcQ5VU
2lvLKwYUMCLoN966l44+acEN7BKCBxX7RH6iFtIO1IdD7HRul8jsF0q47sFtgH3FUfGtUEPOt4Q+
qPpMomBmJO800B6d9iaTUAgqmFUJUoPJNutAtHrRZX7qiSW/w2Iiq66lg81XjGbSx83MXvkRkAjf
rCWbHDen/L1GzP+dhO6fFYVp5OfnY2cikH8pZt9e+SrCdJIDnInNOow3EWr8yQL8VdJiDqAS7kn4
ne9Ix/xImxcqC/OqgMtVsTbSzrWYmT0CrHcUy0GiBO1/rjsYzcoIGZvekoO0btNQBHzeyeomnGIX
fYyUT7szagcguJqh6b8dnIqiWereC3ybaWJRo1uL27ExvXxYxHtN7yKoHsZdGWOVHrR2KqhjAB4b
Jy1GvAwcR6D3Rp2bc3BfsIP6foSJxz05V3gU5yqkGtRol+ZZJhU5aDFG8TIiONEkpwxn5/SWlEMh
fkSwozV4WtQ3sRfkIJ+UKOTJxX2ho/wv+Q2opfB4ovMRI738bKTQTLpJYijwB53u1UsZ+0LD+5zx
VDDezmyziTM4fAeIM5pTD/YI6XHYzYhrItAdpoQD7JoZcbJIhyVWbwcTcoRgOyUsWatBIiEiCqVO
IvfdgRcK3ZCHAW1eNgRvNjXKxAJeLN5Oim0G6F46au2Ee/3ZCD3ZAqIqKVJlF38L74QIjK9NvzZx
WG8fpkG2TvNliY6ymsz/mPIVhZl/6+sgk83cElzzXvHdI1eoZqyy4ZxujYdQUHE8rNp4cqij/J4e
/hualMeZzBngqfOYRqilDg/srGwoT6uWDvVjfz90Y6puqzsJLmwUdfD40reAK2WbToDaZR/e1D0z
yx9FCjcigUBcLUNNu+Q2TzpIzSNeVitYraKsBFD8YC1fvcqJVeYOHBxMdEImkZjbwdO4A8VSxSj/
h5cYwMYmYG/U6ErXxyLfboHOKcyofFZhnbGDRnqBTfDiS9ETGdydpqE2AFm2GXLXKX7c4LrnzazK
672DpNZuzwNLSe65jx3iMk+7w5qohGkRwfVNuiUZi2u/t0SaQQF2FhAhyhw6QEIkXiUF7i8vNz/G
BOK3cdmRK+xus53xb3NzMxKlgZy7NahJTBSjROqtZQCNgOVZQy2wwJbS3fik+qH4krsIr3RgLMrn
+pY7D63bcBBjYAk+8/BabUWz5TYOeGSrg7l4RzL/wQYJ7V/bQu7IZ1g5+zCKoK8Ins3QvFA6E4N2
2H9Hm7AHEMuEBz8paZBhkLwlXNs3j78zQikcYhm6wJtvhYQA0r/5tS8JjUnvauSZQfY6qatW2kYV
FUlaVZHGgoU6HRXUzGBobn9CWL+xaAU7tP0aDqC2floHZ/eIlQ0TjGLaTzH7F3PhhPbg0xCawUja
fendRRJDwFpdpaZTykmDa7rfLmpGrCa1OZ/VoDSsaHO3xHELRBmKerMOPFs9L27r7tF6KQJZ+6D/
0tUhXn9NgWJpIoREVmF53nQbX2hVARRn9mtMjRTwXOMt3lJtPUutC4xStC1TXVv879O+3kEVV+wR
slECYoIG9hUrOEu3sU5Saiy1WXNuJxHO3swyirOC7PdpVm2gwQN5PqsbfVIUtE0jPs2BsC1q0KxC
zkA1uaZe/GG9t6vbrQm6yTKXTcvEP4dlFQg8IzTTfS6Oxx5jJk32JqRR5xohxK0OjjeyUxWNkzzS
xogOJFM+FxzZe5O9rjcKxBYLgzSRbCFYGEtyeuelNwQXbGbndCcfjNfx2cc8drfTqatrCsOJZX53
TX5FH66VoHjdZncO+1QsJHYX2IsVrvygFfpRH3wsdtGR/W/6Dz9ZD7VsMwxMqSK4QeKHR8uJVinN
yJWoeSUwSKRFNHDU40RL3ga117ZgNtnStY8D+RlszxTY9qaEqdzgUT6U/3qonqLpSQvKvmxbQz1D
6TrrFHADk7A7eTVQZUISBB/VXaHdMWq/oS1Gz1grJL3rj+qsmIVTHzw4XHZhFPLe+wesWY0PeBHC
aqgiJYYpEGvo/sbXERj6XgBHFuJDnyHCiQ2q4C92U6NecpfNYURgGeT6+xjxSv2V9JzgielAzxUY
i8zbuT8knTqmO4KY/xGyuWQr2oOwEkXyiKlIX3kFjqq8lY+EcpYizB2c1+vZ1VCnh84h1XY4zhQU
N2xgQcVBICmzSvFv7ku4p9W3rBCsvJNmLR1P27VST/QL58bYhg7L127YK/DKdGYnj0cZmrlB5NHE
XUpmRw/vCOiMnEzp4Y5d/8HtLNEJhKFB1a/pg7eNw8wjJTTvXxV3POzdPH7qCVIaE3QSu+SkBd24
jJs3W3JAC1pVxO+c1BqlDAsFYzAzcb+xUkvH2u5SXYiF8JUsPGFbtGWSkZO8yQpoKXdVAe3irSMQ
j0djGh3ZdZW0JCl0wcanJNCO8tY46ZhyxW6SNZHH2mvg3MR3d90MynvcqQ5GuF3hlWM3JvUBSBMI
fDSq/NwRs4ysQ0RG95wVijSP37v+ypNJC6J708GJn/bkPlcDae7tfU/0b2h1KrvbKtjzAS7iQ8t8
F4O/UIv5ATfRAcLVFJKubdVrMFj/KZXon6o3/b7cnmBGOuXTMDaW/GXQ/YJ+e+1xFxwWodloglD/
YhAn6bBnPL7aMVZxB4vwlDjTWg/SBp/MBsIo2tMhI66bPvYcL1uHYq42Q4ttbnmgC14Jyr/gs++8
zYLAFY4oWmQBMg99esnXGjTXV4fAVVoXesxoi3SExFScKm0jQs08TCAfCxVfPbw8ghl/n4fBnpa9
FHP2+Vj9dI+CPwD8IpAr8gahe02i+4FOqgy9j0oUO2bIHKs+VJO5fC3N2nczdR63NZ6ljzGDclYS
N/7gjtS/2w4JHzme1rnpfPQv7onT8Rgl5NwqaQpGCs+RQjLQspXX5JXPtuDZKOMf04/lMFy6bCaJ
Ebj6hnO5C5cdNzJngzv4Od6kLxcTtFOi0HygVWzrPQRZ0mB7aBjWJ3B0+Y1R8STdEuSXK1MoE/uf
oC+WMSCXbj9bbI5HcWnyGJUPqdGZdE8TzWQcotLz8pO9kqBA5utufBLPhiwhh1oOwLWJpJOjDljk
nekaY7luIQX5mhGMHtr+xuM8Ha4RAHSDCJ0qMx+ry5rftMrc2YuBJzH7sP9sCuADi3jnJZQmA0WH
bQvsjEJOhNiqdCQshCRFv939hSUsU9MMTJcHuXOM+nvFY3ioBVp3N+q+ccukuoOeTBWVY1cn4xjh
uM8Wo0qXIb6GJpYUTdd2biZtRGF+GNzAFGy7WDAHyKpQFWMOLvDTFsTEqDrs9p6u9r+0zO7r1b+H
SEAJKo+0XAcklNKwTZXUv8gFEYfHl/tfoiJE8LhE8GT2p6Ai80Ir2LVn0S5c7NXWWZJ3k+IbHbgW
nv0mii+NdEyA6tAdoGd2k37bwGyTJ2NZuqFcWuuIIov5s6GK2GNsbAaJi7qc28L98vJqvffOUlOQ
7y01uT71NwIF3m2KjJOhbH6/KElliROjt8GR5taMC4Zvqb24oxexD4c++YPD3cLvTKXQPrCL/WeR
8yizR0HJo245PfIUrpdL2QqpoejTbxw/7cyAWNsJakwAZF87+6SKL704+m/EiSej+jmrOE0qURb4
pfCPPzqZ5oyPTNsu9kMm66C35y5Gy9pj71WCtdOaIpV1jJToXnXvrvL55N0fKuEsXp4zRCt/SpTR
KswUaW3k0mBVSx3NDs1iIaGxUoLZdEHLIHjZ0r+EA02a002qyHgfTF90IGWppIKoMVOm5hI3Fkz9
yw3jWFlPMhABaXX1EG5kvpsD+EMAYiJF4s3vAwU8HcsobtwGDRVeAmB6d+dStRC3j0fm0V61lu6+
vaKeT6usqAYYHtfTHHjeAWdEcAzWdLf8bQle47ChMfnMaLuGgTUCznMGu+HdPvQ1NoMDUwljHjrY
2/pPL5WLeBjnnECxlce57m8rI6WierAhqIodeHusO6ekZY68Yw0IV+xderWL0A04EVuUImeDQ9Y0
IRrnfWYqD68xfFyxACz6CjrLgO5f0+h7/vgUhfcE0uHwgmnImV7sOVVoCrfcoMihFSGHveHir3rG
EaqilLKIcffcP7awA9D1I0z8DLMXgEwZbXcaFrP9z4Kndcd6aw4cqSdC8Oi1w6BDVwvAgJJMkkJw
1A9+rVLFvlklesxTk6xAKbZWhblDAqtiTrxhoD0knz5rroC5h/41oiA56uYP59riJRSj8VDoaewO
aai3LdcokER9N0whAuFtzgdhWiWgGoX+kgRW8gXr4E9X3g3oXkoj1LIOMSSwJEge3p9ZN4Q6Aa4o
NrxIHBekCx93kzgx1kEkB0hQCHZmcf+JeywsalfEsZ4N3NWr42mqcR8qGpzggbL6BEGNz/fEIanA
ONW11BUYqCHp15WWUYyukssdP5S5rALC0U1OgdQy0Yr/oyyvKDo8sRlfDpa6TNkTaI2H/2nt6EO9
iWvrcmXSgo5iFvA15S7jMwzE+zrpAiXVf1BsJ7cFb+/v+hKcdJpEsStrPrDz8b3VlojLuYgIj860
2HV1ICOJoGmDRptawDpbXW4JpmOZm1xw+Q6cMd56G+zp7TBI83ko6BcjqWKsmoD58cji5+214Ij7
bCtZ3LGRvoS7JtTJaJiKCvG573NleIPmOi8ZHQD6YXXwE4C9NHrmd0fO6kZa7dd1lbxFFXwyMAEm
e6fAIfuIWoJiA2jQieSJyIqnxJA/sF4Pqh1iNMbm0J3ebtanRPkxC6qTSyM51mLuRDvD9LX4GIxE
UjiwczowL6RG+SREstwmM81n8hv9p7exfhCMSp0l+K25flL2mTOlD2UCBE6n8fiiS5rSW9P1gWNl
4IXSWHjm57ZhJX+d1DI3AlnMGSw6pjP+1Igi/HxQkZv1sxIcHyMxUbEv/kRZG2oirSCMxeabMpkh
1wG+YMF1KhUyDCQ2DjZ7ug3wgnzFEmY1Dy3+PBZA2WP0c8rwKzYPMXfUVCyTCrwdjGokQMpHZljp
bPRiDU1Aj5sIuoPwA0OAMSd/cVJOwvltto4mGMMn0/Iej5Q4xjzBfhsjdoJF4dgJigohUSJAlWat
JqzFU3BL0bBuNi7JQnGsqsaOMHgPuiTIICY2KUbBMHxricKD/2jhZ+ZEXKGWEeNfBRjTboRgFcck
xpJqKeK2jwfUgHpzeFCRXZR/tmDfilbpc8hBJU/NcJytU+SdG7in0E79h5BdCqJt5NhYKmpqs7zl
/IgEiluxX7mD0lUXSgYkOrLQcJw7Xg+MhVYxAwCKxGENJk3fz++VwtA8o5Eko+hvJscMd1sJLDqp
rXs0j4mHQhs5UlzXVIM5mPcbov4isBsBtrsnH7orbjihYcqITHcdRcnfZJGJMM72IDiynzmLQHLz
766rQpRXtDbuVEB2h3E5WcYiQKDqoGdWQzSqua4iW2W9NYBLvy6vSKyXIPmOV4Hc8ZYANjwYOpAE
iETRiGLPhXWl5D1TjSzun6/9iCK1aklf3gnK9pluk7s4DHR7ar6XdqaYX06i5rORQGrRLg6zOu7r
wNZKdzc5gAMVYE7+F8gZ7BOeQN9Jurj5na/ayur9FOtDiz0bZcM/w95wZ6oJBpCRU0RjeTSVftEJ
rnWjB21Curh4S30p/+Optc6LiGHoaFsi+AoaNPm7+KSJsccZGZ8MJ8/dcKd5UTkPnE8jES5sr8ih
fTZcM1q8XaPTXOihoB/VTST5qjFxhinVahzZe2dxADR/yZFJwt4iSWCexT9HsSbuWhc4QK8e37wd
sIPy5EXSn/NMe4F+RsqnQ2cMhGdq44NlHc9XfStdAJ12BCaVrrM0E9Wl5DTxlU3+GiVvQCm8dmg3
LGPAcGcfduLNwmEAoYtC4S8oScjt9SPa4+YIySh48jAYXut9VVj7S+bU1GmLTEiuAOQh9p/59Cl8
oSYleHYCiuK3ht/j+UtypmqeSFJrPpB2KvbF9wh6UScNXJfq0opzBlTLZaRmapNp7deybSn5G7q6
qON7xtWtTb584w6ZWvrBml3sla56fI6Yp2S7Dn/Av28d6L2pvkULIW7P3lDD4VLARDq0lgk4fooM
XtyNRxCbxeFag8BFBi3MGIHmCeoWP6kBlA//J4vUi4OMECl4PDOxXpfOAIVMe3qmJnloPzxuOCiF
eCqvjdfQ6ELCiT8CID9VC5eKfOsnmYTbbXeDFVu8jXxt9C7MH1NO+56/ommzdvxBQJGUH1bLxc1S
AXZHMThXQSVYEhTJ9vY6l09K5o2vHOWgAggzVtp6d8cwbzDFrdl2NtbrlKbRh+3APh/idw32iq7S
UcibZWtIS6azDhRDgg31K3Xt6n6sxQ+usX5ooDNSS3hrsodYgpgvuOoZmGTJZjd3dVsv7bBsjfa/
lI3o+co1z37UvAHwFC8z60+4p64WDofw8YkmWT9OGPCHK9Io7auwynymPz7uxBDJ+v4//eTYqgCB
Bj2sz/F6Db0yrDjSRIRovAUjxdcx0YMFWiXhMGGPFwhWWS44iZjUV375EzlRgBSibyvJKuxQOjjK
G0GIssl540ekWbUXb2Nav53UlN3zwSLKTddt8qC1JIsnwmivbgJ7zYZneF9xNWgc6FcwI3keDuJS
0NH0AffTiXDO1k/VbfsnR+sO+0208kgxDf/5K03FR9BMricvTNEiRGipTcoQgz4DoBeVYchacM25
3OldemUyk742JqE4nXRHoXqNo5PX26IuLECdLdgcz5uYfWdl8kK9M68yQCQsNAHJvyE20rYVeNO+
qHXqTqqmfgd4zhvhhWXvksbpqrzYKm8sFAOiqBhD/I75s6Z5T11NJ727tCX7IQeBYG1itZFVDL4l
TSpYGZyc3nODkuVj0Mq5ztOStpziVvuSlZJoEK+lykZJ2Zx+MJvMt1BZKZoe30d67SgK5T0sUbWt
2bmNVDLSnoeobOs4JIZlcgMOyft5nhHnYpjmjBu50r8kBxMvroc7cKCQSMvOpTx6S7QTZWbW65em
O7Sa70zVguTwhe6n8XEIpHyNBKgCOjNMCY3JhIfV/NvO/zmMlA5/Vce22JI1eHuFgzNtGG2IiSGo
aJdaem+9b/0euODpeSTv7/c4870JPyoCs8D/rp31AOSLd3uF1MNDWsZW/TsC2B6Lud1yMvR+/QBZ
3A00p7B10rvtHbqWyrJPGhNseOG33/Rjfm70ADoyTq80F+qpuP3Ns+T+5KzM9dLwjLbQKVIE1M1U
RZGyAKRzGf8fPg47W7N+QIXOLbSlTDNigdYDtDFM8mpmYMC0nhyi6Bm2T1mZdCsXRffaI3qV+xRI
If3KzBVEmF0U/ZWKYzFeoycSgngvKur9mZsRUmxpbLlSMCVv9Qezo7In1KzYz9kB58ziRAz0uZqH
8zkAcN/zZ9wWWFzc9NmIjoJPmtYy/XW+chM0xbqrPbuO9q07LAxCFMN1ekmfVLgZRfcBuCQ4CSG2
oBL/cL2aAhc2lc7VqPvn6ftGtOSA64dgC1n71qQGVvD2HgVCoD+0QBszoF8rptm5uz9HNnWmySlK
V6xRWVJjK/Y3QowFms6Gw0543RGMxhzxEOmF+wabWwJAHU4o6Y9ySHSkB9XUdgkcRR7kKGmwAUYu
mASE/AZ1NbD/hIpwNnixVTDSq+3i83QDrE7UIryvXwC2vIW0uC14DrFwkQhwrPJ5Knqnu1rsUkL9
p3U46LTKfPBy5YpVKIL3v7D/VKwgEQe+T5R9a5zeYvVcWWUhnsuYdlaeUtraQGxvz1ufGJ5HlC1I
wPrSXBLXC1XdW/hAMUWAJCMKS/hK16E7E0VJv9snsu5GxM6j9NZByTVeqwFOWBNcuLP9ON4ChjbQ
Z8YGaxCz936rAfrykPYpq3y2Sy+yHhyB4p16VGqGROuU8viDGgI4SDPbmY6kZPleig7OMkGr3QOL
iCVdlcp2U3TUtgmMwmHyGCUh45MaUhbkL3yUDJmMt9H0LfsWlIpmBqkcyUHwjd1Y1wtHj9YPGElJ
v/rNaZq/quvTmbDVXLbUKlpKpfXE11TuW1gY1xdwUYJyvDQ7IGCXT4ypEFY0D8udz9XbnI2Wh9DA
JnSGWyDG6lyJWCooB/J9MHBZ7iGTXZlNpClIoP8yk6d85sIlAXD1nEERjsOWPwdTt3aiy8fBRwxU
1IwhkjAYcjpn1U4Ya7zQpXA4cgfP+2rrTCCXYVCz+Kf1NIv++96uG0QzJv5lKboco7nUcOwJo0tL
PdQ0nG43gK/jWiRrMtsHwBWpgpOCNTP542B8u01g2rLMW0WHejVL08ak+Yci7q0xId+dl17BuZSV
n+AzII+y+lsuOLda9uKUe1++1LFfJVJCLGFMPJNhunh0zkMctaW9h30N3QVgu6DIIj6IuqU2ZdIx
5mgbArd9l/pSlxltp2p8yIPegt/08sCD4I1ASW8mW9n53QrKwhjlzULsQtLw75eB930vsZtWOhY2
MSFWAE+APwJj51YJbORuQLwcxruGx4JMD6VnaKX1Cxu6Jx/iBETjO8uepEYg46fAqKN0MmEZ7gNw
YK8C6wkCFdssKkJv+Uuc9JHkd3ZoGXTha2/zrcuTdPm+C0/h43PLCnv53TnOLPityUUJcVAj+eni
6Z9HlG85t4IaESOoT1zPLB9BajaIHl0ox1srTkYhlPRhEw9vcQsrs0Poxb3wjMStzC5bPV2dp/2F
V8Pc+c1QEjRc6N+mvR+b0N9vpWmdEzSsZk1lgNatGQ4LCTS1LcAQHx0euowAk2uEBRm0DF6zNXLu
+vb/kBm4JlfTsZGaUyHCX9PuEAsd4t3JWgeXj4c39SA0QHeZvGRmS0nTBxNt4/LVO0YyAaVmfut6
MIAvndy6Io32IGO332JUtXPGfFCixWhkVNuXx+6KkbyaACHmyL+eoGCdWo87oIdEyx9Zcy2DSOQR
F2Upr5PNz8FAnQKtTCQ3Qr9Mi81I2UMo4I0QA6Crrd2MPKEBm41AQBp74/11ZtR8t2MBrQKlC3D+
AA2F5yZNh8fgZEYLMeYFE3B1HiyFKPq6HgLbcvEsrf4yIgx2f5XsCKlDdjLZaiAe6clDAUqAW08Y
t3nGYNYPzxNMecO5UEskurtY7OcS/H1fGjZrAMMZDzFr2fxVmyvH2VN06RmrgXbuzEDSiGk4EXhF
vH8NJrfW7SG+RKKQ7VJRd/8YxNG5m3Z6ySjWjNPZV1kU0B2y8zOBWhUBF3cAO7wnJS2O1CcE0Ird
0fxigZpEG2vhywuDzFcIl2ZDl7j8ORuPJ/pBMZvQvNIk6Hs07Px8OMqZttnTxK/RNjYEg4qLEf57
2SWh1dU2Tf6/bRfpVO2gUcwWmzuSzxZv7cygPVzNpDcXheMLxZGBW/oQZwlP2ToB/abqwbSd9RGV
j/7wqQp/uDjeAx7Ze1DE/hX0H+ZOFCUfCR6cy/g+VfUFOCWpvQHTGwIvoK/o8GlrkEju8ww6JsC9
0v4ZcfjA2Ps4BVoQTGrWiUhGgSurTpORWeJvYaQceiDmpGuJh5qV6VcySP3DxTFb61rMi2mrpmL1
XiukPAjpuCp/byTum2b0po9w9Iy0L2hP9JhzgiOp/BHsMStJ79tuXfBxmFmK11CaCDT/OkowxLes
7J25jQdHp29IN4UeYapLGBo3KMeo5XFTObScM+BFUVXsc7AkBh/FxT+F3+J9j1B/YaXx0W+HF2mJ
Cu3mu5EmrGeQkd2bBa41C86/tYhgRsAUmO4qt8iqcGnJVlCJWQN9uleDAy0dOib3s6XOkcJIb1Jl
ncc9pglk1M7ihKp5Qj3FkQoPLMwFsy4uKwUragVQUnyvxjfnJMYw0X05l0PGFpMoM8OTi0jNB/XQ
l4e5IzVUllteJDJ8ymCXXye6nzqT5ZEdou/5dqbpE6RxlCLkmnpNufWblG+0BL5qQtH6ATYQ5DyJ
diAWPiPCva+pqAlbMgWXSsOPA2n08OXiUYBjok7EQwCHvQncSE/xYTqeHT4lR3rsFnRSAE+QBC7g
Ya3AyMZibqZNQcF13y0kWm6JpOzAddaaUPxV3nT3QGPnqNifZm/43gz9w4xNjw4MkBnPfHKPGTG5
eLOcqLZGb4GPPgnRR1BKhn28dPxDeKFF0dpXd5lVTtxzGcbIJ1rpBSyRrSqVRLVRTCuqjoY9i3Fs
TyGMAJ9WSmLpT4nrStMbPA5AkKGcK58QEywu4Ovny4FesGFC334YadehGRHFx5aw0CeOCwb5Lp/U
8c9GtTEHh8grp4+5wGGWIPpALuM3Ed7Sn96HyP7ORJ5VHUoptYMFJjTKI0XywzBKQw1Eqa9uGnkN
5sIh0wN2eP5qcF78hZio5AKILYdltubEOLXTTOuqw5VR1d74k7vtTi+VdDGyKOOYyctpZVHxSakk
/2xm3/oca5MVbMQiiqcs/FNUmDHAcBI1IGMw6h703fKIsKSueMJ+R1Z6DX/0uozwa5ntEpjgPh9t
P1ruuDh1ufR9TZMq9AbCu3ZB490acEapRkgRxKdqiV+gynHZgW880g+uErHviF+xbivdXhsKgGy9
Lbdujz4/jTvJKBIXKgvMsW8f/kmCHDFJzBq3n9OZzzoLHLkumjWg/q9mjMEkjukp9D+t4T4dZPcL
EBj8W2GrA1fjC2sCgASwUHC9kvWdltusqDQDZHyjC0/2SwRgdobXgboUPGPnRudLMlesB7EJU1CO
rWs1wzznZRn+P8ADTtf159xQi1YTj02jIjOrAwYWvMuiPx/c0Em17KTjqAoQQus7zoTgmgV7ENGY
kIUO5+UOpGqaXItjIbb56RCcSQTgJFSs7TMd04x5WGZDfJMElU4YDJb6TirBAOea2Cc/bqe88LT2
FlGnnlAfdjHfq8X6/vbYnVtslRhu1HZ7eVdLshtG1c4ppb7KR1oCDfgzEQAwQ1iF+CiuIfQqmclP
CIB9OC1/n6LEYJ2C60mgqpk2wX21vFjh6Ta2kXhsWIrvHULt9paGTN7F5X9+h7HTKXuVZh7adJUR
WDf9nRiNKPw+re3nRbdY2dnaLhX4PtUm5yyAW7lCsVE1rwPe+IVpHnDCZoRD0Pfpu3j2t+uzLf4U
SGzP7VzYt7UDxPrB8TtMPutZtZER7iRVutoZ/WqdrnCNkthvYdFAauomPTcRTPtTL7UEKVE3JPvf
4CZPfnFL4EGiEmdvtlewlR/e9IF2IdJcid844NfWEHZ/SJou7fIL9QtXiNND43tcckEY7TsDD+GF
K5RsHeIkfeW7EIYpZtZkQYKRsVCQfByqgPrejYXlsSY4piLpQbN6jGQQouf9k3p58LdVhaTC3yHc
DMyS74BZR2Vyg43SMc162zOaiK1ov3fi6amOUntFUP+iMyxpjFWIcmVRtj8lAj8TjNJk6dbbx86d
aerwiMy3dxOjl7nn4iqebYuPTMIrEEDF/wdPvaimUC3K7Oy5qkooMYL9O64AlZeKQKKKyGRl8+cd
SpG9SV9wrJiV5NYa2xBNOB5ffondmp1Geauz/kc2voDvF4Wi2t2NTuCBEfu52e+RjTj0pNgPT05p
r0ws3XZA8i3bIm138b/7nrVg4HoezgxlgfE3/5TJ2dSOfM4s2nhkV4daPci/hAlzsqMhxjaOQJf+
shd56bZBwdySWPm6ZBo5/c9jvFhQFnb0hrD1nDZv6QK35+wEB30SW5etzB53+ORnnSiFljduKri7
PrFoAAziCRkvd0puUAJcMfALGOvSAk5bQ17ZRwLE+XLnNUJPVgeQS9NUXWWbsJAIRN4Hu49TvPn1
SXa2cwpeaZpA4hi0oeQu8yszUjbZjGoB+Fj/t6CvoRM8hyl1BSIN7XmpNVRse7ICTq/u3VtyDzHp
GXV/a/QPcT/n6LcXGZx/oR4somjKW+m5z9EOYyfvieLBFKm2ySTfPYcEMxlDbNHa7Z16yQASEoX3
61B6RexOSjE4k38C8jBxaG06XUpD7x14k3v2T/A49N2vq6DqfsIV+JVS+W6a9Glp1bHUteaQPHr2
BEVkgxaKTTxkZNmTRf37sLLdMVQj1T00LBM0cQ6w0GawuV3/U4RSLu0eL3qohUTI7D7SH0RXAl+L
f35sLQkfBKHkOFmkp0ngqbwv5AQmRJ3d4i4niWPWJxY/xHwsOlrYXftjlHKGYZ0l7fnc4FPHLRcC
G5ivX4JwE5qb4UicLUBmLu5FCWw8iaJR+UsJMV89xQgs+wR2NghCAnJFvhwr+mP9EpCT3aWUTmb2
9/4HZtGiSO1iqBN8O4pURHdtSvdKULyvuwNU+W1O5Iz0Ql42V3Mg8xKJs7SJtTkGN/h9XyBoaUrd
Tdp+TG7+ae/B/5HZxArlUVy6h8LrKKffdGN9BCqKxfScRxec32pOLYZAw24SA26PJxjHXqcw9rfu
LtKCEgo+K/CeXB62PoNSHjcAtWE0jch7PNUtTLphqw2FtGgHo9Djlht7g1j2k279vvMs5/FF8lIp
PvDSX4YSZJrsy0e13nacljWxDBXLyrPKoAmvYnB5hWOeA83HSd/DWtCwHCiMU9S2uZuiQhxC7ULx
wPfGIkuAU7CHjKcjs1XQcSVRqMgpZ82CY+SQRe/bhES557txxb6Leip81O0utBXf0nLrtzKrjxgQ
b42CxJs0BkdqgEAiCfRHHLka064p4XmdblwubfNYnkUCXM6/uCv7JQj9r1e3Foqzu2G5kS0BShRn
3ze/3N9D61+baoG2ZuGXp9syUBfl2Ja4Gli32ui7oDrz8EUJNxxrK/3iACNGndvCoIXZevNS/Dqc
dCgV9c5HIedF6EeQ5xwKSnLnJzSsSd/SIADPrcbMiC1IZP8w6msFiLnbNvc3AF9qa+Eh0y1M0wl3
IWWd9AWhRZyxk5IQz0VF9o09m3Vx5/bx4OqRtJPRuBa/+i4TMjkxt04AT49CqgdU72pWL/vdqrDS
7erHLiLtpkE5n4jKfI98TTGnziOkOQMr25z4j2BKjholKobwjThhnJ2nhxsOFB3LxaSs/m7sD0UF
HFZIP37sRc0LAkv9H2588FhNgk9AoMHsJu+eN1Gqfai6CRTQftQDMreXmLH1shdfwEqiu1bFN4Dp
9fkVZ6un+BHZhLqMy8haWprkKa4FaWa5QFT9uGKEyT3/NGJJuw2k6kMmxvz1suk//WZmbSfY1lph
SULnklqgfunjsP21gAvPSN4rMQDshgs6zWGm7bCGhAV1WvkfzmNYP1oxHeb5DuUbrmwU5X5M/MjI
qMZ21VkwhDfqIxPrjrClDDeg4yRd/VKntXDs2b6hZMHTlCTUT5pRjsr5rb/rmsQX2XVzwrHPidvl
5yPjXJ0SOQqJBBtWyVrJahqgJZUtZINQEFrPhEm6d2noegCi0fanGsg7SFUwTwRd7/9Wd7IrwmG6
vJjgdVdxUKKT12P9CmHLSY7o0wSkrJjm6SwY7wsoe2ZrC/5KuBDwmi6yKvxXpyyt9mcWskGC9OIP
TwBhv27e5w4OIoIfzabLCjj7CJF9vFtpQsAUwJbJzdp8+RHDzRgk+gIrQfjcSM6tYydo8CgCuHar
z2FJKEyrbYaGeTiaC59xnTRYuBoL6fih6UyzhnhRLQQ0kbFwMcIP9BhOAZkJeZ3RZ5THqKabdQoR
z7LhGHtvggdoyN5noPyAK11PG7Oly6/hsYl7FHEahMHiGJty0v9ukwU0AYBBVoyjOkYyMzTbEQr+
Jcnzt13R0AWbZfnsAS863JuD8JesK8cAhteM30R1WdA1mUqb5EVpw9aiZCXBZb6cf2Scl12Iexx7
0EUt8Ud7sDjpClmYPnSeJ9baFJq6nRZtIEA55AGmyUezrUW7dR9+f/pIwGGpSZX/YCZ66ZXQw+cw
unYdEqgvBNxUzGVdUXEVpPEsv7xSTudVqqP2atTS12G9pi5+eBkbmisQLP0CZR7dbSP8joucquXk
AbcOsSA3OtD5dInc81M8hT3LonUdsUFnKYjGUjgrh2rFMR+iC8I54tFLVPyT8Vw5FYveh35yQ7eZ
9vbX0AwtBfkiQA8bINGCRPM4XoNf6Mmbh3Za+7oapo9ijNyqCBEiTomVmfUtv2sJbEDJsr8572PW
4pCLaMmsQwzxHbPX5MGequSylZju8VcXZSFmHQZjRUK0qWbrSIml6kQ9Uv2L439XyAZfJgXLgGT8
rE5x2zWjwiEx65rM5TzSnfk1Fkt2jTdJUBDnp0tTIJiPO9O0siwPN2+AXtgF098oivLmIcjOuCXf
RSl4DKwDu7VyK2855n2LJaq2gmacGWDdXVr3UUQIAS7LXeg7n7Y+Yhc58VS4SvDLP41dSGq28Grx
s7B4j81dGwjMdnsib+4spf81ucpxwi66MGglPq43OkCmrTCG9/+D1upW4paT53gyU0TrZwXofGzp
aK+gbQuPf0HQoOeKj9iwtuvKH/gWZhh+MfZvCu4RfAOFBzUJVwTGI86ohNBhH5FuGSP/YV/jlmAx
5PP0YsIKBKuChM1oIPL+mRU8xJHysBQshCikE3l2pmXKYuqsu/DKNzjFrTOXnrtTA+RKKTy8nuI3
UnQGNcNkp4ESp3zeoVoquVF9XHOTQWdvQw3qGeLNuep6OVUUlW5Ht6XS9J6KzRC612eReLUotFA2
cMUjFqhZOQ6aQ6svaITMasgavJePxNCNnBi4IHUpi07ohuLwYIgmFhOD/Kn9KCFk4eJGkgOsVsFZ
u+jsWcHkrmMfAbNtzAKWJ3a/9NUkowjvA7zoa7H1ze9u6VTp5rj0Hw5C4Hg1aneWe2MzM0YgxaZ+
TWmg/p3D8ml7L6Hg8Vjb5ebJyIzXeXSigTQPtsEvbRFGoUKFcOKWCLZWoG2PnLUC7+ySBgpf4/qX
MX4DE55t9+6VgdhebzrdRh3nCcVMM8WLPGMHns2dQ8N0OUXFIoZwNQBTdmzkeFkTioUWFOjes7Kk
IFW2EccQdfXv73cJYRHq89wtgZbpLPSLQyEpQMVMmQFmqJogrH95Vx80Nqck8BdZk5NaxYJx7/l4
gS9Cwb08HrzIrSpg1lhoXnt6h1JcgOW2vzIpqFeJsd3f/YhOu0dxb7aO0O+ASk2onML8qRduy5Gf
0CuNcdQPOGH/wWwkKhvAEtrBdTV3O74/UsZJUDGoX/C4U16xEg0cjhAH/4U6UyXc62MGMthFJqHd
3JJpxx/TxzhvCXrnUbh8tmoPdi30sBObQjy1vS1xmQezSANVC8XTK/+zbjvuP5oMwj6zdqfNZ7fG
bTQQiO1N2Zw1IFi4R66r6RRXD5nY6CeOqUhBaQvDvuvppNErYbeiy2ECMNS/6WSNECfEpdH4PPvO
byGZ/KneOx2RKJDe9PLWKrja4z32rtT3s+cNSSeNjlocqQ+5KMsFsteZg7uKuc32ZyBltAxUCs6P
9DvBcHiGhGukewN49XH2tNjLDokB6WBAvvO6j47WgjKqJwjj5NmwhXcMiKy13Uif1AV0nYnmjEm4
R8r8QHunDBp2emHt1BAFp9VX4OPvQ8YF3koRbvxIXds2fO53T/WUiYIom7xEisfiHGx7lCZjJCco
3encl37hj7HeqSP3Yif0Z39rwjjlUEUb5zVwEkAQhXrHnhCZQBPVv2vw9/FHd9n4MKCj7r+TsCOa
El5dfYIwzHkivul6+uFMa+sBZnnNTUoIVjn6szK87RHyyqu6yCD03cQXQHJuMzytw09NnPt+4Fd3
d1rilIWGIsFdiKY1qahxtx9uHdkCaH9C92/WV/XOASfW73HkhZ7gahVo16oF7smkH9kjRbJogGqK
TPnPGCZTaoF4rYnwprOvJcUS/BMFVkhwbFJoEDMRtwqRMp06qO71aAKTfcdsnI931hlSzT01Fr/t
vyh1Y0D1euWV25VlGndkMd9bVVnC6qHGBlN/STNF8GhP/rV+iKYY80Ge47bR0Aou+7YCzmXlyGQJ
6KRWjhNU6iZh4kBMModR9MswRiBhU4md8VuT/TTCc4k4rP7QSisqlnc260WNHaZgb7M02FLawxmJ
utcYtrIihTCRi0U+dmi2wF4i0r16XNHRaBlGghKiJdpSHT14ZJ5+vaalan0VTr9pTxe+e8XuOSd2
G+69R4O8MrQ1WryBswNQo+wTKqN+68JJw8Pu3vqiWP6uXSiE9bZ9iu5YsCwdqFAKsNfj+AId7gQh
HvrY0BYbrI0Ioyd5XWEXvgL2l/FjLx+eop7xLD5CA5gH1fPt32niH/Xpl2PfO/XTZKJhZVrXYutp
lve2JlK6IGoFx68PWW5+olXO2ApvCslaNEKC1x8b8gTrC7fUQjylMsxAaGvbKRaWM765K3QpfcDK
MvSXUtSAd2Hviq6i45XYAcqgAtwUd9eQSTB2qBy7MVSl/qIk6nNAzLh7aD4OZgCxpc9WhF2XcbeB
RI4HVAJRx3VVtH7zXPe6XBD5LAFMHI/BvfCJmf30DWiIi0X7ISMXIltMCcyIkojcpN9InYS8rVIa
abWEHdy6Y8Kw3WK+eAOEmH4ZvZNXrhp1ie5DvfAnLcNycdXAO+1DQGs2vMQSy6epmk9q1JA1RsRo
Ks8ftUciH6UIwKReVB/YaGesPE5vXNYXpLlx8T4eI/xFBoCXVQaq7VVN60v2HtZmLhWwtt9CdCuI
LU+UBXfsRlVjfVF8Z2h+5vPR+Fu4fJp2B2NGKvNSCtKNbNLe9QTwWJZLWcOWrdRInTbGXLngZB52
Al8XLDhOivBtM8/KW+2eyhILwrQLzAwDzQTK9RCjY6aHtU6YDoKFk6onJr9DIjZFe4mPIt4JhbNO
nwxA0mZM8Bvaw/8A+PmcyQ3Dvb5bhQrdcdwCFYlNfJNEHYwEGY75WfBvdgedbjI2Geig2dHBqNML
8RWD43r133/KAYfLkpeTeEw8BsOA7WhtuYmU/X0mVtiNaL/EbdhfJseglgKWQoJrpHP/DrFm73LF
g4SzefSK4tfRidXaKa8kit0zf1MhU6FLj34uJ+YQMDNzwCd5iNoukP5BfDKaEX04MrcK9Av6c3TM
aDxAkYretk3J/kiJVd1xCaASjUgPEiN22JocGIC6jcjkUWko+5V4iIZ428ZrnUtLuxR7gutsjUiI
d6lIRlP5VxCX3MWF+hDSj0zHWSqpNh/xk8AreYRw3PUqezUX7bsZDMEY1E8P5mJTPRErPl4WyQ43
8yyFi3QYXhy8gNDCNZ2lLheIXmRThUUsZmPSgSapZbTzYtKzYb8wEzM2BdN/foRUppVlCkT3DsVQ
BJq8oHxanq5Fbe5HkM7ioEu/TCvzQ6z3hiaqUK+3CeZw5M2KwWqh2Bp3WFi2/wHXd+BiNn2bikFP
/XDb0CN9CPXKwy9iKUxii0Eqks5xHB+g/pIOTLklO3MRPZzOxxjSwSHBujHzQjisrfLZ4JVMhcyd
t+YDgKByvryHMr2UpZ4Rgk9MQ65vTv73u/jQroZzV0RaiLEXRZnzIpXY8WhLfyyAj44h+9D95+/i
Vc07bSIEvQJO77IN7SKpUBX4xS9pMFuOeawzE6uoclBOlWPYnwaS+a1fj5uB5a4Ihd3cN42Zb1UD
m3oQwPQgwz74kp937U+jZPv21ygb7kFSaskIysZcQew9U8XdC17JGscy/0PuqySqbsAJ2gPbY8bw
CRyifIVnxLXnisKCs9Fuijf4IoISuIfbNAEcoTJpLxciQPZj3Arhwdw6d7k2BZSZyYpZIfWX+Ds2
JG759NNn2TFK1+iJoje7BTecrzgEhP6oFJAq8edbOInCTOE17JQu9nxjbeZTn95VqVXImoFsE+AA
prVHZ7AeCE4fSYIytQu1HewUHcZs5rXaqKFk+Unyn5KsOrbP5td8ld7HLTzNhrEFqeyxBfxgXnmQ
yOaHIcbzijoDqpADoHC7AZ2wjEGnh+czljl6pfMD6hlybZ1rQoBcnDJp//Yr1/7TlNBYhxsD4sKH
F2JD3zOz+AP1WSC3iqzBO3zgfEQERE82wfFN5jc33RT1p4OP0q9RfHgXd1KmnJzLdchWAaFF1X+U
L/useqS5jQ8+e2NuRKQmYjAyn+oqFGqqTj4G40nvyWB1MC/++Nkypwb3CL4/ssc5Pf0GTZsch5cX
KqAwUdEuA9RGtGC1MFc5SRCSI9j5g8nIpcahVUfuxn4xRM2TXdWvNLmoViD0kFx+0Q5JXI4DvEgR
UWWWt1JK7kFHptbHpGId+Ukpf9U2ab4++VX96cyjkMocgGKDMZhrNuNbOUcQgGswBKUPOhubplqf
zCF5eRuOUa9DpZmKe45wRRvidRACCq2UAlzrsMmpUKgWgY5aEoR8vNeenYT+jV6iCSR/zsxDdbmH
SN60F/brLIh/bWyMpS29iVNv+8Fqjhrhdpnw4txVeDIAIRAiZym/x0BTb/OmpBod8OaGSk7Sc6iY
fRFW0YDUjxW8reV9k2v41PbKRb+hj405LQh1ZOmnRkoi4ESZ78bvYEXjgSWU18obPluUtAkWQQvO
S48UJ4WhsZGLjRUlfks7CoMmwcnGVYEX3Qzww69tFhXMdVScoR/foeWrKEH6l2TVV3Suc9NFASM7
+Gj4E/nZk1gsoTbk5MbVmQXvlosGTNJXd7wDFBE7FQ7lpasy2KPSPE/ok7bK+n5AIDvJI7Exj3fE
GneS90gwdBU4Whnz80xOIpEmiEZtAFtOmK/XCJ9GagJGyk/jiT2jJtvUhpqoBuMyLlKUJ2ToDp3G
EHkuuG6dRvwSo73Vxunw6kJ1rwS1fOICMp/skme2cWCG6T+wVZNi7RAfN69fooJSSoeTf8VZwG8N
RZnIyl+GyFG1g/AzUaKyQtSVHgyYlqEUTHWDh5mnxom2InxhoiG1vW6K5A8VfsctcF5AxZoTEEJn
8Kfent3mboADOnS/PBY01qWPwc5awFlDh625RZlYtekNo9Uy7sVS0UZ6UDA7vMCR64UbdND3u/AY
W2viJ/ETw0ARr/vq/5BGlJm9v7J1qM3YRROz+uap+YvYDrEGiMWH8QPmTBKNArEFcj1UrHnwKKRx
Ej65blLvpozR1lr5x4pXElJHRDa4DoTwKO80gd2c6OaCCcnQWwdDNM61cPcSBgNtcl1pIKsZ6BCn
+zq/H2Tu4P14gOu4JlmfhKIlPEpVdDrsgnmxqrl+1XEPp4gPOYiv3RkfjgrSGXRzX6da7MrHyeuw
QLWDni3cunPORe8WKh2lGHLX9yMLrNGr93zSDCv5amcUJ0OAe0IMi5IL5GTaxrklL6Wqbcf85q80
y/8w47R7kZMgekWNMJDOAYt/t50LnaHCxMoE8lwFGdWE8smzhvfWlTfE/MZR/hba205gKEjYVbbS
PuUOmw3khlr9pVKTpWuzTACXWJxW4Jw4ZlOuXSSDqlm8nJrBfhkZVdk0P9WAiNwtGdmDO/9xz6W6
YkS2hJZ/3g8HHmUPJJ2sUnFROIxhpR9wbW3R2oXED9ADNkQeuYdW5bKLVbGUjsNaInHzRJAEVysS
KSjiVh0VogJRWEN/2yXSkqRD8altfmzHcVYp8ecldckqw2FlqMSJ9EpjamTl/LtWa9hGuxhcPsiv
g3e09oOxqhj5JARrLLZ7fv08GegBfQfDb7dVph8VZsGgEUHvESOxV6CcZCdm2zkxYKV2lfuRYXjG
zJLgA0mlwQCuuQkbDCTl4ThNIlU0UaXIEtqXqexgBjNoMOwQWL7snyBbAYQ+fLqkER/KEstuhyWv
dFPwx+s/tkCETHHp7tVO/wxlSNdn2XpOSks1dYXEULZOREZ0IS5sudrrTChSl7SmMEMr9T3xmNZ4
1GGye0ao8zajh8ElBDG8X4RVZ619PwcNZdnmp6eIKqeLeOxcnFfxGp0hXDyITGQ7ejnOTXUdLAo5
yL992Mz9YtHlL8Uy+NyYkGhT0QsePtr4dx1iZ05Be8jg6o/uwXcZaLrCONaqjwHcyj7fKWof1K5b
Wn+jlnA/kt+6BSxx4YYD1NNgjPKwfBhs44haQBJK/2LMroBAhQImszzxSd+rG5XyeSXOyniV8tH4
aL8/tg8+HkEXFrTMlBzNAUsyiMvnwhGUWkhfdbtAyMg4lrzOFoISHTRJi5dSIaxVfABDN4GdyuAB
/7MSkqnM1SBQR6Eaa+z7eTKUNQOEtdCqcpePbIgkDY2gbUnTURSl/sziHrFlVI7C/jaXwE17V9mE
SL+HlNEIHZKXvJ6cu76LBAW+YdfXYoP3+tB7Kq+ASndewuldvCzzH1kIwiWD4bxNlT9uDQbSBisr
PlcvNjr3BG2vzQvslva/G2y+XRBSp3eGeh5BH6rMb9m04tVJzkagpbF0lDoSh9gMrd+5acKDA1YN
wnrLDkdhbPMt4f7hriq3eQSGc663AW89fC6dIC8ZLaVy+djIqQpC/OQhqGRocL/QrEkg3dEcBRDt
wfK7zdAiMTPlthAOY/XeLXK7dPwtA7voN+X5z+3a3dspqMUVI9WtWutHLeo4O2wnYyxZeerSbL2W
7TMkHG9HwrDxhz282pzs2gMbyOBXnXSFmgRBgwoag4zow1UtlVHCIpb6ZNQHN4ms+rHFV9Wtgr8Q
xmaQuI8aUGRiqDUWdiQJjvqJfsPXiDyOWcqtEE7UQaLYDDqHLq3A4jlhbass7bG1RK75SrY2ZNQ0
ZhiYfnnwuGuMHYxXO7eUkZHwwT/j8i8Ur2sdMXLDadjt/2c+4bTWeGvW5dOxC+5rjvD08K8wK6tD
51DP0Rr4kfUWJRARQ0BBkkof7dZtC2vymmYK1wo02+169YJWohWZaCVIr1+GoEiDLO3G6WGZsMUs
3FV/z2V7JGnSCmz5DP6vk0R/DUA04//vvgz8PwrSCut1anwNXoUDGkHbXpDH0CVEGB2dbYCPIDPz
RZwmRIshcJcnqHI13y7SC3EF/DcfNzyPsY7lqkR9ULTYlTIgC89D2S6vB/KGe4sjOSc01Axa8620
ItvdPMcRoXQ1Fz4afSGJDcgyNRFdSNqbyezOP8yjnXkRe701vzGPHV5HQmXgH+HrFuPVCNv8ph4/
2z/qjXmKHgzHZJKD5zykgLoA66Hr14WDW3c0II0b10+vHxdfWsEHG3hCHfNkyk8+sqBth9u47lRP
APB00QN2f+O0Cfv31vAUzeVnrgbtm0PmnqF1BvVtsJtOd18HqtzDDP8KZ3qgD6xhv4is7Z8yWKx2
pGj7Gpk6/cciv0rv45IPP9FtHKkhL3MOXDYFDq6ZVp9D+r0mhrpEyBEKC+Zb9Oq+EEDCZaBx/kiC
Xq9/vqaS73mthiehneWXH5sPJdqXCmqdZ+2fZwO7eHmIvhU1/uAZmSFl+ExPWwIN6e+mc0Jg8oF0
DuN9XMTiHJ0R+NpdxmyA7F9NmswowRklW+63KCTgNxYtmiWeZKfVEYLjdasn2jSL/+OiiRr73nfD
fpXP/9ReOsZ2A96kDpzE6VNzTanrHn1xNH0gnICNXsfEWKkGfnJb2XZGMHzL4sHph/WDjL9cWg/N
KAbFCihL2i2oEuLcVmUT+sv6piNz3TO+U3d8p8NUgJDIYg6HKZcWGZ0OnGQiRgb6qRzYIUwz3Pjv
WSEgMX6c9D1uRxiuDOygRiojRBJ7ZWomV2Fr3mDRlvQEfn6OLKIjwvJ2wWgUAUQbSKbzZY4s2pHe
zVEt1A+qctoNFQmQlPQ6ANH4d3UtY/ECsdHjx8/VBMgqhVebYu7KsFvtg8YmOC72BY4XQUI63pMD
SNwkfsY++NxEnRjLAiY+//dwigihI050xWF22bbFev7QZk2v3ltlVTNgD5y35oC8ww8kIgtzl5TK
KtrjqV587cAK4QI5kezbcdhil9kIsTR6qoSdgMWAkpQC7Bji9jiMPpctNWpindPOaNl3xU32eum/
stmZKYMA6SxJwIjLT1PYSK7fs0NxKqLBz1ehJ+LFjfptDHXhwodmlQlfDEwcv7fd0NK4VKxuxpVh
NsZHw7W4LiMRPc/khPjF/IF+BiS1b8UfPz7/UOIrR92Nz/MZnBEMy/q+yTC+W5AWvlDKFRobgBRF
pgwbg1QLYcyoAxVZmM6a9y3gNgJhgrdmS5ov7HKrg8YIkNpELsiEFdIH6mGxifRkmeQIsLaAg13a
9yOneC+FNvNX0ykXk6z1nBKZ/Xw6S4+b5M3S2Xv44/UeiRIZy6UKUTZE2tDvJB15u8OQYHEUT3Bw
r8kk6mBhoBD8KpNcLnAL2cktQYpsuX798wgOxdqmF3NaKUG1kysCK5dORUtvu9APrC9v9jAw12mx
4Gdl1NpSpkcEbt/ELvkcFQn7RRZ6vpPNY6yaMkWWlZcfJGRrviuPhqDiPsPm669vhz1HFoSEQ9eI
Gp0As1AxwcIhvBqdHbWDT91+rPdwruy65/LGzfCwJnYiamzhtzTocIQH1FHr3xaOVVV72vXgzXno
JCXHrOP89I4uxJTSrV8VupCXi8gsopZOhC8JvOyON8jQpEde11pZfnBJyNaYoDCVJHJbYIZGqyRf
1T9SBXLSTXOVkBZ1lrLjUGzzVejB+Zmub7rwSUByVpxYtPa0LOO8VAjgHFSOXnviEPFf/ktCDg9L
jB4ML35Ir22H67y7uiWKahYWVu22bhpFMrqjlAiy2yMfvPPYCCd2d8p/LA2CNNYmK/QaR3AzXBl2
QM6Czkz5BCE+VV1NEcALzHFbi3X0icUG1UTP04ltnW5kPKXu2D/ZL5ZZcBlL/ig8pi7zNuAilCiH
aAwb87yts0JzbF+7ZnYZ9Hm2k5CHR4fo1WZR8qQo+LRstDw6jMiZ0tRE8SkirRAEPtCBrQO0+Yrf
LGu1VlAX6cPvXf1NQHX7YJGRAQ7VpiNEJxQW4SZVhDzlcDOzzK2McpGXjoQdIHH0zH6pjcy9qr44
dlEVUNmYYzo6Uj/+7IvZeXPs4HdOu60d/hhRNTKvROYCV2eCLTvpr75h4ySeA6zmNoG4KF/Jac5c
A3K8v2c9jDkT7zW7GUELi5kPmO5rrXcoBDA5YZhgqKSeV6ZsqzNPJRSpJptDzpCDEZ6SR/OVrDqK
i5XvAnURjhrVjyGJGbkhBiczXCTPbAAdL2yShsPZwBCNDxVJLqMTTgjDO2tHUT0xqNknn5fXmD5h
zRJAQTf7Rr+XK1t09iEUgsmpM8For1enxr8dy2ojGA6YFsHMIVk1fjIZUfcPlly007khIE2gGjbk
brCSirawtdZr6hLZGuHWYDIm0YK7bIjUHCyytkdPSAl06R5A7YF6tltWwK7z/LQVIO3MGxLzmg8r
U0SXCjPwkGLGqwBcVtvVG3vihDDhZlY5fip9tRPDQ3qp0vQjjmlvCyeH/4WUm8lZ9d3x8CL09+7n
8+lRRqgz9CVV9gItQp30xFh0ExVX9oDHRDS7x4r90jHtryVlxSmi1ayZBO2sSp9ViSdN5BFuMyfo
sm5PUG8d42Y0Agox7yjD/iYfLgLMsEwixp1QtUqm2d/XhvVmZ6CZRXnDqQA17zxJ9dktJ27IyWbT
4QsJuyyX14ABU9RrA1A/VvSlFcfT3EzeUhgVDWw82d/17xDMRdYG8R9MwTvbJ8Piw02Ognjf7Acr
XmKcmlyQk74EIrLGavSZ/yvHJfaPwdmnju+zbZmjPvOj9BBauaOGS+PsI7A4TglfNZsJGlD/H7N7
H3NNRI3y/keZT15d2v6ZTBVI/YIi7NVf4MtZfCOGHwbyQSempOnWjZ8aYzcyWoPpyYNxVec6vvrT
Z+8uc/s4be3hLxMq4tDjIZwtarH6v/UoSq4YRcarDutVPUqX/zbv4CuzYbyl3QPqLpugCpF+OpdA
WeQipEL64TVQVVXQe79mTYC2NWvO2Q3r6tJbHNCm5MukjC3SVai+BWNvsfcgYKrlrBpVyM+ziONn
+ZKtpW1w1czWBuyxSzRHXtq/ut3wuPgiprsjaJcBhF0kIjZHzHEPUthvCUUTNYo2tYMIh/njJsa0
sgPmiB7ians0yZqw7+VFggkS2jZt3lQsDp/5RmY/NfX5zbFGOlj9vEOt2wFdgQh1S0q+IZkvFimK
Xt8Z+qCmNXtJwWS6sDDTTwyMSV1a0vTCa0sG1qnc5rYXu7HodLCeNGHLYI67PfyHaisYzy74ZRfM
y5ODiD4Wyn0FO7HDG1z7euxyB4bU9oM0+WKNL6WLWYLhEWHv+52IZvRgnZcNoTPsyNbTax6N4QjV
EziBSPmIrmQrLR1PfPABA4kway82+6GT4YgUz6VTs8PQs5g5n8awDEAQbsoQCJ/T0vcG/YSFYa7e
n+lLg6V0cvGjVmG5NVNCyqNvxc7547za9lIndKFSi+8FJy8WQ2j1hJ9fBlOFgFR/QLbTVbewHAda
VH8o+pnXFF75aP5VVL6JjFj1ji9n6N2ZGTlhL6LDaVpBtlPH6ddpiOEewdN70WGc4ur8Bx3dWwlj
7UE8ygTZ2YalQfcT1RylAszlvzPrVOpuZhd+zMJigGDuKD8CZJ/l2X+le7CEeMdOd/NZ9f7T7C3m
SzTyYZCHG4LG6NyowTFDC42wAIbeISEuwxa/dkFTV/dBwxoIIuW/Yum04Upt3fP0vSRXifkyW4CP
Bl2GTqqKWrIbOKvdllYozEoFYVqjLkjBFWj7AnsOT03NcO7BMnv23yd9CDon43vQj8nSNv49UDZn
ifUsKY7VgBP9wmSQ4xDGv/QdZO2va+pU5smSdTmP+kj0aNlVXqO82HEopEKriwDCemwPpo9LtMnH
5C0gd759CK983BWS1Xvi+tkR3kyYDb/u/jPXx/ITgcNVqqSmRyytN+3zfW/bqbzm8zG5WOiaQoZM
1YQ1fI0xVoL4bH8I3C+kLt0+tECIXUypX+AIvk+T3i+AparTABYjwd31NGuAvsQcZsR0UWACwaP1
9TaOYBJGYKBc2WY/04fLuPp9TQfC6lhp61djOMqr45Jg0IbraowPm/TfsgyfVvz0I16AO2C7/SqI
dMmHFzEMyeqI6VWtuxYdHdg7dMcBU1dtjwpGgp4zAH6x0vPiWW3Su+gDgW8grcIH4Qu+4EUndCFj
aQ02m/MfO8d0MUT6CVTINls3cn3L2kJQXLUCKkM73S/N+KOSZ2CS07nQk42gZwEOkOpnuxGzOyxh
HzxA989N8FkAwE+fHDRQiwDZzvvenjgj6w9vJBTuG+2fAF30U/ut9O2Ec39cgHPnVTplwHQzOeyb
AyrfJDmpO/CJuXr3Wb67ac2DaQatuXA4ndJ0W4Z1rDwEAHrAA4X438ej+vbg5GtNgBz7tJDmwYqm
getfApXCElTcehW3FA6K1UfFGONSWrX69CQh4iO3ZHfVZ74oRLx2dwiklP8Qv30bQCyGkiUiaVXX
a3g2RHhPLDMKSkS2M8pLJBVtAkqjmezHy+uP19CZq7xAMsBZQ/yI+Oak202uz38xOq0rlbfpiM7x
goBYGWP4f7v+Kodfw+R+LoQoudOPEfJwIoEyMYTAn/YSLBmAWQO6JI+DZQxKKuCv9jUBUYN0sk5c
6HdnrIloRCENNfLueVcvRDhdFXVvYlFlE159nws+XPA2ZDnnA8XBYU1yG0r+SoqoPoVBzXJyx2gs
CFn9KFgHvO/1XKsnQiDjeuDAlOTi2pwJGhm3GH5wjFP+Xegc426+xSK4Ro4Ch3b7i29QAEXwIflC
uZUiWH8B1uK/i/UKUgPAdiptyHFPXajwFVE7CDPjpYbcfpDcLreRP4U4q1TJCPAwmdaR1+hN6rcF
AeTbYx086jvdK46MLCXzJiPc1xmLnqISwoMJZV+mL/pWNaZXWigS0KHhkEGxI7XVl0GPGs9IcBYY
2vshUurucfwSAHQzAZ2oB4iYmvzfLFme6bnMT0GDebhZazi29sW8hzAAKGc4rgcxvgs/vAZqo5Nt
6/J8W8lS4lGwZfWn/ly//YeJB4DIsv9BG4nLjrI/c3d9bbUfuUDujjHnzOEyjN2UjxELzERKFPen
571mLJqEIa58oIMKXjdKGDWun93gfsKeUjBqP5gpDiBX4bkvT3nhzsVkRtowpMU/6z2BKauC5DzD
xZns/q8L3z4GQ8fXTDLrybGVxb5P9ND1wX3zZMFdgm4F2lP4zfhp8QIL5levPCaG+Hy7o6+W8ZIu
QRc8zR8gWQVqrfkS9wklqFShgQFE7Ns+w7UUxphkBlkyWvjMCkID8uFtiVLxwdf6N1cXH/hx3zg2
Lh/Cc4KpqL8HIrrEfOqHbYnOK+cLMhIleIBLm/1pDvEnF5876HUO5gsQ+iRxCsDUUhCqIt95f6Ab
mFbsQG4Du01kT7Hk+23o9uU+X6dBKdwWqAKz5avxN8AwVxVSq4Y4yXBUH37Tya3cHjlpVMQVzvGG
CN9DvWX1J5CBbNfxWGaCXPapRBBp8Xr2+9lnswbLwo4Py0rhqe9F2qm0/9+CA1NOha8NLRaKjOIz
7AxdcQmEHd2fMjgxQirr3aPBaPJPwwbJiwern1TJgr2SfnIkUa3oovGA5ldnDgMyhNsQaog96czA
ih+sBFTS0lXf3LxMFeeUDG8VEgQwVIWwCstXeANp8DBG7vLRgrA+c6/ybQoNh6JDkLeLKQwEF7SB
sURguusvo0S0jCCBD13gqMx2vhmLJhbSpdkz211Sgrh3a/YGHztu6lGVhW07eNxuFQuvcN58/Lpa
zR7enk6fL3el/QyxxvFvY7ZsvMMM6088frwyjC5RWWNGLaSS4M3sdb9nRwgG2etkxsxd3lKQgsjm
6GSnDhr6+kXfA0fOprqfAItghVYA5k7wda3mopMXutK8k9DGo+ndhkJSxgDMF3YKkhJMtzFtTgm+
r2Ye89MjnEtflZjOcrezIxg2jPf54Rt34FMDFEDDhkENwiyOGoelYue0v6qVunQ2uQAhEWJFyRA5
+r06shHXUdIxBw0t/YJ8XAxjIcvCIv91Ox09C7dwWnCtz8/SO+ta6t9nv7zGAKxfG9JLdAnHDe+x
i8tOZKIFdHdi9Sw4BUxzDloDhjllSnSHgSw78yr8MgOr3EUtHngqb6fOni31mrtmz6lvQee9djeV
ECJOy4+whbPm3ILC3ySPcZsI6sUTGS09+a3NrLnTX30UKy7yOm8PfIhRIn7PyHya3kjJ8DAsXhHk
Z3n8zrqqNoQC5R/pntIN8f/oRg2cRU/uKPxJe+maO0/ONrXaMgb7XoaSwJeU5kCDyaopf/N9luZQ
VdV5HnrQnee58fAhq5MMTukHTQBa+28GB8jfVi5iNkLb+539QEiHsSNhNf+WecozvXAEbSayGsqM
tX0xPTa0LL+XxDDODYZDdf/DDDBFAONwmQ0viIM0lvN0qHwVzuAbeuc2QU++++PbBZnzCHxEDriT
U9sJZIaz/u7zHoWAckPM3BvmXBQQWzHcazaecvZ1+/pkYQVMpdo+JSMJbYNRZ+coIq7iC2xg/Qqp
liFp6rZlmHPDMOvAkfJAngfrVsUAYoMmmDfBj+hAAVN9+DjS99ef0grvkYAP3TLclzpcLjbkTDke
EulX2JPVHWjK8/It4wYfhGMmEw5p5dykindT8CDwPXKf1/bpKwvAirMRaLqdNZV7KoP6JW0WQTxp
5MdLzXLamLMnB/rohhGrKKK0nWNdymGjjdHQ4WuLo84Vs9FaJajn4z3MkHRqN7asCM504uPaHFYx
rrx5L5TTp3wXK6Ka/ECTlZKqX7BfueY8yeSe2FdW3iDRqp9oalc4+zwNNQVjM25rXz806Eb1dXrG
Ft4OFtY6G+bxQhRz4V605cSxA+NknG7pdek8NcwyCBE8M86FdgSUwlx7XqU4qUe3DGd9NmTpsI3v
LYjAqbF9TFnWTDBcGXmYQrmE+QkTRbXev5G+ZEdn5tBEB9xpRjSxsuBrBS/0pwJ25sl3J1h8yE5O
PzjbOB2VODNFu4zX8rrRz1EKtogjPJXig3KV1mnpjYpBJ6owFn7n8bU8k8vQkl59QIGsk7wZSpmi
YjNnv5rhybqgvYRA7C1ThAy0M1CNadh2JH5ZGFMApElcU2gW8oUT8t51Lo2bALOr/rF7Q0KkDtxe
brYGkF0/E5Bx3yT2IxxViRI7g5Qy1nqajNodbgr/vY9MtlSLLtfIsinw5iAQF9OY5/OiKT3DtxHK
Yl2JXpSbYoTgqm+riBzrY3HrKevNFHLwnfS2jyplwL9ONiRexLIbe/sK7XZcLESAiHAQbmngeakq
YFzOloKQ/p53UA5zfXTV/7Yd/BVp72OExcIRhHmzbJ6GnSTfQ3Xtxdd9qpJDNpZXXxjSJ/c8PkRw
13cvjnPZfGIIUu0A2v8qy6P1nN09x9Ap5C9/4mp2w65Zgw0pgOBz5IYqbwoR1sXHvVzEX2Ipm0EU
DQvR9XXaQ6BfRlIMRKVuIdTWojl9FlABnQpkKSi5zxMrPrQSM7ixGkQlkfkno/Hi7Pl61Q1TzENe
cLvRzW/vmMWW3LqHYXLiAv3ZaEDnp5QsnDjTtmhknBfu2MpOE/Ccb5WAkuhdgXSEJ/Q0J0KujVZk
+EgYT6Kq+8ag7nh5Th/OcT/u5ASY+wVQml9EDpZX7P/CkPHN2qg5V7dIgfSzMsfb2pDo0JDotRvr
F6VJMq0TumnuHjleW53ZxQ6cUpweHqZtUIPyQ6TCwkyucjnJT71DfLO7wbQW/5NM0YI1MVJEPJSn
KHEgPsFtw+TnAZbepo/0C+/QkY9xwgzMbSXBaxZaNi3G3I6Jikp1g3QI0wAIJGHjCDOgVDFS2ldG
IacaxJjM+n3bYdAGw0BYx5A+O03Vd0a5arwuR5gDCO3LE0LHdMmU/+uw/BpFCvIIKmRTV/St5qik
53tH79oLDTO3LKpmQAsc1+q8vFWZ1YxvQvJSQEnjOlOuzyG2/TITTukbeExoMDrwW2hCnZ5d7wsK
Ur9PQv0JfWKNmYb8dusfbGhhcaHhIPG9a8tLVZRwt5JHmaBEpepu1yKyIgeH9U6PV6bQBs2GD0Nh
Fmo6BJT0nEDrqv5u3j3qMWSwZZ6SqI+i3/zVdLUOVnH89Y0pB+gCnOQhCYaNPTrdGNZnu074lwkR
xf7iOi1shMlsVOq8mW3gbsspYrs7rA/n+aLrCuaKksQyVQ9YklFZLs6wgeweGBRaz3hKRh92Cawo
U7YRxQaLVbspoOSa/e1sQJ0t8GnB6z+yJwzCPVVYnXhT3gHm2KDAq6SaBxfq0+J5a8fQfIZDiSiG
p3pq6NLZVI0i8jI6muNRwIQs3RDaf3U4oMQ+cfWOvWtVNrjACnOEYudln3T06PFxZhHmX8P15NXK
6erUTP2oW/U/BeumpN5E0S34XXa6LzBbBPS95m0EdzP4s/BdX36DtO2cpb9wK68kxb9E/EDfFfr0
jALfZV0zgdTU5UUBy+TDvZ8OarWA131ex5bBNJOfFGQ5OqRNk6VPHxlOrF66BU9Qp934Nq3ECtI7
BqQyVmxJFA9TSttVOCLcz1sfZdHKrdUexFgQTjxWniiiij49yMwegg8VIa/hCk4vSx7uXjXbQG3L
9gsAut7n1nNRRlZyHKgC8oDLshg+nMpsRr8PSoxJ05gD9AQmvAqG8lC0s9rCCQImQ/i0yL1Nngpv
T57rAC3v/uHjLx/PoZ8eDqK6wSWoMH/VV7BWtBZUFUdVc57bXVNZ08UVbwZYKUwYvgcZrff7DY7t
4ImhFSXFq322eNBeClYKs5qJEcKZ/TmmmziWBo/asp9QdKs0z0J6mEFTPrwIPliLPLXaU79TOEkh
aQCPv7Q7oaWuY8l5SXpr1XNC0WKDMhpnZDZvEQ0eZsoPUaFNQ4Nne24mpEE4XIcELnPMTpVjMMFy
HthefOiqJG+gdNfh64sgvTaq7pBCcLVgrrE0VaAh+8QZ8/+Bu1RTIHBNmfSqRGBolmZOF3r7LndU
IBOwRoPpR0niUQ3qPQnVVCL5QxbWUZBVKKLOeCVrAa0I4um/6cfIpNAp11fDpsrY+VNnq+SJoLf4
hJ0+WY6v7/Lp/ekGOO4heJb56s7otfS+49Gfdb4WZGgMw8le9mTByX6UxpJhMSDnd1/wTAplfymU
ym/KXuP+wlsNqG9JS9TgqJVFOgI/2fyGRGc8/fLGY7MrqDPKhddNkcDcWkgjw0gxeQhq6+Wk0sEz
YfMUr8XHafulzzhU0YpGi+3GuZwSAQ1gGlQRzopQ3EYkXBiAeVHcW5zWkKYxvX31IClPhpXVPEPg
IO9kcwfWGU+t7axq9tc8H75VIqh138xhtZh0/OHasyR1Wz/GwDYYv2VAW4jjF9Az3hDfcC2AMNl8
0WyvHTTiCSXoHZagIhJSp/V81DG0HVLyuan+WBFztJtWXReKF4I9WmakjnfvUg9Pn602+Jmg3EVn
2qWxly1q/LZZnz4SxJlMA0knfzKTpFyNBmLaMmcwP/3gqJ6Gf9mewEq5oGX3a8GJx33NgMtGwBd/
T+1jdKGmnt3UT48eE8xIT1SqKkBv0dHNWRp/G698cqG10ElYt9sdNH+3zgUEmwTVE3Jd1TZD89H6
6Ci4DTWaP5MBjMZCRa8eZBQosZ6+JmlduKqa0so79SbIBBf9jIKxJ1+hNz/jHW7j3rWu+CpdM3j+
lvIdMZiRbpEkccsO5fVyTkL5szSfhF9D4sE4hJOWujH9sAVUk87OXwnccpCuLNiL6UHo76G9yCr5
hKyq9f0egi3TdJF6IoYSCRc3hyGXIUHvl+ZR18xwOOEj4fXb0j8jtkags5X/K5EHY/uMucMoMQRr
gBgoXtYfEOrwlW0qHaimlrn/9HwDqMsNfijOa4NqPqPSoRTsOwgdQd4HFD3oEDMl3c9Blnta9aao
RPLQCwxmVA3iVLMFSrKqn6rQySI5Q4IcQULmnch3Qoox8H8XnqobK9UyZru9oWU8rToJqkaY9NgS
DNVV/cHMV4N54/EKbWxn0poiXVGhx5hbBv2JPKacnayiHIq6iNtY/0Yz5TEnVzw9NSUMt3rB20IK
8BaOKSNOrVF3wMALbbyZD8YxT3rY2da+7GB2M5r7ZaDyq16clBZfaKW9Poioo32HCtloUhycQsAZ
8kwK9AeExeHmoWDpXD6tHIZXJ9xX43VF90YYxmm3naWDXE3ub70ZFGEc3n9r4ZCNinIHCLCn8VzF
MN8yHPCOFko8mqOcg9/AU+nExLluDS4CQPAujSst90uDTd184uTlSwn2keNZldeELhP5QiG4CU1a
+rxEwjji5ovmaGmZsWGZWrj2unczW9BkPty5Gr/WSqP3u0p3yVuBfv5E7/44k1MtOVzOws0Zh9Pb
1mVefP1ESajvjHFDkU92hzapDQqFKk3e5BczBsvJR5kL8V50Ho+gbe1fCT04YOZH+VLvMsmWDgsF
9owVxayrLmhRjAg1LSZk+BUv0pJmVZvH1FIgRiyRvOLC/JikMNmzFHSx0DQ7n1K5OhCx2eI8LEvH
FJrC7VMsXs17diZqbBLythGDmQEucuuwJENnn+X8rxXglkNUSYjNEk2DurUeT70WSZzkOELPxSfk
GPl3mod+hD/jiAb9MuFgoR+LZgW/0VXt/yusExVJ+3CMlLieB7NCLT6CzRaPEhgHAPiMZaq4Ry6b
DVtA6kziuCe3IMFcoZND88PgpkUgdK6nDGT2EKUW9ufTNkVsy+xDhVM0GO2H36sC/5tih2LXsxqj
90PU4+nRnWOA+LedbFiF03D5+qNMVWG3GM8qaJ9/9NQkUTxALW+Yiu2JcbESQ96KIFt86LQjkNxb
hZ8rI0/Ume5zUlLILgiRJucEQ4ey3Lr5S3hJkM4lb3nMb+UuafZUwhN6Y2yD52OswEfg2cnoR1fn
d+OVZF1eHHXsixQ2m3iZ/aYny32A7RJB07C1gRzmKgTlOpRMIzFM9ZVxSYcA/HqSLGRVHDX2M3fg
9T3P4fdbxyx1h+Sn9JJAO8DYXx42Z9eiv6VW5uQO+5Nkwm9OMTRmnS9TGB1orW1L/b0EhTXF5Sb9
5F7y1I1GktUv5+PZ6a4VYCvbKDcX/nWONN/fDxBIpiD0opdHGUe/yEW2hXMkCwZ/V3oW/QJ8HaMS
+cP3KdefR07qi1oAQThuu4oNN/mSUM9NKagVAuRA9yBTZjRORYEasZ9qgR8kXCL4W3WmJKFcZwFz
y+GpPQIrTjgqTF3aTKZ9HKPakBKFqEYJqFhxESJIJzQz0DhoyLY+KcS4csGfv5PxgnsNSJWOJJfn
uC8k7L7AXBgYZo2wzqBBm7JETMhqijuFbMXMJA3r8prd5aEKFNinBTwxmBCm9S6bzl47JzSegfRg
nKsexi6D9Hl7or18Wgg9pI+Ej/3JXjHhvA3INfFzmAqzRGSGXuUBsdyZmuHt8o0yFP8wghBhKb/n
XWpPA02aufxv7EXJVtZrVSuLtRxWTSEHSMtiY4Ewnnihlk2OOH7rQsdJgbOBhchVTzW+n9tvHzVm
fClNxY76tudBQROLbVgvtr6nRfFwoMab/v9TGkJyBq6SRasrwvstLzRU3CZQzPgASxzLo0CMHwPK
O9uL08fy8IYWjXv2cLirJMRpsMRFv4f3d8hBgqhLwx4p7ny2cdWar4JqJL+nCDosbLIgqCCb+qvO
RM9/fWXfj0rjw7PlEyLrLKybNgWY5OESTWdUFHj84M2rdb9VJaJ7o65fZEZ2n3IeJUGZ+GZy2EKV
Igh5VhRSSuc3G7jbc7I8pUePuI9JrTGvyePXO6YMyuwdxWoJteVwAfwVLqt/JZZLy0024NWxicpj
OeIMbONz6Uh54eWK62v3KnRKLajYC9iPf42eTjt7cGSuPtAAcBOecG6GgIvaaq0xynaXbEOgQFqp
9+3Yw1OJ0epsw0gujeStK2x5rv1XCapIFCvi5SQGOeHRYARKB61Ogo211h07RgR3Fhfq3LfTWaz+
OTadumpitKyMb/7hDNCY/+Uohyhwx+67L27VFmId8JcNzvCdo3DGQYVechoMpy3iiSt0+UF9Rw2r
YZZexQq5ofVsP8eOWuUbOBzbgHG1P+u3njro9T1SJffrs1oyES5/zFYZ6XngFWp5oZy44hKLzXa0
CNDfnU62lASD2x6Gksff+qyuvc+FoByBz9vl8YFtX+qThjvalQHcXCE3aBvU8A+Gc42t6ZJOuXN4
yacgY0pPuqAQ50LV45mZZZkSv+COnhHXcZY4T7KUF1BBjVMwKwG6zm3J70A/xrd/ImO4JlbbrdIf
F6oa1GHhyidxxcuVT8pinDFTtOX2IVIqjm2BbSI9YOS+eGLPlTb1pNtojwVcdzpTxMsZRxSAw1Pl
MoEY2GeToUl/saqp8Z7BVMv/0+BLblhvijxPHcQBOgWbVaL4FjLNiEIdc8Nzf1TnYFySCtOsUPZe
Nd700DDeh9Z8PDfbqGgquCjs6m8eGnb2KVq33gEDs0ibcRlGcps024u/EluR2PuFQU3GYEYKghAc
g3T1tXXV2HvXVF/ZHVXw2NaZFvJYUoHaLFCp4GGVvO9o0lQOZVxlWzQT3y979QQUaAR11Kg4UXTO
xWpk+IzOv3F2VxZBR981tjqJpjF22WetC937dttVwwrQNhm5ucf3Gt56pP4DK8uxFtlv0bJYm51j
fN7oKMojYPwmpyGB/rxVZPoWaoleEdfvLQAsq/QTVk6Nsbb6QlryRiaRo7LLBdJRluI0sXKcZ20N
Wl543cN3LEb78ATXVXLFpt0H60dR9yrpnC4y6b+LZMkdQBtAQNbdVRs2brrGo731ZbScC3zUPsrK
NmVYEv0/f18k5m/SCoUTEiNpy54DVtsAeAG5hgU3A0GEpFqACsb7OHvUrrBkYr2ZTnuaFNotSZPV
3TgChEfYZBUwRBEk8yQZrt/aGdESi/UjMurPHalg/EBF7CEH+VsSxEiwI8Prb2zmg/UlwGpzJqDa
0IB2aFLLDxJHrYvqNZCXSvWGt2yt4OI+He7BK4y6FhT+iCcvM5Nortf0AVEvJxIHuxrvSp4ZQrYS
jojqTiwh9c7A62/94qlegcMjL3J892F3zODW86Ukxubm3+QDiv5wgfCODJetzV893om1fcDPSDKi
ciRberlhwm7I8xPQFeZA0fvfpv6Xufsta8hMiDBmaXraLKUf5fkaN5MCAHFlSmHfSN85nY9ZHKQK
UbcgrXZVRUkw/s5rvqEZjetIqKEoQSbcHMpHYSG1wee2ovoI4i11TWeYSoo3VIHwHBdBGJTqOwsP
xwy069wj/6ljogfbqsExCUvhhf6WhCPkYn1B55sGxsSm2VXNtEuiwvgqpzw8LhzOj8o/7LNIuoVq
grHorqqRcufa+i1oIzI4LZEyCGZOK1yBMK7WDD4ICsLID+0O8CCKSDBw0maSwzLJoPE8u6t3zob6
O0T+8qeaGflYfFlykt70+OA4G0aKjpCZqIFaRuV/C7SmsWTOLjScnh+WqmzQbP0qcntDGx9fXk05
uOQMQachNtsWycQOWYXkW54jhaPlEW4uYBONK/77nIKALiWmMJ66zFWQXulrlQ7Dv8Hos1wV6TTY
EyEFhtqhxjxGOKc0AjmV3DksKQmERJPg79iYW95gBJ8uBT+6Spmf//oyVK8vQSAB5vL0CFH1vMz3
sLag1Jgp6kvVW45MiyZGHaZPneLvid6+kD+I9bDvk6ZPMyCZN0wqGu2hUua8B/x/ei4AFaq9ySPy
uB2Y475hQIHK1LMavj0xL1UKfedy0q3+hqEW6l4WR2W2EYR6jwcsmu9cTsfpBkRkjeXb7wTGh23I
3XLylRc2NCFfJRC3rA4flX0CHjnLI4vE04fLdG4QEHLXJc3ns+SZjzXBrlQX3BhtDI2BHppo6aL4
/LR2hhuPSdVkQp+4/MC3GH+wngkdBBlD5znr7uBlfmvla9mfTw8xdP9XDy0rXt0L17mvlEPaNjwV
SqIrONGVt0oQiiOzEx/G699d+4VPfd81aqr+7UDzhaokVx96lM+/pVlTYfgr0DBxmlOZcVPH8vo6
6omgl/5VCSnY8OqYu8tv6A0C8XKV1Qh89uPD1hXqvnWNRzkIC6S+GAHZGH4StzPjfZPiVzlrCS0g
kd+6V8Twh1K/tLCKpI/A7RLQipDftmX9y3xHaauLlz4boYY2ZBNCcWCq9IJwccwhexMcpA0DB5lE
0At0f9J1/B1TEyYC7dn2Nllg8xtNVKZ2w7IP8TKbdTIZ0maZ6ZfH+WHqy7Tyg5iHh4/oGwsPGlW5
Fko+qYqcFIap9MkgmHH5T6lc5j9AQZ80QrEl12U5Q6aCVXoKTb0Xr6TfQ7LNGukZvr+d70y+9NZH
iHAFqdzzLebZfH2a+J6a0OZBshBtEkeqpeRmoNXvoyhZHTjSnsA2QFlmtMM81ugkpXMWbiAHz2po
qrWKoy1NnxP7hDbax2+ZF5RHoGMsbDoeI5Ae1c5b5G4OVqmw0Cn7mv0I530U/rJaLch66MW3F1Xg
dxZ7plWwwBYIsjK2e/RVMR/F7eD0DQegUjiCNnwgdb5CXgL339JAeikdOBpZDZFno0Qz6AdrPOVG
LZL6WY01kM1dvqf6dfL4rtHztOeR18OwxG+3c91e3OWsAeayBFjOQyLWu/tdJLL2si54Qo8pyu11
e5iZdr5GlD9nwK+5qjdjZR9ZtMtuf1TwbkJbMoOR9DsRHtrshrs5fo9wCvO1ybI7awvSWtDDIoJP
3KyYyPo/Q+hn019kzoq0TslNW3RWhQNZ03cP3lim5MYsgc8u28T1FJGK1hppOTNreikZjVdXQRpJ
CMdHTMZEah3mlYRKmD+e1em/iT8U4vGwN9GosIOpMVgnLRwHbNF07M4+fplBapRgKzMcMBVFtU7G
DyflemuEilMWnZzasLFfbAWWYn3RYA8iALG9LC4aP1XJyjw41BPIHAwRloB58vt/zfr/i8rzk+6K
Ezt05d1OuCvn7nReCA7LSEW4sGlCRCbaNnbIflhJY08Z2HbVlaXT5HHSFhzpVSpcmP/YGHd4cZpL
Ak5sB4K/0S/7clFIRfbJMf0uWsazWTWaUfCUyJK+BBVuY4yQv9YQkbJ2fHho7vugtJscuk1D41vu
zq7oztQVwSIpK7DCh7RXYwh7Klq3erAFe/zkjB3ns3rETG+qHfxtKRbMyUY4tQaNSCn1nj4LN8iP
7WHgMEYBnMCKcbqzh+vhWXvnbz4Pt8o5E8lbUC+e//IT1lcZoKRYxrQaiOX4hr4IdpJWMZLk1db/
zJwi59KUiL6CuCVY9N7jcYfiCL1KRFRr5xTBkQpQ6sjqnGUzDFsRxDwr1vAvOPmyuTTRu1mtKOTR
fYSQ25N4oDF/ldo9Ew99SAz4IquzqiIdJxnVyYWNn57e1weHRmTYGUHLygCBZjELnxZRjuiUyOk4
djo9dSaClw89QDywTZmwZyxpEHRn/j2zS+htRR/MFUkI9SynIZjE1st1+FKx3vkZYc2zOctlt6jK
EWkdFTF9KqfF3MhpgKPHaVkJ+lK2ppKb0k7D+A1RQQR9/ivbrsvZMF8Bi+meT3IhiA6sjS63z3MZ
yaKtTldVt2tSQafbrQd+IP5ps4+eXKAG45hGV8mC0NQzqS1tK3GE0FrhTdAAYIEtw8a5YRjt+onl
FCvBFLnj6MDcFIAFLDoQa8IxtyVHpE930fN9TBIUzi3xUAqYtJ3xXgvHgYiHgaB5Uor5w/K3786V
NqM6Myd88yJXvYPO3e6H/AvFTJcUYQZgRKeXHTUey5S258ql5oBd+J8r4sxHiVfx7iBu77xyCJRW
/pd+eTkcJ5UQRXtV2NokZQS/A2sQR3LbKAjmZNYC4NAj0NuJajEgvxV+ymPN097H6czBMOZY7AsL
UvdZXen/4gAIrHRJGedL0mHfLtg5ZqUA5kLcvtvy99jf832Ije4PeuEYa3+XMzla+bCeqob6REhA
Q7DTJqA/9V70ayCwQVEwetLITsVwnae41uHs4WV6xDwouaceXNV9Bb3PFGkHywXPeQpVrhFCAp7G
PBfmZ5POMIunJOz4HLjYCfHV0QZfKzf9E3C7bZ+qmJ3QbemJ8B+RsYyL3gdeA/ABcLZksc9yjedx
A3oMWx2rzT/+iQ8lMtkwuUeHfcIFxTIwuUMYEQUNYj4T0in8UKj2uC9PCdVvjRl+fWkfym7gwWzF
58bwmCIm9l0JirgvjIbQfTSWIyG2Uu0LrRz1L+/lgfDXc67Mt1kgJXENHawmf2VMIuBZyBscIrqn
fx3FQ1f1GDvq6OKlSQ88xKjro+iBvzYGzdr7SJ9EVFCdySrK+0F9cZcQK7SdSf5fZiFE9hbXs793
tHVrJBPn2nntSBjQa3uUEXsZxnOtimuHYwjbWnBcKGQ1h1RGPC1Y8zPIp5wlwWjv8fZHu4oPGdtr
522SZTHkXkWYCmVrtgUCXfI6kTuC5Z6VNSaR2lkQQDqbAKGoeEqzm7BYdrdjQr2hwLCPtPzKuoe8
8JDwxgG8Ro2YPautUuClf7b5f0OFlFNwjHGSvG88W9U/VUuiuB2vLRxMO5oy0qkZA0ll11EJdiIK
rw1qWWHgBzEUQNkdTO3imEuZBSvExgFLqlN4+fxcRSnPmS+xCtEKCNtU8QtPGyUOEjcysPQN/ztP
3PgrdBY4vdiVCiwVhhy0DLix8iBPKDBWt7+3PcO8iVnpIeqMWdEAyyA04GzKOzRH1XxaN10jg9De
9EGACmjlAUInsRk5qabHSn4pvP/fIzuOs8Q0X3vhdyujUsDOs/ObrqokFjtkkFuJYL0Lud5xsopm
8gP0esR6+0tl3m30FPv1Wg0+CZLMljqPiwOaI8gSUa0S7RemyByhPCMvt2466lmiL3PUHyWVZ3i/
RUxMFSfE9g9GryvdSs8mumMWwkq4nkGKke9WynA0DplTnuyFOl7H+GE/eyIiZu1h8PTNewAXvLQ4
IuaTpQE+LfbQzt1RAwDryCC0MJ4LMHovT99BjvibY3iN7KWHdNGgyB9+toHkiiOXX/3PXUfbLz6Q
QVxBWN+RT7n6NsdbiSjbkoS+YbiUjKOwJz9Rq5FkgmWJ7S9Y8h4cBJiCd0Sny2vrkA8Undy6N8xu
DCv58fMdm9gImbuyhG/shETv5eSuRqvVXMStR8Py1YJ8lOUbMVh+sxoAEQksHnYxebwYk2aUT5nR
PAKvWTvnjCH+gIonDS1dqnpJmYReVz8D9n8K2wYn11x/LC9LPqzvbK0GHtLJQFgNql+LKLyoX5jy
giPu9H/RGiMPneqm/asBL9FmVmHRv8T7zpjL5XUzqGKvs7kjB4qc0DhPR5V/bpPDW1ywPYpS5z5b
v9JuPiB0coTOn4h2KC1XwDQJLo2pQ9SaGGZstn5kLyippR1vf9vBfbkhflRg1koD0BS2wTHjX/vT
pbH6/EBFrZqAZt0Zf+2z/ADLH2Fv08ih/XvP3M5nWdc+1moOivOV8VovyVZZP+7iG7HuRgnfROyd
ZLdEk3OWniz3xL1dAah45cqa47vIH4pwmXap9coS/lvJN9BRHQoifD0pVl9I0wh+lGAvb4Xw/Jeb
e1CqBa4wg1ghJXJOxRZBOIqII3O9cZhN3y8TqruIsHyDzV1xnp66kAYDvLMhi0+SJgXYZmbWiAgZ
nd7cS0SaRK0J6JcFHioLn5KAASsWg/MQo+vsaczY5+hNFZPdcUiVi2qQYnGNyxqzOEOCCrGPuw6g
L42tsEQaE0u5zRTmgr6cJIgOv34vwKDw5LCdbH4/IFr6f20+MiFnTUnmvynQHEMAK4YtK3E1NS8d
VA7w2ZhnnBTE8cp5gnzmhwLQc1kWbHgBle0SIbxGrG+tvTDkvuGwNgB8V3uUkcB7GQYMxa+l+E4T
EhAtveKrtDqLMVVI7qAhKKK8IsVG6aF7tszE1cwZyDuwldXfSPcsMGy3wjpAuxG4gNpK6cDnZJKH
MDwWkUM2OXuQs578tT3XJongQ9FZDkkhDfKAskHpdbdDzUdAm8myZhQEJsGX5pm2ntslU1P5fq55
ygrCsrhw19Z92OhaTF+py8Hf7BATxmuETvlSvJ0kt3A6qXuA86DaCupOLPLLnp1ymmyJ0gYpRCYG
NT9W+bwT4NyqyfMJGIFybK3QBwLCxBuAOod+g0UAIN9B8ZvssR33hjgsxtY/832uH8Ox0zkpb+5g
/Ql/HyjLsSzHh3hkSSjS+Ov4BwQu2v9zUSD1RSO1DRrmxVS+Y69xdXeHQq1TgagNXGZi2k5MBdbl
Nr89Dtd59hq1NkZVEzZX6Xtc4nGGnHY4GwPVY6pKDMjjcbBsy5MVod0LQlYr8PBHMjV2ymLQeZG8
v0ku+jyVA2671Vrlml1DsfSMHzwOkQ6ziRcyTa/n4GdNa2ZvRK9/VdIQYG5fLJLzLIOWWKF2oopO
6hpo6yLRXVTG8E92pWdMAJqYZ3QjbAH7+hfObPnwlmdTp7TFtw40smGtLScsLollfXMKsCdVjh9a
PwX2+FE4D3EAnj0XaMGJS5vR/7pmn43CYcCrRuxAyHW4xO+8jYGS+p1Wo3zKluebwh3NBbUQR6on
w7sptDpuTEAj+iy9fC7Zp3dXuCYdCGyQoaASX9vLI6a1AoxZ73xDzSPOrVEcf919smShed9DrSOj
FwaNV8aV84rw67URbE/MAmuy2+ubNOb8Qdealy2PJDa3z+wzj/wCcHBpr7dV0KVjh6GIUqZBKkca
79UmNBG34L7lvL/bRetCAdpce9ITzQ63vJt/0DfhVOknbkddLqmTSdfhb4MBEep9w7a/xl3JLx4Q
3E/tNngLLbow1wVQX+Q8SYCmgqnEmlyPocSH6WUYqW5aokILLbTEa6U6cu75S4jjy3VoHN/+K/k4
BnJMkrn85Ta8SZ/pglPi5jO9z37M/tEuNSU9+BnuGkcPPooPAtnqQwhTISs6m944Dtvb4EGaStJ2
vBTjy/RntT6rMSKBiXNtaIWoUWpP04yc56TiEjPBpUGAkG7jv+bW/PLmqJxLYXroL9yxYeP3EO4t
fW/7k+YKf0GJf+mctg7s5lGTClcraBUqAywzTO1AgHxKndyA1qzw8gbuPUCFS/eGh7Aky3B1kPxD
xciAlka0eumrD1lLyT+knqzLIsBBhT9EEjXGWNJCDq0bP+KoFlVlL83c5PeDuZfLSgaHNwLVInUw
/Spd9jOETCt4dUoxYjdz5aTovGzp2D9jYdeCdYI5T40x3lB/0U7ByZmDI+4UejZIMQ+6KjiwqSxl
lgcdYDmpsOoqn6putT8PCg79Ri13CKsGbxrROZnxjqqr/0+vL+5gDMT74j50emBuNBOoJ+4F47CC
ZgqM4thtmpP0KSxqE3gNCAzlTf7xgyyl/Kd6bEm0WhSrxmJerkIfg83sUkKvRRXQlU53KLeHnpqI
06/Brn9fAAqqBfjSIeU34pK4v6bJMiDE5lNZrAd6s5emZQUqHwtkqWzQbYlmiqjSR290oxbNYvS1
KeggLSN0B3ut+XRfA6ow57EFAvi9uPEYY2Byq9mgCz+3Thuh/rEHSOvsgvEPyK+uC8GqIg0oVsRT
dwiFbWw1TJcQP0pB4DvErdcBacYQqWhNogJWK163mntX45P2QwVK0cnIJG2ckeHpwrPnss0qInd0
ylxtoGD2UphDY/n3aDEkFS61fW/jwARN4lCu/jySR7NzpN1NHyiEH3K3ubCvNj/VFpGGADJb4Sx6
0GBGlC3QhFalghXtjDPW1FCZOCy0wyUgtP3I9d6jdkd7oNExNL8YTBbD6qBfEzsJ+uIlobN6CReK
Ym8y6AwMpAF8435PNmbkWMSwqUTJsfTJGJbOgA3rdRXz925DLMQ3IE2fmBilHuDoCoCQX+67ZZvK
+VSb8Tr6WhMC6tPlE+7ktQ0FcGWojt2GVy7BlvBnRJ/5o9BviRfPjnTBvp+IcGa4VdCjBmR17Evs
dp5TEsRC1TLvwkxA3ayA1dyGl9pGHfLKgEJIp8IbJoKuWSip1O/FdyX9hZ3ru3ZYRlfqznxbpj+7
utZVyzxkPdoqTdCVHI9lXtAz5/F+OaVcD0Q0K6PHhtHegtD8nEKN6EVHQW1upkPihdNmsJu7yD/r
MsMpwczF7b3ULFteG6jD++ESRou3CF6uaep7MC7NjHF924D5FVciOlgQ0L2FUh8x3HPagQ8uqhyo
YbNTT6IEC8cf6M6fYIgxodyz8ttGaCS0QMeWQSuxFv3Zc2a1xl2s/k9waNb6O48bjGKF62KjE9ua
+saITY0+GWdoqcafzqdwMjyTi/1Rv7MG/jhv1e3ujRBHTt00WQtzSaMa9V0ubeF+nEoMTCTBbkpr
Qs7yaEmu5bzXtbiUEGZLUW3Eytu/sjbGidddrXnhPOA4ZXX5u3ai6exaSPEQ/vqwlplQ2BYPQ/XF
iZOUv87MAISY5OEa6e/PQj7ssEGiTqjozA5BDgOiiyGwSzWni1jVxNFt4tauyybXcqLkxBufCeiR
bWrKtqBvvNtZoopOhotaG3tnCrPtdyOiGgstFLXklZSFNxScYKFI+WleDRxljfm4eHisNzu7DAW6
K7TdJ9Gtb8fL7auQEhvoUyhdhlhadGzay9xujv2PexSZfQgggScEHmHXFbnStnX9A0xFVvdnIept
pTBD5FVyjNVtmkD+e9iypAsxqNji0iD2leh8vUjQ0V7j+46/X2lVXX+lRLIIu97eXU0mTnSgGwy7
wDhARazEsFd7isvOu/rN5ddfUrp56cZkawjphoCuZcBvFYrQjxCrOklLVo+yoNcWsZCYw8HcEABW
qVC1JXNsC/8KcF6w+zHRuOTJQdSNlS5nzh2mTydW9KxXW+lswO84ncThBwsFUtDP7pBjDtkS+5S+
B5Kyg2LhzZml39HvHfMUZkaNgFv4Jq6H4nBZr9hhlJSwF6XQeGOgD31ICrCEycSiCztlB6N+bOII
VZDhZOq6jVCUvE0RVqohtYVj5PAnuJwm0uKg7KTvtBqp46nMA8yWPm1VqCktpyuud5d7pQUrOVFh
+mZg+EQGQLdmZAruDJHW70SPuZ0LlnQ2ooBoKlxx9Qc4PigVe2FuT1RJHhg6pXV652gaafYgE2eh
v64eaeYLLM0YlXCD4csPjFdIxAs5E2IH09Xv7QJu7qjprqEVN8qwzEyIUgvG/LVMz4VffnFN4ZpG
2mblR4RtLTzaTh0ReLL9bWSt72p7D9OneLhpIeJQOc+bJbM6Gg7tBd/z8gvO+aXVCl+KV0O52wtL
DUO/pdLtwoF4P/LjocXnguyUByq/X8WVMrFul+doiEJkW0cnqW76iYjaAQmzoPAmb+PB//GrMuxQ
OYiUEAUA3Eame6x6HM5KWs5XGJmv8KLQjy+zevEOPuyuguJZSOO+fNHmtZyoTpgEr3SZgfUfTymN
1+XQCmfc4u5haL3tAh6GGauPNDbuF+WXCjAhY3HTo9S8q0U09g/1EmDb2i8d+H5Ey5cB/UUJJ0jx
aWNoCUXMkiz9W6oPkC7ZPw949DBsd5Ppesgz7Vv7t7lZ1Riv/0QwovOHmqCnYNewWuuEJ2fdo86j
v6p5Jc9a5oYBR4AACM70Nw9oM9DCMpV9EjGL8hEuBoX429s+veZgDNtNmUJ7TgiQiwG+yel1aLfg
tJWtTPz8vnePvbevL5/PFqcGWMqOm8SHJcM6Y50dCscLG33jiNuyr0SM9aIXPKvK+h7uzqdt0Onk
lDTj6lfKHsVaq5dq+Q+8bcG0T1+kEGSeNhq2yson1CdKxtC4KBzY2fE10vY0b3fOY841IK4mTFnY
TroZdqv/nEjPySDWXsReSWDTStsAdlg3hx6UlGVN2d6NObFJsKdMKel6dpGHqK4kbbb8ZZYHlaem
Qs9JvCD93xeP6nfTu8MxCb5CwXCAzIO4DCl6vU2oG/YLZKtnH8y9oTO+Xk9TeW//QatrFuyWtDiP
sMa/0aFTZPQ2YSRLdPC+hHqyGLDOiNcWABULK99c6Yb8nT4BozgLJxVMi3MlW8CArqSkmax3CHEk
jNt3K/jbKD9nULqq1kDb8ThqEKw7PC5r+CcPVHdtzh+ieKOVcjUxchAZPImtM3zNmLlVpoEw3xaw
IJYVlrBEgK/0bGs0XShqzvpWxhupo3BzfT4AAIiuI/TB8y5d3ArwuZGjKEQUH1jxOP9lEYZHYeOO
NbUf3IHr6wUWs+tgXOlgZsjIJmVp8/PUC8XzhqLqMpNfjZULF3d2YvPWcFJIjo8AMIVffirMWS22
EYwlCQdMqCCMVd2hOoiVFDDLxDaQMr7U0mw6pljzYLfLmErts+QD5NdSkbOQK0OwO3rWqHJg6iYV
JJZRCEh3spdUZlf1fxUurJlgj127JRoTthUqR6LCmXB6GCnyGQu1G3mp60BgR2crF8EIxiP4gWR0
ivt9CW5NQrB1+oU47EbY6CIBvqZ4Pk818XGC706O/DVuq0sqGd41GTcoBaAN1VIi7o3UT1qQPNgM
KHFqlFaivexE09cYQYQO/SiDJnmnY72azx8kBH/DtikTH1MjIKDcZB0EuaeZySGoohjqlAWKmyVq
NhOPeLUDan89dkP56ZP8vPosM8On3zp3NJ9UKUj2AIfUcH1/90rhnfzWn06LOSjgEYTAORwk6Eeg
95iXOBmvG7WVgohux26XWiQsmV+5jqkEAPo+OtUSFZbTfOxriFB4XOOBIUo1l8lk7ESi5HuwvMX2
JiR+7nWANiGPPrrw65amO6TfTrLqbp3iyMPCJ3MuvmeCN/DAqoZrh4zwgj/tAGbY8ggjEwkgAiYP
r3AcQA4uDxarEUWRgwjZFN/Eahy6aT6KKUmVf++p7gDcthWMukuZKgB3EEpCs7xynqnSFSwCR7yv
786usjBVhTInovKOGk36RXV/q7X89KuKaIajUuyojDDvJP2j0j3Wh0PEe8+3wEHtfMfvmaBBkMYZ
h7E3FY1MRrGEx6NOOf8wFbKJCCCYTlJKBhVa197SeeS9FoEaedJvZ9VxzM02WmheVY0hDs/4Rcbd
E2lFRBECqKecUMoez/i2XUa88BQ1wTqCUr3rj7NPobAORelvEcYNxzAIaFgSPsvYpVGLI1z/ADja
D2To3Al5nMPNDOGSv13bdCufRbNV4pAb4LtenQxGyCCwTM16Pok9Slt+RiGRVWZFwfmB490IT1T+
g26+dXPlYRRLet1J0R0ECCR1TBFSvt1dZt0v5sL7g77lGke61z40qs5mwDmPG1fYtHTPgHekKP4/
8JmMi1ytUq4uvPPYBimNnofANzfH53A1bDQtIJsru3Kfi77/E99ExKl0L79HjfJZkT2PPEvV1QzH
y20YR1TzC79mwgAYdvqR9mdeItk5xL5WLArwfV2pXYA2Of7DIaYjNiG8nePS7gCEp3umG4l3byLC
qfdnSNf4kEPfg+9uB5LjXyGgE20eK91oddW8jE28bpIqb9hFBumPfjsfck+kanizgsIQtSXPaRPq
kR6WWkLrkY9/noieNz9YO1kZCqqa1Tfsm+ADkZo0r0phfrdAXDRThpg1XqSHzrVEvn5N2P8wQ6Ws
YNO5ALUYZ1ftx0KaZ/kOOjdALQtGnkk6wyL03eAQjhshSz2S2rG7oSk5KMGgMdcgrutck6N7XWHb
RRhrlkSSk5RakKn8ZGQwXnHbL9ydg0SIwAQnTYTTQTRiE/zMCsyOGCaVwniJ97HkW/KRr/wlDJkA
ZL+J3g7t1y2wAXXiqaDV+fTB7H9b+UABOPQUchOCiTeH75WXIVDVcVXaQCYlBJk4ZDk/pXGh+CNy
tPOgLqI1MNlhoB0fGhkmt6boANk9QNoKQ3sqAOJod5hy/yULhH5jgzx6zPHpzZ+lMsi/jvOP4Rzl
tlptfxW6GFWyj9Eb1455x5ofvlopp50fcjUR4nzyqVF8yUAg8LNLdjwMwFylkTNDCa1N33JkyQSb
ctB1aHeYbIog3nxtWc5MryQiL7JMWcnt3qkHbFtUhaERawHW9nETQga90sSR+g2XWmVe0byeKG3K
TSMz4aCYoB/nPUTDDZw6UIghcPvmHakBMyr7/g7qwrfFcYfOqWC2XN/xf2rG7lDh7b48Y/dzDKgL
dqyoPky0lXjIINfIf55UnMJTWxH5xK1vAb723AXExE4fznyiJeqGazdCtuq71jZdcFgmu+Qh0gR3
c2i2+Ox/IUkf6+BHK3etHCGtSGMaIPQGrWDyNq+TS6zSiWGd+1rWGiuiX3aw2nEYGgQWxaPi8635
SCKcNVSvLDdvIAv7IJ2mylrZ0BhJ2cBwAGECh2YFQSbFNqn+Ib4hN8bBVCxUEHkl9DqM33R7sHy2
RrgyjPdMxbU68T8tDqZYe3IUZxt2w4UIFjfvVDpQQz79FbIf8fNByuR/a6/R2x9E2i6cfGqHqw/m
5NLFTBlhsUJAZQmXsQJJ9GYG8v8ghj0MQAFvgiJd1d1rUv8kvMYXpSL6dLmcZ50jqhNqv5EPSIzy
nmco4l8kuztZmeOyYVpciFHzip+za+JkWm/nwRdfZW/jhvfojFagJinQrGrvvHi45hpvuWrcZU3U
FNjURP4sNIeGpp7kJbJeuSUSnNMiq46wX6rBekpnn5c8bpFCrD1L6ZbS9F8g+qv4ZkKBqgR+/VrP
McOKiYV/lCIzN9isoQxc2u1n2Xx8cQ+dMlF3/MVslVRt3x0w5XrWOUIwgjaSjHFWWFYSUpmvB0T1
9LhkuY3cRV0LNHbOJLiHTRoqqdeb2rgSLNU3ILDOq/ZBz8urYUUqBe0KtUzpZ4YQMXdu2Oh5f6Lt
300328NjDyJ0uxmSCwaiwocru3eHCtAF0lqblXpZtPUVbvn+YFGcS7mrMYTYoxD8QFxaYdyjA2aR
oV2+uzOr0lu1F/UhbVoqIUEe1mVDCLAoN273aAPjZlXrY7IPD0z0X6qvhBNy9q/1khpH3CjD/qKP
H9TZXksTl8AHwTKmC5E486wbFWlBYPVHG5TcqBgCSh2NhMwXDT4yE8xZkSFVMB5n+DDYRJ1HYQnb
niS5W64HbWSUPH2Xv/GGEuDTzZjIh+ZXXATm1EnFMLB8k0qopFfEVEvDAUvb70dTqTlAZAQpCRNU
tk082sCG4EqGyXgbvNLa+Fl8m/EnKmzBWZXX0vdGC9h1U/BrqlC56QX7EKTGz6sHPEIVsr40RILT
4OBiRImWPb2qWCd2V0dkv/wsTUnyHyHg6G9kI9hfgnqJOR9DtJZnRagOHTnrxASHUP7pU023Zgd7
okmgQTDe7DTtLRDGKCiadRq6nynrXt8VisQqO32zO0FpuCU3Co/Ref6a0CX6h+HrzYI7zWYZrbi3
/FcfjOnD91shEA9+53lRfUsRhENKF51G0quHtOtx3xhehXnFQnZefwrw4Q253GQUS25F/RzFAite
IMyu5b6NNBR7OPaqntzMPejhLA17q1LWaQr4zJFA2+mdQQjDAYm+0qZDO5tnHC0SO6LS5Fubh4oi
2Oc23W/81ozym2H/ykocYYSmhiqnUkI1VM5sxC1Y0xb5DUBW2WrI0hNyiZLFeMoJZMgtzaYgePZ8
9dpdtWvhwtIbkYWdQADcpzPupEXeat0Zxos/habKwWKiuYqvp2pBg7Xauy8lCRfrro4Luo8XUn74
SJgu34rIUKUkgjTH1o9FsPNss7Qqbg+LF2die9pPFKXgB9WKV4UiSW61ZLwEl54vZ23+x3peM3I1
Kxwdr/6GZ+LuDgc5iKmCysuvPtEV5FFc8q7V8W2bUgU0DNAyGlB8pwXACqcN9X8l0yLnzTT9b70w
fDLJzvQ5i5crF6DRk1fWKG6TVrEOUul5ht/PXZ3gt3LID/G7l24QnxInJ4KUUoD+s/yQA+O/qGiT
EZai5CFThgpGPKrJ7LCTSdlVYtlm1UYxjyh7tDz/jsb4bBTHLR1ERjB3w89Eil94owNvKyLxz5Aa
OaPAfA93AfV9tpBXPCOWQoA/Jm/8TeS60roA0++YYra/pZF41RG6yTI8IXaQEt+l69yhzkZ+83lU
ImTN4ank2IkhKSUm+pLwcEy1ahlMCOD6tn4rhTy239SvJX+Y4QFk05ffQ0IdmzRy5Y6Eosreat4s
Likg2Y2yCKkl9lCDHRdlvcni/IQA9f6AJ2Qu3cFGL9CP1wChejczcNP6JhN+C6/9YhCKlb0YvNto
zC3uZzauad1gnHEpw4InInTWB01LemY2i7A97xF7fpCLhKBLPzFYmno1ClLNXaTvHn9AcpRXylY9
3FF55kYX/WaTAAkujEsNLNxcbeRudaSqj05Ce2/C3JhnPJ3hX3PLJd8WHmcdWvHnjd2bH4vILTqS
qQU4/YuRCs/pv4HlJkxdjwmkvpVTXrFEaVTDYiiJCfX8ca4tnFpSCIR2IYyWoy+lKk2k1qwqnwb7
YykTPNCxLxa6er0b2FQD03RE7i1oJ/wlnlvkyuVsMOsJva0h15aps6d75NIbiMc4J7rMIIWoqWm+
dIoiy8qfftk9U50mD7fVboUs7Je8SuC53NtldY/lpOgDlRca2TB4/x7Rl6LXCD8RPipYAhhqMmjy
nBMEZ5cqTfTIOFGc04SMWiqlw06WPUKmfSMAOr/DFUFu8n0kt+4ZLyd1jwrqKBfn4ROfW5qcV53U
ZWo2578N8fOEeU46GlnE/2tjy6eMPm+MMBf42y1WxJzYLmn0ufBFE+SE3bCc81EH9Rz1SJKD2xFC
Vx6AZF46SUEgZ5GOwpTCcA9eAZJAQVww/Q4VS6yLF4b5iPw93bJSW0Gu5qjEocX0lxeBDY1JVJST
ixA79Ip3z+MUOF5+1VGH64ByYZArTUTuADr29pR4y9ZEUJMDjBp+SOAJlXSE6CBtjiMUPxCahWJq
3JGFsu9TPcXPJUoa4WwSrKwN0Q4GafRhPEjx6GsXI4ffv9bX2sg9YxqHETL/RKy0IUE4txc9D6GI
KOelFT/HasI4PcgrLrkWfnTD6qA9EprzwE3NZPoldGfvAPEkipeekNKZo7tnPLHZeLEqebxqh2pX
fdbIUBjcDiUXBw60+E3yvZoVQKxD3zY3z3wHgIelgRvD6L+fNZ7CSdMhEoqiAYuCpUgt81FCAfUh
EPTb1TfwfdyUyOLmfSc34ETnwwXf4qodWvHKNN42CnFVh2C0q+8+jhzM6K6ZCCvc7/LrLzKS+xNC
GXiMdDklPRiGeG5VJL+AoQ5uO1jeuyHZYEmxLoFCo6ekKa4nJWbW5ab3HevlpGJ/O9O//1CKwXKo
+F8Hzs3Buirl5yGzSl9d0PgMK8yfTLlZRfosfypAqHpR+vHKVvC7MKcVjlrHrgDvFQab+q9gntPq
IDzOvhdvvkvmvnu5jd0R5NrV3gAf1V3ijMWJlAFSnqkv7L/hkThZiC7eSEe7Uo1L8SjEWhzIDKv3
2ktGGY3UXvNddyad7dX6ZsUQ0Bqmk3VG8IZkTMtfQ99Z7+bpuqsuQeulZXL4+Lnlsd3GExUSsvXw
NQ70w+/ZPh/8na//mObHtGQu1mgnLJK/8O47Y9HzUcKDAdUfzDbKMqP8Hmr08B3/wew7zb8AtDaA
+TFCOVGjx/1EbIfSegRvQCW3Ncrtjq4ep0LHRV5DPNCntjaQ+dW6LXgzoMPepkn0ZDx6ApXkMxgu
pLBk4e4OIk5CmUJkABVpEKJLHGHgTyhG2KTPATbg0idd67P7nsQw8wNkX7K+vZEJX5oLBk81VdzA
hwSH5nL+akKzBKCl/VqgcN1oujRkYDrS2DGRLzj64hSTs8k9YqLo//t54Kcro10QYEibs3gVtWQF
lLlB7n2Bc2u97SkvErFV5zHnhk4dTfYsLITGFjNgPxkhUb3AqIxDd/vrBjgJZSDjLoGmdT5yOLDP
D6gbacQPoKqv4biaYiFAbVQtWtiZvO9jzyX2s5OfHbwzm3c2Vv8ZKFpW6ZxF6imWsVIMjYBxs/aD
+N+7m/dp0FlWDU7unk+3qrsbsXA+gX3WCqRlqz0YE9xZOHn7w4wAlYlueidaJeAdrQFxPLUZ7nu9
eAdIMfVaL638ZFDX3cBOehHStecPse3br4Yj5BIib1uPySLV9NWFqZTeA/oRJnNnaArslyEHeTdb
s1ErnOMTn62gBb37irfsgYqWDGzDHcnxstpvdvhNHDr2dQ9JMghXtJDYG7UtJbZuj21K1xkJRo+A
x0t5qJ8aTyLmiozHBdOJN4kVABWS/4bc5PSrAdbzoX8QAg9SIQEGmyTVEwxKr9gxcm/o7MzFAChZ
kL1QsyQTLblrV2UJAkRXggJbRGrgVXSsVRynKgHS5w1BD1030SpXm3QN0fA2tcqbnrYMWIjG4mdo
pogmI9250dQN65qjIOV+qSMDj1AqIC7aFjOp9TNK+RNFePRoriOWKOfZNJ/IRNfV3gQ6UxFI0G+p
Eg4H/J3LfSqBnTM/w/gir/OmTZOczc8mLdfJ5lpnwfLrMsTE/mr+13pQBkRp5R7xocw0qMS3Z1BO
2Ry+pwPfDlpLZNyslPUUnmPZHw4KlWvsda6//MD9xCVznOxbe4j9//fg0Ml20SxE+qZbrpQU4MXx
dScaWc1XiMlNQ3yFVrUtHGegV5kkox/zIbLR4zk0tx9p0wl/mJXP/7RW2MrSoNKLi8p2X73Zjn+C
xFo/9rwONBURu3iTZudzsSz0KEfjcKkG4ONi6e3ApglIIfLrngqRviyyo+0mf+ZGDZwxQ0qkPGkO
DsX6aeu1M/EWPuVcReikG6Ifr1sQkFvYhGgnat82cRPSX+POB8qmicq5kjKx7XD+CCcftUA1K1Ao
eBQYcojluCn4fmNv3uJSdnnJG9uluT8K2Q0AAPYOD3iRAdazkPVjUBdoa3iEMv6/vhYPeajSFN11
/v8bKF7qgkcDEgVdxzcpFzaKw931Ykr1Zp0nuPNcoANLT97wTxbWvPhq7R/qJeFQ8jrHaTCzn+SR
rlVFKVC/PyrLfkKedMLfekhcRV8Rq+2Na+4CRUiJH9z1wNh4RoEq+Eqixz4OqYvauadB4G3kgkTG
Q3GBn1ex+GfjzWSOgxf+yqz/+TngDgUEODkuD2WZV2d755QJbChcnk/bVpR7LqOL0sOT/wcyi+9B
UGvyp2zNx+kkBMNWt8vaI6JghHLA/qQ9gF1gS7xzVyYlyN129Pw/IEXKxSSmYQtTbSYTBIX+Xz9s
cU+24WKId8oJo7rKNFFFA98lr7Kags02lxuUkXAuavyVpeaIRqQ241/YbfUp5qlqsRFFHoJ5876W
WVSejXFWaHM7YzDyitYB3ap8U+qrTNFla1ygYwdWdcVFpQAkhpDLNPEnUAsRb8e8pD4G+79KD74F
Q/itLbqBZeUUjDY8F7IgN5SdBJ1JhvNUBpQPYFXj/tVQM7jPYUZ/kr6/XSAeS0XH2irOVKuR940j
WQlOLaprGS5x2cqODzl43eQWlhFhfQYnoFkNtPjfVcv5lj5hAy+fmzlAEn4DyUTztATpTckOLk5h
X3GonCo/5kuuNvhHpQ7Qu/M11R6ApvpT5LXUxV5iRIpLj7xkadj0gd3DOwvOJ4vKVHA/JENyudgB
cVzAV2D2dplMMxKUA93sPnGDPQ3SpleOsORwUslucE7fCUlcwqDlCCYRJlF6gPmBs7HmuIyDJbBD
hfU9B3NaehbutkT8KsKlUV6bzEff8HGwPkFBDbjXVLY2dl9TllHazxGI9VBsWxRoeMrRYog6zgnM
G28k90/T1LkqBEomD9zGXxMcspW3fBINX7vx51/c/eCh8vZSOhEKtsdOKBcFE5Ol0ZptSUqsCd63
zDuaHrGUPdBwXSYiuD49hRDkPW5BmpzIY4rfjEC6lG7OebbooPIOeqiNowk+/icvSA0vqu6s9bTC
fOMD+VageVK/H6Ody7MhD/twUHSPeQzuwifn4cv0YpvVMHlXLNaweEzh+fO9cdSk9oTJr7ZcB5fj
7ymcGNbRkyxVQU044zOqbInCKUJW+dkffHu81V2DyXYA76O8puSSTOdl7kEqGtrjV0aKhbY9srG8
jXjgz29vCyjP0oi+ukOPjngOpCfI6gf7dxvcV0h/dj831EfHcW1Lz9hVTeaADwsTVeBIq+SwP6Pe
fNAaVKv5OH2KJfvIuSgKEtr//WbrBVSfNAv510q9poJK6oQ3IcsTMwUozWSemcXCurKvDGATUizk
uG3DSzIT/q+oBjrUx5t4D0jBXVe9inHMlEZcCFY4J/x07xzGNqFhrQ7IBSmLcE9soc0rDmtcAUC1
pnnRl9kstmJqLLv8/z+jbqWZLN7wU8WQ1BlyKL5TwyMChKP+ggyJr0xxc7zU9KLbNi4Y8cGju5lZ
SPB+KDYAXvbzXFn8dhNL55v0Q/+mwn5B4R6hgCmu9m4OrhKoPpt/ibsGMDU1F5Bka0e08Mqwzxkd
IjrsihuyebQhXfILjrztbd5PZZ/zokbrTQbJiTmUDv1/pyvhzRMOlXLqUeDdq694dVovJxntNquK
Q7lmBHcc52WwSP8vwKjb9Vqzr2T8iCpea38LfEJskIv7x1sNoiIyYR5UzsN6QLbIOTUssU+OmCPA
rjQblsesJl0LXtmjx9ycSNUJ7BTS995bnLfMOLZN+ClGLzDxh3cL7mUTIxDd4fZ61DDisFwsqreC
oKIrPtutIc3bF1pv42pQxmXjbpMHEgJw+6BwCFgdl1z9vBK+t25buuS0ZGv5i76K7iuHlHJ25L/L
fjWAJoEdiAIVHEKjh13UntWSOjYdYQD2irPlxHTK1JASwTm4i/WjXtRYMzOS/qmyg6S1aj5s8q3K
hStnxBlZbsVtw4bwc0D4J5jmqKBXFtty6XlFT4COS53/8qyWDhsYLDHviPSIb9VSYY4+bfVeZLa2
rf3exct27NQFgESjLAV04ziAP7j/0ioMI9ejm60FHIvjLOjVTiW9ymrsdysNPZQVe1LDIWwadRoo
bAD1fPULviUZu2HAiGKsyASUcw8LcNWzJFKbZxPjnkDAArE0E04QGt8fQb/NAv0esvT/8nsfIf0y
B+soyeg0GxeEXWwlxXSZlZ2YhhZmtmbblXdZ1C2QAiyzwoGvGymz+MWXD1HBAkEAW+6bWEkNdF5P
alsYIkafwQSIlO9BftBiC2ebCFeIPoTUw27tM71qFMsqkBvrUpUVhNGwRP4+W8RaabiWKreDcylW
08z+zg+Ax0cb6+I50cfLyIFPrquWnTx1Z13nndf3eZXbgdpEoAbJmBOd4PjU2Qz53/SlEPF5g85T
JJgXbTEtfBvq3Zbg2MHgwRr/m9GzivrZAG752+2cnEeacvwAQ65nGTlE//OObuSjyTRU8k59ob9Z
ey1GECTY/b0O9fMXW2fyVrUwUElG7CvB1qH02pAAM93RocmP1EvUdJqXradC4xW+dPNREgofzFlr
Iouz3xw7v+gBrNIVHZlZoITf8V+5maGwCp+wTh3g56RHVsI5vcNjQjsRRitKjyvYq131SeHxr1cX
lYBLxF1Sd8UaVN9yo4xzihQ5GUGAbuXWE9JPTT87XzCaoEuXwMw171n2ckKUxV3t9nFt8aJoNjTx
ZhmJVfvIxCRs/ZVt/2lITIOTTelBUIknHxekbFAusYCGPoWrqMRGIprl385Yp8q4oYQEl404rhPh
0tJO/h8IualDKq1FHsIvmPdh42vCmueTB8siuQ2KburaK9pLcmSh6OYDXWGw/qS93bgIoYl4E3Ih
8ykU+Ntfjc/0Y1nOVRD3T3hxNqVEYnp96SrGrsVwYJ1FR7lF/SJGS6lpBTE8UCZA2cYhvCTD8ewK
3Coyfh1W7yJxc957CC7dQWON8C810KQanRF21cTuPo7lEHswaSsxi5cpTYgkIOZ5OFHTBfvUyOMU
4HML1ZJkfe39ePvxGbtWvM6Is/KsxL3pMmYpSW5J3jkQbQyUS/M6MJm70Nm8FTI1KJN4vLLvGEM0
Sqz9sNHjHlSV1entMIaeKqiQJpMNO9k1qJXMYvF7zKbDqmzEyOrEVWjdPzCtoFsdcXTAVSjK9PC3
psfswftLStu2wdE4oGZrFGQO2mHVmIu9Wa8mVa1nbOjHfiGLXmC6acEpvJmHUIiZ8UdVSU1VnjFj
FEmrYwVyQFSwCbAezDGCEeANpXA7OeK1CJEhnRFi5rMhMIzNoHGyA7/6KAuu6fq9wAuLA9ERAVpN
24EzBmVvS48tRk5HdF8U7JmTPQyw7Y+jd3S+dF1hjGJ/wFd9oO29vG41Kz8vWMfPhRDghVpp57mo
jZQPJlotp99QBYriEAwEBcPCS/slP+9tL28tPVolfCyMQSpAyW0kVtm5r3SuTBn6P0uGsEkbbB7b
ximXFK7vHHJ400RZkLMIE7/07q/dZKGxaVYPlr60j64qdhCsqO3WoezY9mHFzV04L/HVw8iEOfHb
+yH2XMBREwcg9L4qqr7nG9U3PEOB6nWOVHK2kjcH6Aye6himuBlr9ZSoOBUI8vi9gtyAuSrCpT2B
8Zg5sIvgmGKZJ/jQLMtA7R0f4OByWXs29DkRGqPUdikHtQqkB5B61w5s8d4T6sPQmI8nvb8YS0U1
a3tGiP5/RzCRBO2PgF7BIFeEY/NGu/wwoU5LHln3hG811xo0LUGe2UYfFIzlciwslcJ0dxjtwuXx
txWikQ8xbixC5QIAaaM26vaiybrnSeFbW28q3ZCYUqqyQyPhEcL4WdU4c/MpuZXIZ+IMffdEfhmp
2DKEOHkQzTSBAQOqGlIvZNyrOCOkghPcZ1WjUu86+jqqLtM3W0LmXQ/N+G8e6N15g6YfaawbBu7X
M5yza8BCcDMsSWYqMuk2fjTYgme2YFWISdK7WcfwXFyYQKy5EV79/0g7BJvLhLMPLWQfeO/zeZZO
8PeFuuvXrb9nM2gv5y+J7zjE/ll1HWb7T6k260j4LCwH1LTQeAoy9C9RgdmzNeuKxYvxBHsyCcJ5
B8BZd8CLmKOK3iiZwH+BgiKIOFbcO9IOZTD41H5obLT7NP9/8bVtp8JDvUbnLhZzIV6fciLUgOjR
HgOLTL1Lc2pTP3SlccMysowLB4ScN7ReECOaU4InFNJNZ2ws5/xm+m915sVHRQjLtQ4CDzJwRvg+
W7fKt6/tF++q9DJ8M676zlupqUAfR8xUziCNljXvmRBQ+ELfKASRMSGNRBLMn+Ke7IfFWcuyiDIj
U1Nj6b5sgHwjpW9WITONhX2eULv8k1UhAVhg/Pq1Neo9klxPDXJSRVaw20JyKR6+jwCDxQYtlmMC
SDc84bGGxZweRRtPNr5uXIeEafIUHqp7j93Nhvi1CicP9qOiYP5/IXP4PQcgEWfbBH9BWPItr8WL
Kh6oUxQwaVhZLIljOoBn9dJh4Z9B2Sg2vPxF35cDqhRNhKFD+oltBdGUQyBolGXWSOUDaBW+Q2v0
TdFEYSepi1jQlCdRiNMERLCZrbOBO9mSNENh19bE54G524ddiD3H0KDNpkcrLjEaQgMxpCREyOwb
s7IBJu4oQOfPvcx/+nmtRglNVJ+S1r8YwN83qDGZmRAYWo0Ivead2cyna1bt9tiN9eHiRLebNEOL
UAnUcW3DN+sqkcQEBX+YiS08mj8xSI2uw6MZygi9Vye3YxJNTpbu6Zp0zGWhk5vIFK7YGtEFk4C1
CYdeNg0fqLlgAwW6BCsgBLJh+Zd373ObfRIL8j7/q9/J+lzO4Kz1cf7fznxHe9mqkcSzAqUmvTJW
qPkLNl+hWXTXCr2GhwdeXbGiY3XETeSzzdv3+SrqHZ4YRCo3LZq5gqxCD0+kf/YKWIyt1mDVC0sW
bNDIZjtStE+XEIo1K9yZ+QeExZj78gY+FIMe5UPIw3Elv9jKdffxe1ia7aglAFSi6olHD+TQS5nm
0DRZJCALtF9sOelUtjI1r6dOkpjBwBNO5CEEz9a/qhTeDosnOLeylqNEE/2qqNass2NOJwFzxCcP
FD4NpjK4SLMsFqiJccrsxamuJxqov8Ce7OWmtjgycdyVgYGJMUgM8zwZizeVPp1PtdSNKacJqDwz
R8zVjZAuVkW7nlsywuWYQ+Za21GJqM3ItI63GpO/Pl+kxlLMWj4qj5UvVoOSlV2QnwIC3yAH511l
5m28A8+Q9dhNZrGs5V3hd13jLTo8C54Gtxx9/npeE+gUcA7q/D9FAHQd+f7bJB32OC4HkUiDK4AS
vcsE3LRS5azbQd1JnMh8NvkFUcKHMOStd3ct9BZno/BJxyNYglLXQIx8rSnjlcV9DWzEalB+RpI0
Gseh+ItR46GOSo+9NQjbzaLYOYoBNhuLB+liuDjH1LK2yzm0oN686VvWkPYvF9z+aIQCWAnpe+UR
NbXi90bmvQ+FzjUJwfYSkwofmBNqNRXKtwxNI8I617ooUd3qAI0BEq8Sa3kEuW2YSjSATUEpGDVY
x8sapab5uVxfjMrCWom9V93TP/4oYEpwLlufLtLP2nUYzStmCeOQjcbI6WXvh3oJUk58pn0BqSc7
9Cj2lvkajxPRFdaxHaDtLc+ACFZzYXMYlOInY8qf/P5HT6STvd7Nz0k7raPBehn5wGZg1fZpbfkF
h1zmzGai5pXIkdIQtkqJF7Z8uI/traMXU+Wh0qk0AibqmW0cHE+T2MDgca0Yekv78D4F0OFE4GJP
IqvFRDuiy0taaVzm5YO/o3KjHks5T/3J2hThDu+4NjJ8VgI2O3flTFQae0Geoia17IrxhQMPNcGd
+CftxNBKxLQ67h1BAgQNhR37KXmYj+nOr/wZYTqjiztLz+uJnXDdefUL0EzOr8/YxDLFawzQWmox
S4d73WAPbI6AmVuc4iQe0BX5N1Q8+unF2md6CztUHJHqm8AGZZ4fYdIQzCr0185dvDVdhr8ZtijJ
puqa05YCiRkbrvT05gVKTIeLemJXMkKcRbxQeYWE9+sXQAd9G9qF8NnHod5UPctTUdsq29edmIEd
g7x50c1o+IR/BqYjvdxOZXv92YoUsFWXRXp+gw6SXj2pn7noRoYDNlNQlRA0QJp8hEHdQKD+Lac0
hzwaG6x+pCBzk2ysWQ0OLtF/6jXXup1y02MRsZqVVUNU3UQzwESJWBQ9w/+fVM6tY6aF5PlkXQ0F
+SE31huTgh+A1j7yFcfUkeP3suvd2R3oHM1V/Uu8K1jwEdfHGFOH0a1NBAcNH5xuy4VWlLfc9Kqs
JoCGmN3a1u3vmwxIxEKRi3vjFXZOKM1yDqxt8QxH1LN8cibIpFuXwVg6SO5CHQ8jGaCc5xsuyqQe
dBhbhpv/L6u5rdYkPGky6Yb+1Swx+zzk4TR51NpNky8wYyjF/6l3qEQfKJ5WE6iVCz6+Zl4MFmLt
YHaQvFERV8FFEBoPVpMrmed860PLhlD5erZegJq/G65lnbE6WDxHl1J3YAcHT9+PbFQqaWnNPX4W
0kgWKRGEngMdhbu78B0L/LHy6ktessNhbXTkX0EDwCA0t2/CAGJXIqiAT7cTgt73+3AYJn+IIErU
k6MoZdkJKNHUexTWe/8V9rp8YSWgkct2LxausopGe984l22+ZHDizboLM6dZBNyF1KtO/nsJHYRV
niZa7GLHNHneNKm8jpwcWVxQEVEJAy0LJUddN8jZWmGdy6WJoCjpSZc9wrT8iHaBfjZbM6irQq9z
myGqzKMXATL3i3JktoBIlMIX8CFsNk5ntdlI/hkt5ewBrmcZMj8lIextfXUXELW+o31J9+mlxHMz
T+Dlpb2ho5wR/YdcRFImCVFFlf7Mx8HJvUh7ZfPCDGKh85VCTBFDcljz4hUlteXcpm7u/s4ibSLi
piZjWyQr5Vbj3HPD/XYjPC1p/U2Nq+7OhmdcXj1JEdI4KHbqP5K30QNdH476SE2GGdhHp1kdN9Ex
n2edU+Y7koxrWf3JKZojbnZwQmOyUxbXPgPtpj7JdS/RUmLWYwYvEJQxrGy0NSC/QnvgPtD0KKjc
ck5FVJuzyI5KLzLQWqGLXF3lHgZtYA7bCU5cfVdsHyh34dIvdlqm9uEJqM1lY+JRppInJf0pOpqL
TK9tM/Aev/2Hs7Ekl84dQpbAf2xuSodH/zHBZUZAEYa2T9KASLUYq3JTgllU0IOnOZ94FIN4MQJM
4qol5007qqz9YW3R26wQAQ6EWQHJePUGZnG8rnS4+oh45py923TtDlsmjG5TyFhh6ns+FPHfGsiO
jKLZLh1rv6WvNX7vDqAKfXhZFFCMdQc7ZzMc+iRedlbqYEbUY+dJuf8feLCGgp7w03j2sSSmxTaE
x/q+1jKX32R9GeAz7hXnt//sjsd5tnQlsxqyXDePWu1TD193RTEc4bLs8fBqGkeY39l8KeIszppw
dJBYpH3FDd18Ar9hT0PWuvA8JiJsSge8X84PG5laqe/D0KpnxNOyab+zi96nUL+pFxjJ3Q6j1Mh2
0o3kErVWL3bonrhgvG02ZUuUU+1SGOIkqcArgszEtegvQocPo0UZeB6luzgel0nUWjfog11Hm7QE
QwbMCgB6Rntf9E1dyvXznPc6xxmYtKKHGYoC2NnTjr8GMZbeVw65tMW9yBW8K7R5yxLqM/yWPsee
LHnBGn5FjssFmCOO9KPYD6WkVUIJpAjBADAoU6R53uswrN/txTv7OeQtPCt0xzKOp9pb6GkKhKvA
49iY3qgqKlQYwqLRUpDgQl+7BbfQPw1X7wpoHBMRe9w5le8+zGP2N93DZuidXCh5JmkHoE/XFzdd
ib3fiJdIYp/zU67j3VoFaQVqVBB3dnjxs2ruRC2nKjl0XLNMizqDcQEPHZ34olnzg1oEictxIfr7
YLa237YDFPlQKKeH9ZhyufZ9l6xKLzNVArXS+cj55BeA0gHCHYjTFUDPDZczx1XgtTXkTMXLLcOO
Vq6NaTkp9p0/PB01xTYBKt04POtLK/ITflZUBvbTtYNv9TeKgAlJ32FbGiQHQNsIP1oQvIgd56Io
GBGkgnRWrRKJPa3vzgpUji2BY42DgKt4/n/ebEWPnjOhpqfhBM9BgV2BrRkgjY6AxhRIDcSGB93X
+yNiwM+Kh6oBDs1OefdMUPYuuV4r6IxUuV47ovQhxjWVbzR1CMyNzgXaCtYb1yVNpg06xU1KbEc0
Zj03oEmsolKC4lLvWi7wq0tCleW7/aNu9lwD46qV/+g+q8UgolaaOXV2IUq7+QZYqHk4L+SFX6nJ
ynFZuQ/7xZAFrL2GDFpEkag0O97RV5OprOx2YneCV/rEG7zDfu4eiBam82g6hzwNBRWCkP0/NzVb
S0hITPsb76mOgA0TwqD9CvbO1ra/Q35PChqv7RC0TYTb4u6Zd2s7GG7z2yn0/cBiBPx8yzgLMd8o
UDzraDtY/30x2WfwSncefn0Fv/kUjjbV0QtEK0n+3ewg/huOyqJUyhupNEqxqzmTBHW+zVrrBzAd
93vvs/e9Zmv5gFI8ITL45wnd51yvTJErOQoXTp8AlYcxpV5WlRb+d+BNelGpazlR8wPOBq/dW5Q2
zja8zictuSBsE98U7Jy6FVegfUWZ34QeTgBuSZl2Pyg6UieJ2WJbv41fQLiwhPm9BYwnWHQb8/co
ULZjeR/9IMKN2RiW2i0LUCGAqtug8vEY1n1Sb/4DMPLbskZs4KTlA7ddbjuA9ByYOEi2jRJZQn5t
X4OHurJqu9Ko6MSyIc+I5ydQbhFpOnN6zYIowpG1loCbFkNdpALZVH8MXLFEX1T6SK3CsXbcD2HP
1l1naeRtNmggOmJ1a3s0xBMz5MmJ6tBrcWavIHBQxRtsiCrWCno8qsPw2rq5+HqJ4LcRXeno9Kqm
trfbh0r9jmH8ojTO7uQ1SwcgGSh68UJrcvzhfcMFQAY3g7mcboIOrX0nnE/tv6t8v9VQoGESnsXy
6uFjr/dvFtavja3+9jb9po3AwYWc6yaEOmSlaQcGk5uCgjcyfADVWIlcWqloaV27PTu9DYvhesFy
mr3VE1uHDbgQEVdLIiafAVTcXsOVb5gfmptJ1KsxaIPmdMOm0FIepCl1ziwL7tvVrDMzp8jO0Oyj
j6u76BQApxzaYREyAqJTvgNt4o5jlz1DhTwJc++5zfHs/h34H0PRvrh0R7+dlkABD1cjVZa8XLhO
dmcLrKTnZSRWr2J6V/DfYYBeixwNgpgrJobBaYDte8ZIeTWNxCxdDygCLQUMkfPnm4vT6TupORPk
5hHY9X0HrgDUu2WrgBB3ZNp5huEvIUppgQZ2eeJL6AfXbySCPtHzdEJLu1VR1gzsRrAQaypczHpc
01t9Y6tyYx6Mdxc1l+5z+Mm1ppzSp9rnSJLIxJ6VhkGQs8fdt34u8RqnUNXVMs59xEHIge5uuUrM
WayMy2qCjpjw2S1aaPkfTk/juq6jjRgB6iFtIgCPQUr4GpzvW3lZLufY+e799x8wQL4LOCjPjxoi
eiwmMRiJ+cQ5Nn3nx8qb0DOazBFAQRX2WTiXkIHt2aijg2v+GeQwiCsS+Al5un418NyQe4VYvGX2
z2wKRJHkN0+Rb06mxpdSH+ZdjicBFp3VPlnJyJ5FdKncLJTnTNhKh5SRKoLUpW4OvzDu4R0qDPdC
ygqiIiEOgueXP0c/nFXsPJli6eq5eZWU7jMr3Qv3ZJ40BoRp99A6U/XVx3WbSaZkO2EviBBa7NyY
phExNEXk1GuRoiSJ8nlnBbitGHD89AqThIfqGCoVbFUg6iNFxUcY020XuXXBiOQKYAj8zMgfZfVl
+F9f550cFTY5NWu33zq+JVA662A9Vs2UlwLxtKH6dynkoAKieCPRFgEA/nzeratXH2BV5NWyLqyc
vVR3u0fkhrRy7UFqcrJnUAITeVRKEgIBYoyjjkkWXUloShXCWgS6pllaJaqLUzyiMGaHaS0h5R/6
rAAwsv9baikvZbTDY499eA60vzODbQzxKXv+u7uvJryW1D46vJXlKOoPh88y1hBAnziCxowQvGbH
02dzN7kCcA33pqsG3zenZzqsLff5wGH3xg6lDxdnGy6a/nD0fxIz4OwduaizVwaQW184I5xJ1hpL
htMntXHb6+b+OFgky/VET4weKsefqz12ro4sS4pK1fdDiDPccI+sNamDcWeaP8OPU8GnZxiQhXFL
OF0/okbrKlq4O6xG5u+dNm/AiQh5/maZ1+Nt3+dTfLa3foApcgVa+4d0vu05jL9sHC+A90o1BT3N
Cfz8ZsL1yruSir9KtWU3TsDRXjs6Yv2auFDKb2WPDuHTiTRlu30odfxgn2sfdOIjN19FXR2WzRl4
pYgB0amAmZm1NXnoVk668evIS/+FwUfBHIAIHeGSgYxOCwFcqYdTOMKKeqfPDrSjRa3JCevoEoR1
xpqoWSEPK5iNJ1sMPBf6cBHclCQI1psC27mqqVAg17ohWoQujZV4ImatMAoyN+Tab39QoAHq4lzn
bdW3Xl37fgnBRts4IMiaTE0DJX0gGDCZp7cChd3s/nYXIa7RgyrA8GF7a7sPId06cLk1SXvd8lQp
OXT++J5DlWD2Je7TK1mVQC/RNPUsYBvdamcwT9XxTj1EUxYx4vMdlSelVitDvtGpBO6k6ySLHV1P
XTS8+yf0E1yfR5HEfxZ9859qBvexrgUpz+02Efkf3H/9iYCkICPq+Nj29Awo5pyBudOXST186gIk
dzizjQ7qBtiGMFQmQCjqQGRDaaqgs+l/GNAE5pMHWLy34KeOTEiMPYyoGlgX2z4kRD2aM7Tk75K4
Fd1O8udaSWepy7tyxkMDj/VjD8WXEJaYvI3K4YH4JQEoIaz6D4RUeHkUx5D95BJ0Nrs12VDhaX+U
nBIvH914vudi2NHDjCqG0+xI3cyTL6xgJe4fxW4mWtugRqyJE1KdYW8SmwKtX4y5hBtJ4lL4Swy0
t7UQoTYYHFHdPUI2DeY3cIHikFcm47dtPUu9d2KJEGITbMmptOuFD0W1zrTBBG2bCoAKxr9S0S2v
CCFU+9nXL8CsCjZIwj/jZOjl13RNie3oRVQ5WFXNgBncgQv3d3x46gdNsAyvhDZvBYbEpAMp3kO6
4k5YwuipyEXC78SvDaSlQkuZnZFSCBPGcBznor54pNKjkmS3snpMNnghnbefGbAMxThXGN967sxD
bz3Qh2shszGF5trmBhqqyqGxrKlsc2Rt0cPEKHxCW0Qmkw6XZ3YV0V+eZJ9aGYvmHCCFwaanEKj/
AcjQRUHxvyFfgggsy91Dby4l5LAKwBuqm+calPcp438LCyf6m1BCMEGQi2ubH7JE07Q90ce8ME8V
BBS99F9sagC6LtGmiygsyFFxZYkHiW52xgj1BxwW92doqYaZgcS233u7fdLoixfJ8115C461kao2
QnsqKeSe5YmZf57KVSu6EgPA+yj2B1FIVZNqYZ+YkCF+BhrCF8d5Y8DNQOxVD6iBM5Yw7dPrz2vA
NfTPWQg6avgfT0lCMrNWu4HSH6Zf9RRaeF2wyg9559+ruxiX+B7xATK7cLjRIkPTSO0z11xWml5b
v45iOgvR70DZl1bsDbQWVxatCIlUYNYF0Feyxb1dN7LZAw9tZ2nyq/T356x8IetUi9VLH8ayVbvW
4K8X2GdIwAajX9Nc67zLVt4To7pujozs4rLDGZQprC6b5EzM6VT6m9XHMKGewTi1DEePTSeDHDzB
q2jwZ7YNAf/jhOPCWBh1ZTWxNRIts++ABw2GiZZ9VgYni7IbAWJv1iGZknHaXQhs28gPkuAFVGzE
j3FJdfMp02jBIXk9Sq9/PZf2sZduuCpmcviE+WY0XbY1UA2FSUUrKInn6RCJBremwNd63P/qB26O
+xabdRCyg0EMUqMNQUVigTTCWoANAKsX9z5Nv4izoFLBPit/2oiO8JLEQjGwzA24sa8yLXyOfJqZ
6pA1X4E/8epnSeUN8OAz/OuPSpWAnsycpoGvNFelt8Wvzk8hgVc+HMRPDFmVWEBbXymnG0NBPV9G
hpVku+w1MUjz54TcphUGaQiK8KXIWePmeMT4IplmB3uS8fPRz4cgl+OMlWdDIV8HXIcxvb7LMzV3
qJrB1zQDLvGwke6Za3vZ5S1/Mp66tzsW9wE46lbbd1oUOxuDMjtfUaatxcegrF7pGiMZO6DZZ21b
QUjgxigwxwFZeqXoOhEXBZ32MlNR6lhtOGhJBk/J8Vc9VWqvRwO3z3GZJaj9zldHzWbAKe7C9Z0H
LW3nRlHbSC64TBAiZQ36L6xqdJUb8AFW0QIpnjzzJLkaLyIZr6q7vwDlp7PKxvsfMbv5Mjok0qXK
QmGsUEEV21JiurP1Yc6XPqL6eZdfz9+O3vu5Ish1rPB4xOpG24yJBUasgYmi6b1WFD6/DvHYhz7r
IXiU2ldXIFuIsj2/k+q9jz01se+/tZiG/btKHSnHBL5nuwpdYPYBy5KWNznmjeh8KkBLp63iF5V1
yzY8VaIkyFcqUNGnscEr0Q5DBb/eplhyAOJBLP++Xzn0GaqNkgjmEkdrUAESOmFlrxINneeg+3AZ
G75z+3vCsJgpLwIzYv7RHYxE/pf54LMFCvzMWWzyaMfo8FXOZpskYuxqN78z5byyyvcdEyf9Zru0
eTOkYMfBi0G3gXG1awNfiTkgxykWCZlNS2UWow/8F2e2N/+gfNUDh+mDdqF+u0zUHDJll5JUikdF
zbiNFXjtGepfziS+85+Po2l2VeVfAPy61PeZrESFAVB7EB/tBWhs4zWHXsa1hzH+uLl5Lv4OLExI
71EZuBAXGMe3gDie29+iR15tULv+chLndTTZTOVgReSrYSRSYGBfFLB8aLRrRS9YW3MqiqKbfAXf
29cQtYkCYnlUmcScoBkAYxyE3ecZXIJ3Muqlq3Hux0DAMR6AvxcVjCDh9EItL1aQKeeq5jxOJc7N
OdztzOoiFd6eFI+7xiZt24ydPSoboso0kMPTQimT1TspHnlkZRqDIc9biSa7DAjen2V8aWjKLDl7
/2ljsFkx4YNTqRvbzR34c6zHaVTxzFsNfKZ0PE2tftFxof+gzwJ/gCg/Wr6rtqpfMxJEedCN2Pq/
u6nVZoielFulzuPojHPAMgDdoGoKx8/HuvM+gYILtTbhGpTd7XuXYyM09t7+0F9dPIEQ2OukR4GK
YyAa0fNau1Whp8OM8y4/i//LMCCyBv2wmLok+1xfNZfPpB/vwQiM/G4c/yiL+4hPWN0nBtXsPGIY
u5cdq3saEw+Xy4WBO8UB2vi/vp0d7cgRMxyGpfa9y1IEyK+HsA9/QZoTN/ffdFJkQPF+Rf+UXvTf
bpka82kSBTod8S2XXjVWrb9S2j0Q+4nO0Muhb4mR3sVc7rjuwujJ/68GzLEQTn076ZvW8Fe2yKfi
qzFieS7GMnhzvl2RCZkZWppSrzAU8JqfSDQlctwb8bT8RHaca/Gbc5LiuppbwCMreRPBp6jsaR5U
HzWl0JwKVHhW4p9jgIzAq6vHleGGYvBqVzszjO+KX+ksDZzxr9XAQ+p+RdfKkW3oeNMsqmkbwC32
p+3khbfQydSu1fdfhFPdiBDTE7yQ4Az+9WIU8TxB74q9alymvkEnC11+6s1jHnuCWLnq6C2Cz+zX
rbD0h++IY2NboLBANRRAz/lYWbMCV4Yj1CLnpukRvdizq83FXxbXPA4RGL7fSk0mIDgNVgQmekDz
bGCKC1DUNjARWUf5ZurkVagiDrNeJY7auOoSy8Ebq2uBHkoSDDd1PKtOCSs3G5ifZzysgavgeHOV
etWqnzW0NL0uYt4K/cCg6QSOr1UDEeR7ZJPBHFnjPhpNHggExte0fLucrhAI3MuWDwKP2wMu/6aQ
MegJ0D9R+fEuHW4MCoTzkgp5g+tv+ST7uA3RlOTnpq0juOw7LQwznViapmj/xLn61XK02YO3kkJ4
te/6haSnhdI7+861sUn6xhieMJtK23zgnZqgW9MOW6sc2+LOQxztBjoUgiGvfdF5d3ymy/0qZT86
FkLSD2Vr4zC79vr8M9mksSAWHjz2bbxtYC0AiryZCq2xJago99gOJMd7WtpsGD9iD/Cf9pX40JTn
aaI3ffIEIs1qMIo+ZatYy+DtTbLKNR2uy4Ima+JAfB27iiFIsx+kZnW7aJBdJfdpUCAY23PD3kd+
pPuUkhcWwTSZdo7X6BybSqK68VNQJD4LCMA3xFhLzT3oL0P1SdxXZCHa9fIeV+7vPX/kbjVA0MKU
tg0ifHkskM7O/0Zz1Dk1goHvJbdjsH01j3KSqCCN4YTeagZCoMZ7K6QaJs0IFBAmXFL/ja2gSw+k
5jhH5jyqEcrg5NJ2c9hJnrP7YZYOEP+CZ7wjXx6w6na1m1euIiliNNUL4l2jJmFd5E9AnvIKDtdG
lmmt/5D6WbezWEqbDHsam3La8k7l4oCL2pAfI6z/GItU/vq/NbFZs1nq3kO/uJRN9oirUlp3CPkv
4+xcQ6bzjQoCU22iLlcBtWY8+z8gfO+hdsZcuZzqjHsPx3p7MnCCLVwk+NFZotF0VNzVcd2ajSSd
SMRVQW8xzgcInJFNaKMSGUlYtZvRnSxESHIzIhsKun0/BVdIVyRA/ck6lKR0za9i54I8Jh126zLY
bQe7dHcRLtecaxJpM8hIaZ0IkYc65/WiuKcPIyNlE4tQqjKMmosFLWO2culohi14djDhguCADTbD
6gL6vxZfFGSw+MFq1IpITIJ4H8J3+CgpDOGEugUxKi3l2AAMShuey5rsZzHI/BNNCsxcUDnkJDSe
/Tm9es/eyuBfz+dHrTpedi6dh+B/FvhU/sxi3Yy/mw9PsBZ1VsK98KldbmVf7CWkg7pkKyyIvoGX
h0t/bqeofobp9PomHQge7hw5m0hzZ1x+DhsFGzj3C+TLoj6q4H+v8V3HF8ew3DlkwTFTPKOc5jAS
lP2JUQtX4oGLVugDGMFXLoBhjvUKC82pcK5X9TBLkBOi2vQJU6BsrL16lK2+PbsmmEhEkPkMBwTH
nJvRB9pGDhX8TkcX+bLMlpzk6qHBdQ61iDQkNgcQ/sSWpKchhLcIiiXs0pp83FUH9AHR5dwf0riF
Pv+Dn2Q9LWzPJatflYNYcWa+nGgi1iYEipbqWpU2AMN+pqoaOtNJyXNZDepsLwibX90mu2AWzxme
zC71kJP5xRAMDuiz8oSI+OYJ90AgZH41Q0Bb0OX1DSTeSDnX1D9qcg06Kf/Uwxa1IQcePHiOjR7k
PUUpRNHl+/jSk23CGYLm+7Oo+7Zo+rXoSLvfx32XsHbloitVg0vPIiFUTqU4t76e/r10B+tZDrP2
vsWsVI+hNEz2FlDW+MEH99zDoYXIBYEuzVXM+0JbqhvMH14kWKCeIHbjv7Yla7mSF0N597+Yt3Bt
+yLqBrGxR0SzeqRUg80/Kwu+/ZiSm4Zo5ntOvkAyP4ikDHkqyhi5MdnaLisx/Qz6UPHvfdM8BL9b
gd/JGxsd7785zGjrkZF8umYJVHZ32mxvYIVAOCjtqDhCH7k1EXl7e19NM9hNgc/4iZhOesInAWBu
JDB2fFdvmpOFcShPJZjxM+7d5hJ72vEaViuL5QuWjQMR28wvWCuUnMGvaxZ/GEWfgIzoLNZT2acs
NnYXKMEoCuiJAVZimw7dZXgEuHBLXoWTzVWGlihgkvK5/Z/MeEme0Lf1PNiz0+1r9jRouDE/iyuj
Pz8f2xysBEO98I/J1jc9jf/sHIDlAymUNO4thMokthT/x9qqultwoP4jT634nZAFNl9BGLhrobjG
xRrlbnzCdp8d302NhWqzSHc5cDhaKVt5DU2p26fbwe5b4MNUXRd1Yz8pjl5hA2Qv4RuqJuvuU9qx
lKVZnjTyTfr3JLQBSSE3NnyAizCHOmP13m4ZJ4pFghUvImeRnCGC1D7LLIDUMfhtnC1yt3djFTLT
kQzkHPLfIFiXh6BrbtYwkbMVrgBl6m7ndDvYOYLSLPHD5m35ToeT7bHfzDJEDLLnvGEQ5/NpMYFd
sKbAdM89rWerrPekZbl18XvyeWnerzL7/pLrBN+KVhd6dJbnmZH4T4FUGOgBh5bkrCgf59MsN/ob
ky0Reg33b7ELOgIPYJLWCh1I0n2p9a9LDhB/A7XpoMN7R92hLKC79tJby4MHZRbpNxOfHHsSFzNf
Th/paORBSo6sJBFqdltFbqVPrHznbAxc0Gr1310tBuzcTmoi6lnLP0soI+jDbSLhUNMdnN1uj746
MX08G4wV8LOc9cEGRE2XzZNX7TvBZvPbi1dsQ2D0m7Sq+6Vw4GL/0OsKg6klV8maz/8pUmhH8xRw
umKeHaEDdadMoT7rCU5CduUd+JFS5zO0d24hTqtcBfwWvWQYw8EuYPi/0BsVN8oBM+r0zwbYwBCU
hjsV6hcULj4gx6pvbxLxjhpZ7BAmZx31stLcPNZFVM+3MWEUrjBnbcWDAqbDfOg6Z9nz/zaXq3W8
7B1pYOqVDmJN62+Pqoc1gaB0v0jUCvhBuWJY+dfBNoRZOTLUd374BITt84Of0abbA8SEQQVzV4pC
6acz3oaOX4npOKb6DAgtsrRkb1OuyAYKc6s1VHVTxqLVlSN/dyXx5XuMuS7rW6UJojb/Ikf3IF/r
dqfn1ievhEXwdbCjKfPMYeIOZ2IOyEmURUl5Vz5gbCVjNZvEAd4t/XzGn9pqi3pNuvquRS7pTie+
nWjk6PTux7GjBsnMCpl5SF0pueAmgRpAFX2nZ9ysFr6+pCQBIm9fwhimOtYUm0v4evRtFUOnXh0n
bS8xz2glQjsxHQDMkCtcMwRGLgipOkr6x/WYrgt6OzlMRXkGqzqHAGktVkXvtrR4LbA8bfUskFoU
lCLHUw3EY7LDeNKv+3jA+epcLjJpNHyYpw6hQ+jbXD64XFE8t6WkKIhogv7K591BvhVkngbzHBI5
xD64VBXn32sm6+Ey11j0J1F3BygxyGzuoPX6NNWaefx6CaW1y+EXY1Ef76VM0ZwI2Ih/HBUJpv7l
fIHzVUbjITNzBXeSUxpQ5+r7QbYlgXwxb5nrttPgwCb6xkWjD/Sr6gLecFOUCvkPqoZhGtmrQjzZ
96CzvXP+rDm/GzGERPYCbr03crl8718jsj4UybePx/xzeWNN9nBaFJwZDrMQotf4zuMTlA0ETJAf
j2eFhYQYGS53EG5nhNKE33/F86Id44+Nr+wBIOpvhId28Oa+qq8kcS0am/zURbMoKL/o+PjNzmu8
Evb/Xsa/das2gJTwJcwRhQILqrQSay10utmlrPLd2FLK19Pwy78ZzPP0vlmru9nPTfNY8Wuw4j0T
9TvmnkkI2+m0bUfTkHUemSMS1eUinBstCU52ilgCZA5IdfIEffSWHA5jNY8jQBLIO6JoB+nA5Ft5
tLQpbpmKAzcfYV8mSWF+v/kzzAx72d2LJ1fQFIxW67Aafwrugg/CF2Y5D+pysXYxNGUSBMX/wgi5
vh8UI02ljAYIMUjLTfej1hGTMyGFi3IbSTsNIV0q2VM+rqnSCcO/OPxQanolhICLDIpayR4LPtQ0
mDEVTe2uGFP7mwj8EIGmZJ98l8peSXaAselmk4hQBTEJBObc2H+KUNi+Ui/T6EoGh7yHUqE/lH15
iqdm1cSHCuCdKu5QtRjm0CnDdR8B1S3Bvd4U7ELCORfHeY3FHef+EIdcTuQob1TJO8mZ3aw9xY7c
grdHL6D0FMal2GmReXORm4dhgL47dwalaA2Hn/J/imgzir/YyTXObSo0hGNLwrUUkkGF1mhZjGRA
gUvwFRzBCG5D/6yhRc5VYcKEnFN9KWhferlKWFEuf0uabKHwjUWtJRdOajKieVESe7zb56W7qfgO
pjQ/pz+liy1V61hzOy8i/jOR9u4U7rQ01KstTEaU/I/NTkNhsw2Jg75lTSZtN4Cx45uBQi+1SEXf
IwvmLNhHJM0s+ahXOxvkC3Z3kNebwu6qpYfWvSpZ0kAxdcU/tDd57z9vOkG0x58rizpT6wwhnurZ
mSdU7/p6DVvDU8pNRD+5q7BLRim46I4RBiWeEgQCR7wpbX1sXBw9uuQt/ZlvhnJFG6/cWsTqC16i
l5qqoU7Sp4SpPZXRQk/4UarugLlJlRL8u5K8mSc4qZ+oUbNh0Lp+gREED+sqoThlCPro9Q3AvfjO
b/ot2lSvEQMUBKqzFxxunuGBX048JpIjAxDDlGdk5fPlUtk2s9NtQoTjynEY/MEnTCrLCGdpR18m
a4slrDxfCXCflchg0McVqKBX9zfMAu/R/4AOh8raIkp07cp5q93TWIVfCPPXbxwNDRFMCDA8OfFs
ArfjMVZxRlGujn97PvzI+DPqmWg93K1CJhZtRPLpIs8CtLkcuRcLWQv05ykioVMtUS7YODcwBlaR
WB6XzTSHyuCDFkZskCpI16j44iSz7HyuOkcySWq3C6d6IY2sW63SqOML96CD0VCuFdccfsmlZTEq
DH7a9DVW1AxWTaIWc2/jefmVzj1nSrPutUIaV1+jS1nmeJEVUYdVUmyKt7Ouc2ruZhTMaxQBiI42
NRsIpOZ0Vi7tA9pRrhciczzfwqkLtJwx7PhTjUg8DAJxcJR4gVXemIcBkrh1/6LAPuQhbSwjPFES
+pIdFIRJOUuTYAZTAhwm6QXtBYuV4XsDBM89+839HG29XY33BzoaOCUWrXjLY9QqBu/5RT6uTakb
4gxf/3o5pNBuQxuJM880O6eiD+bziK4NbAsbXOVaUvJQnvo2M00rJnMfiqzcUDEeoLCat/DzmLI1
odLGQI5k8YklcdtxKmW6oGzbA942cOsSuV13fOdtCiWzIAId2xPzFUshJqJfjxBDnrUshGPOCebE
fYjY0MzrcGGaG9OcuGi8KFd1mkU7McmwfphV90ocUzTI0cW0nRYUQBaY9L0thlwdAdSW8sufClmM
QUBIyQgf37FEaL9O9GneangYChSmjT2bF8hX/big4DiQAkwP4gnsJOyGy+aHX4kIbMdFwFHwe/UU
1msfxDHYdofBoQfrCc7HEQskg0uPetDzw36cbU9Hqo6eZc3K5+6zuPwFHHDIGcaI42NgZYQH0wYu
5yHOHUd6zj8mwUeGewDCz4jibae+KSaJJ5NHNbOL0VD5t+zjIkx22uaj32ZgJMjgEqC5KTlj467G
H8YmV5ruG0SL6EOQ3r6fphc3VlJyPymmjObIFQAboNr4w8Fb3nst9yRyrGKgy4d/zW/QW+bbaTAT
3BjUqSpLq0x9q2eFG1asD37MFAASh3TA0t4snU8fxAXJzunVapOrQpiAeu9Q+sOurEdF9utAYSQn
8VIGEavvPV2LJTa9vZfEv8dyLefBNfxldwuKCmNBrBH1yY2ocsetsW9iLJpHpGtofuB7y/wyyot7
xzPc1lsZn+WrjFojOoUGFpGYc7ANjjbBWyPcOQrb+XV/MuFIaPFMasCBT3Ja2xt1ih1DguRzT2xZ
79iZ/ZfNtLmjjVMQEXiuIlTTfVY8+aI7RHjfQlaIYKQ0EGiaiNRx4g5ZjHaMKvUoUEjNHhKdRQ8p
AdvIdBMjzFS2PkdNguJq9nbGzokRuBzKm7HgUCmm5IrtpcUTck6zNh/BlOLtjtcn3nxD6y7BqeYM
cHyGH9VOPt1l/2LU4sAtdW0dIQd72VoMAruipwmO2nVdevRYO1op154dlyQYSmYuY/cDQGpdytYa
PzmiKNvChCrI8WbIQIfj7VuzRQhnAxGorCfEnSlZEfp9XmBlP5icQoWhDAQzNFalAnt8/llf56cX
2ao/BTh6d4S+PwBeAb58S/qrjMjXTynCulxGGKJQkedV3HMATpQmrn5wFZbG7tXHMzWSaVTV0lHG
UTR8rMACxvouEFH5RAia3bTtP2J7rSBcIGKaswxJXT38rBwKx4SPu+m2ej9Wecii1s/sm+nIYJaq
lydTLjhnv/f7hVvz566VH81eFWOvVwMzc71vKe4vnkncxirZKXY+Mqlp73vka9C12+EtuUKrxajh
NMF73v18y2sfE2D5aRSi6vKvfIvxnalTD+N91DQzGKrTUeS4H4VwXZlM6CzrOGX9cqE3rzPmt873
Hsp846qUvdY5LeHeZI5okcgfScqKG3Rh65FcG7fIfyjAJNaTVT4yUKGU7UFk/xp/I0vgN+njUlkc
2B7vlo3LgV5UG6arS/l+YGGTe++zzHDJZZxzlvw8o65wZbkC5n5AmEmcxFyjCNaVkGfntBnxY8fY
sZ7JzYbGg5cknvn4WSEOJmjDauTeawsedzugZAA6PJs8xPav7drX7bEexQYAMmA2zLJjW2HPJKVl
W1Dsso7kXSzbU9ZhzrW11WDLNOhn93GaigR5OTHreTyl6MlO1T24e3ih2eNu8vbGACogmAoQIBg6
DsP2NPpxm8CQ554kr6h6HQJbptYYTMXHp0ZXiHA8XDxeHfOyNtDkaMDTzxGXazKwYdQ2JHOfAD3U
hzAvnuuzjiIdBGUqedbfNniJ6au6ZG4YQSKyEjQvfqVVvQd0EngyXHrs9T8+FqHiPW7F2/rrWiOL
gk6/LD3TfcKbv6KA3ePjM46QPG9PLjWK9Pf/K325UCGbLCUxZWzZxcpwZh52bkZueqdA4ABeZ+2r
MhjiP2sMyB/XZXfMOdatLY5vGq+NupoeM1zaLxjW1L/W68274jjvOEwpeMVo1WVzNuUQ72lk+6tU
BUSnmOp7MNqehJlany/hV3r57IsFUfLbdaM0kT1P4MixyK2N4DWavrO3xXKBsFKfvVlUvkTJ6Vgu
7SWFPN4XazqiOjQB5razx4i132N9WfIQdI6z5+8Zwb7aN9b/1+JeCJm2F2Hu2PnJAJ5XijTr6lMk
21rXwI+nPzML0W9R26WyCFcnVuIGk0LJ4NsDlav6C+pFL9mQNEM8manw0wQ1LYNHYrg+5yQehuAM
zh4tKckLokN380wpONCGI6i6IhNas7ohTwE3VHXIpVZhIbyS5FsR74cuZZ2Ufccs+byq9TINIr/p
mnG681/EqsOxTS+Hv/tOUAi4f2WlN8cbRTzfDg3hHsQonRF7Jcrlm75yA2u4+2Ozz3jipScZYql0
u3LQm5rWoZlwjauNj2HHeuP9T7gnKdlIS4ufRPn8p3pFL03BxbI+Rnj3tkU+RLExchvkQKrpquIM
nwLFBlB+AMKvk1FT9+zJ5s1yY81FuYmzjM0/pwc9aDracfAPA21Ov+MHPvM/tmW/92e5jpyjw8Co
CBOaxJWf6vmJt9+je4RsOydMYsy6dzLbfXtqQ3JB2sAGqU9dJfAicXFXAjo9rAE9qpDAL+FCFh+o
uMIibMOU+aVmL6iWVxbWGYm22DWoXO92dAbfyGnz2XkqFCVdeho5pOMpY+hqjz7tZplKyhx6pDNX
3EoBINpNvzwDmCo7zOh4Cce5hivjHuYRw66mYqYA+G3OpQ8w7FdmlxemijnauzJYuDgrP2yC0mDY
rpJBbpV3/yJSnjwUhzX5b0tolj4yfCiEei7ZbgDvm1/nm9zqwADFwNeL79xBYrJMeIv6IbRJp7WY
POx9k36lbBYPWjU3ODnQAQXURHdXG6K44pSnlzbiZ0DKXg/9LSMI5cB+DNI0Or+swDZyq9BRKB8F
qscruokV9/ifzfMCKC3rPXVAwi9yRCY4GxeXpXkR6ZJmsIbDaqZXmlhoUKoalNpJ5DpZUcwVkV7c
vvaqnXKvWrtVFsvv7BxYoXvw0R/TyXFQqD9k+gihGS033tPnsn/j0pIx0S7LC8FIR8RFesv1n8Ld
LINCKjE53bw1Pht/hrvy3ghAdkHYLYzRWl9z8mx5URMR8E0cs23Pb8l5+fa4phl020cotZ3TlCTk
GMsQNdqXT1yz3PDGLgKZ2Dq9PyO6uiiT1555Np9xR+IJ5ptkcwUAvrm2lBcpEl5vTdoPgggGASDU
f3OVNvFeLzCQENRCbFmwgLX8Hi0TcOu71jDdyP8AgIm9HnkxkeAEe8ylpIDcZmyrUGutaQM/fejt
bTtzzYWN9UUA0Z8M1pIvu7JCIfZ2AW+s/EtI6fS/XSfJGInh4sJqoUtNI/ymXy8qdOb9VD9OZ0iw
LvsO/RwZAImYfU9K4ff9wOnpMtD4tCW6UMQifX1PHti1oV3oe9VXHrvEm+B+kYaUQkSEYpdJJ73b
yAL0iI7+ioYUWVkBxNfMqTdU3FGZfn2JpFQqEY0uqrduWVIIoO32Z1e21YA5TePLpDrRYrObw3RI
6PVLKGB/XKxhkO3TMrqxzPwKYC2F3jvY4Pu8plfkkmbwvL645Ta3z2EbimHmIebfSusaYiZ+Hwxl
QotCyNCvnX1YWMP0W5Sx3WmNhmjTvpvlMtXOkawhmiyUf5FZni9cbxgJ2S9DLBoQcexwshYiPr/E
BLHVQlNY8kMpLE+mJX/p0YhWbRd8OdChCqxglwxdyXOPxmehp/9y0xKDCMFZL5TX07IrnO3AgYup
Gfy/FsNksVqL7Pcu+v5rn+Ynb3dGWdFZj+woKSbk/pBg1lQ/lLQ3zYH1QlwHCuZzkIEdGrtrt+Nh
yqqP//J0SzQJFcACOgPeM+gQPN4b4F6C0we4eFdM8anBqyPFwm8XrXtzux6H6/fuEwQaD5Tkb7vU
6/ziVqjuD1orMWncGklS7HLClzaXV1mt8a7pErBMRve2Y6x2jKu+PfOb76r9o2Oj4nyznnPdxebv
G02fD/w/M4CbSlich+oYi0BKGwNtl3gEr3a6GKVjVmR7tB393cySAhA8ug4Vk97vk/aWBUy4OmWP
WjHFu64IfH94z46/CidvSPVSrygJPGteOrgPdsyxKyvyjPqQWHiFzwfWBaHuOpkqaaCY10nJQ8hi
HKE4K1VtudHQVLi0XgeQMSJM1jo4xFjbGj9xNkrTSX4sQ3ICx6kJJrBhj8MZkxo37HoV/4z2Gzko
9WOu8rDz1EF+Qddbv4+2FkuaEjLn5O6ypICssZpNxpsTavc13pARipR+b4qUr01r9hNRmS7aBcGk
wvE3oEncsNhCPWFVyShRjK5ddOux+i5wn8Iu6msLr5JjUZPhPMgeB2rOxyUdyw1xDSCUG8nGF69Z
CmmBHXWDIVJ8rnzfTbmicNigzVuTzPVKoeLzq66n+wui/NtV+9rMvJeH0u8aUJ0ykjSdokhSvHPQ
lrXSzqgfWHRYcZwca/pTD3/GxZlOOK2OiA2nUmtMztYDHu2lsMMG7mr2OtHNz0B4gvWMFD+OoAgB
7pEe+/4MFG0o+YOMSI3HfxsmpDZXlJc2oQsgktvQlbJHpxfM+0hSCgCfpdoipWRK+4tVNka4lzK1
obtQtLiZMlOdHIoPwXf+6m5trCMHuzMn2j2XWlrc8Y33VZaoU3TeJX3UPBZzSgeTOFrrXLQ8YbDx
YF0kC8w9GgHD6tfvy8R2IrfqA1yTuu6kM4byJuDjII+4l5Q6OVQsCMeiO1J6Gj4e8XDuJqTSC+Qa
RXekD1Bk+16Dg3+vIdlMD+1njkmjlsuu6oPPQe7C3PsXJOyklodtJryGDuocabyiJA7ZQpdVVFOf
+LXIm5u5OHbaMgJE03QQtUJvLSU1FUr0isODS2nl2DLi4jE7S8+CkvuQ2V3WC3vp2wZout++Z75S
a3k9E5YLsM2m4eqmIvX9kG8oc7skSXRnYmLoNNgqO/3HS0EPN7cu5HnnnA+TdlI/X5qtEwrfL0zH
y7nNeDeQxYP3P9ktdFx4b61nAEVx4KIcNLS77ddvexbmfI5iTfiaZ8xKKQgfuhN05MWgWkDAD9of
CqIuQutnQyvGrTTJdWNL1led2gnelxbzzQcFVelgnPtvfLF5b5ckdZDKsUU+M0oA4gs1TVVwguCK
0n4eHveGeMddqLvWtjn56sc6A5r1rBt+z9zhoNwTfkNbvKlSdpXlI8xHE5JK5R4xIK9cUQfcP1S7
YtBfdv83Tp63ASI+sv6pBWUzoG33msr5OFVeMUsarViJGzkG+ycwQNz+mW0iUq/tPAT3wLhtousx
h5ktZZqdWP1Kts80ABKdHQFnoPA6s7r5/AMJ8n5jX7fy4kcJX+Dm14IGPnUlbbxxLvqINLFVNb/k
XmITrX2cl96pemJfp+fJe8d23VesKiXot3P1u2LRfWY1bFwQjjyQw56uVya6sVg/lRxNtpdhcLZg
JYx1p0eMdlzJ09KiMBevW1t03iGKnSdFDispnNLVIevyZ5koRXC/hqe4f/s9Lt9FYEUPU2mVIe6h
iTyXTbiHzi7vWBBBcsxB6lVUgNuvYhAwhr3gu+u/9TSoCsdtf0vDaL31e+8/608qIKQ0FMur3kGG
1I6BMNtsg5zxH1kg4Xfr00p3LscDg6Hgq0g7Yn9PY8BbHgHTLdBfrVGiEZZJdfmDd1HT/KhhtnhO
XmRF7wwxyHoh5TEyyyIL4XTN/hwbtbA2WB1FyVLSSS3Jc/xpcDOJGIgJBBJxk/Q7fUY0uqKAnWnZ
R2r/nOEbdMcY3ii1u3WpbgTEjN01z6rabp8SFHYXQ2zPsD20D5Arzp/0GuLRu8KtMqptmuMAaVkf
DJ5CQ1bqJ/Ib+KXelprAiuNTDpAtrXckWNSGFcTd4m4HIipZQd+M9UF2J08AXuXDR9y208iBm4nm
XVFk4Tx9ppPUvHfkvv2TLS7mkdvjVkzmTgnN2LLFkYb1sgkNcbuZQSLbQMPYSsjvdM/60uL4mgJi
wyxl8KK41R1Sk/FC/uodZTzej3kziXzJ10rjc/lNqHkbCZeq1D0aA16JHFJwQezgPzkiqq37ynuz
YkAaNZHBGkzme5+OMYjDSRj5jQQGYUus139b6rLRXQWKEV0LynAaZauxZf9n6KacuJVXIjyMTyQh
L+XzCn5t3camj6HzoFmAH+ccSZEedlGdvJ6gukc4MUmjBZM07VBWtvXcPXDY7mpkbg7Equx1dBx/
GR8FUAtAqamQyZ9VsaMk3cYpHBtkQY+XYcEbfQYJ52xWxK9FKCnThbEBnAPhpRQJVjD1MvsqfxYj
X5P0vm9LPMBzVboxK9O4Ew0ifn+Bb9BmLkQVU7NdfeMuBM4qOBZcM1meN3LSzPBn6/Ojfkm4NpBs
xWTi+p21E3X5TomXkdTxLSu/Bc20bWaABk1w6UAayJNQmv5BPLcTogVfbQyjvJRsvG50pHFEXayP
Rdu5a6VuA6wq0rywwbx1ZAe0qnfQrO5XXPDubJxs/davmfj5+C8jBfYTa3YV4ni+usjBDW5ZYHkw
b9EFqb4Y7Opj7mNfU7shTR5fgWLvtVBr/+jyE3sMsF9t//aGIbHznVH85agKAVYlcgAmhYffIvv4
CBMqdmLFf4jBIe337iX37kPpIw7OXOQ/sja50AJ/EBZ2EaHnY15cyzEJFKRuXXcXHYsVacWLHSls
yQbWfagMe9siFcMjsahE5vPv5ePOh3eMNLJ5b2ihimJlwO+2PZO3IyXGn+Ml+wH6AaMMGTwcE866
2dxSm9ZZpWoBqErQNzraVUkq0w+K0iXcz9eCZAIT6rsOPffTHrsm0zReFOLLlz8kSmtXCreaRJE4
obNpRy7brEhjLAxkajcGCm8kgWy+pGbdfe0EpDO2KY6iavAmM0tqyoS4pSTX0VDgQHsib6tfb02R
fULks0WYa4v5mIM4se2WZ91muZbWoTPkqHvI6qrI8w4g8cj8XMPXB1jy32AGLdZiEsf9dERjMo28
DdQrJc1j3XnUTJAO2ZkudmPmo6NVRDNNp+LD3vM7eOcAWNofgZSjE/wXSdQRyPoN9SS//iXu3PYl
bO0YcYMXvHgu98+Cqp/WkAY7xAIRsbKc4oxENUrl6XpGO3kuY72HTm5e1kPhUvmNYhY+pUlbmdEv
9BYdKCiBhoRpkqtuuHlcM5wwypxQgLxvaGsTsm+eZvwlQx/F+5YoSMb3FQ/68qXzrTeNnTBcFN6m
zSgHSgaSDae211cG6dgE53vEW5EaGW4rpAcQNQYPC2/l2Wb4NHVi0CHUYGyaIWSZJLn/pIhorern
UXKzcyt1p+/UTIiS5KnDJc5cU77K13lWx6t1tbII2/Ks6+TQou/5Wv9+2YkLHxhevsuL7p3ilWWn
mtCbfBDaqzepWGuaf8lo+shzXzLCmNVytUw/MVQMrPHI+iXnCS1S0NTZroYYKQdoECCIGpQIpOgA
ycdzGYg7uDpjw1GUL7y4/4iNtSwPW5Cl+MWL2McXnWlAQyZjQ4M8ls9EN2qk4i025rWZUbqq+ip7
cnaWAuWTeX5Nmsd+ZNNwtHSSPW6iG+1QE74fmVx/LtqlJeUDJfHu2hEqIvGkoGny7WX8OWPFYQbN
M9kAUImzG1jQpewbN8FR4YslhHRTX04hmfU3kd5WdUVMKk95R3fECOlRFomnRLykcAmJJJsy2x2w
2Ivn1JR/aeYPOWFHiyX09IvbwZ4LY+bUEBtrglDHVbz3EKfwJrKWDTvN5vFzlTL4PbPtAm7HmF6V
mWozqRslExySDbL/Sp7Ugq7VC2aZDCPbVLLg9lc66ZinMadHXn2WYrRnAIchAYWMuk1qlh0oH8qu
lAk8WC4lvTcE2lZDfO3DufG0dz0jNmLjzcnsULzgzW69b6iae6GFGtDMJ4LXeabepEu7tFplmRNb
pcp5b3NXV6Sdd791HTjW/bRUzKVU1qzJIDjDsVqTJjX6ILiv4pgtk9PpDX/Mi2EGkOxBjRDEMQ4a
nwybXC2ZhRZk1XnXvQpIhthBa6709eXipbNXLsh/yAmODiFthiNtVsgrcttA/wS2NrlEmYuOCXeK
3IypnIjMDUbdgOoctL89eYB9LqXDiA83GIqrDvkxRb1sfotFHf1qMmHv0n0hp0t6d8rLEcjXIP7p
4MtZrxHYyETic5Qvq6lOKQhcui7ljlhRVW/0t2Cb6TVQ6ENsE3SC7aYvmqsUvRXPt7d1k78ndgmS
8akYoR+Edlv1pwkWjpsizR1HWQxLDBEIqA+51elxhl9PBNfj2gemPFeJcSmf8ntQTWyMY2zZkWQL
wqVMwrD9KG4DQa+rVJyvS+KiEOuoLTV0JGoNBdBiiZ9FeDOt6h1SdesM2UDJoa5/nu5e13L33P/S
sq88l+cNmKkawfa/6oR6Q5Kk4vF21KtpVBpf9yye5OBY8cnieud36MbwjmijxF38W/eCQh8xH8wq
rMA1NeRaOIJZBnSgu+CDe7BCeYsWs48LEkcJaXGxIRkgVTx8eau9egfRZbfq3gG5EKT51O7BP4/w
x1rU3GCGfL+qA5dSBEXaxJM7DBZdeWScUDoa/0uWHq7Wlw2ENan0kC1ZwThNEFU3g5dJ9K7DO5v/
RLl/czjW+nz9FTTCD/d1Rslb8C64HpY434/VCg86KOD7HmN9fwHqbfK5lzq4+txGY2XwnoNt14XP
+9M3wFmb88eDlTCj0BbGMbere+6C5Yw3BLx3NiS80wZa3WKHZQvTdiV3SEf+VzdgclGBVh7eG9tW
7gXU+FD8d7hEzxEVczSoKxlzEw8hrn49vuk6v5VjoaUdauWZZHW8rX8HsHL5xANSixPpK0B92Na5
EG5Q7pcqSos7fISEHWWZ+rvTYidH68dRW7yE+yScUqrCaXSRKpKeVJjTwKzMpBgONyI8pRJq8Gmm
WB9emxxV5D0PSyPMrUNDL1rk8zFHumXO7nMk0KOYzXhhOE3yru4IpL4EytvEa1GCqJt645oy7jVI
nV/AGn7EK8LqpYQ9j0XBXcM1uKOjl6f0+rtumr8LezdBTqSXcmHKstbV6Swx9wl7wSzX2aXDrSM5
QXT8egdgsAFi4Nut9HxjAzttmW2NaZncWN0jkzTF3WsETc0JwbvbmnlXvcvoeU0HX1REnx4VbnCb
EyO5vjLwPA0hV3RG16aIgJYIa7W98YBO3wWSjB6ORK2fYjwxg6khz6uVuYEANLmNtiNaCTnm2M9F
Ge9Op3wgbyOLe9x1zFN/VxGoYCAQAKoxuWDf1Lwy1UTf9JYvJUF/s59ZRAmK9TnQq+z/ox+ffuD+
y0AiknrGA2E5XrOGkeDD4kh7ST/OaV8olwXoeEL7UEbONtBi8syKjZXvvEUkV4sU9gGHrI7/Vk+g
hZsEReVMTM4FkhusvHeOcmcpiuSBTlP86RrZJgyjK1TjTXW6rTzzckCXw5vyfVhIqKz3HHmaj0Cb
e3MFcuD+BZyx8hJBBtS9+4elis/7STZAKL54Hdh3wFxxUxMkI5QxF3+4qYVwZF3d93GYsm1ucRkv
AD2jhC9YDhNecNHcRczB4Uj+gmH/ub7ylC3zpyGRvsRPrN77gM4ElNoNEkgZjw1rl52/raoEmRX9
mh4b+E0tCNxMc8q/AuM+/dxAIzvJ5kj7JE1ZkvM69ho2hitcTXbTynV/i+8x/Zfp7aW8cwjiBREp
yKQYtdRf+7X4VZEdU35XFm+AKichLALdsQys5QC2hdnt1j3CTvPjaAPXNq5L5Vh48nY/LqxJ4jSE
9xzvYawAQqmMvllhKfJmBy7pfw8hY/3HchRKV5A4r4byL8WhTbbLAwk6NbfdXXg4nQwkQ2yoIjUN
e0tbgRraC1zesZnvouZtsvmwnza67sKIQ5mgpNVi3ER8VjoHZcNx8bTl74K5viVlESx9Kk4CVUxL
R3ySNY++BV9QuCgsyD6zrQUaiwvWQfoegDm1ej5QQq1PO8egPdDo9YUS5Nq8eJK4XhcWE04NNbOT
nuHRXdPTpQRW9sh3DlZYbILKs6yorlTsbnjQ40wReAnwVw4sfk7EFzIj28AV9Skk0/mNGHxuX6km
gy95aKuBvnCHChLQQ14368YaI98VWYD8Cpr953g3Ry0miT1t/jmwtmh6UroSq2xQ3t2HgslgT+b/
OE9rpmMCp8kCubRBOKv74S3OvNo6XJqrGkzPGdIcJ7uI3BDkRF5eWRYcxPevVL9qb/2blQAtq2f0
ZtOABtXG5Ntu76PYjRAdmLHI0jSqMBVWgjgave4Gmy+9iOQC90W8xHNG+V1CHgUENdiOoqw2doAr
1cHo0FqUIbN+8RSIea19kQeyrvo8U8jDgUdFAO0A4GnkasWQ7F6LRRuxxq9fXWn9SUx1jQ3d4Doi
9JfvYVptXjFbc6Jl0ukxJ96/KrgO1GJw7wZihI2pid76xK0AATyY+6ELbbMlT0JhtZh4X/y/NC1Q
hUkOVztzjFYuZJvrbSlsumUsWiRfrIsuiS63PRhoa/TGohUgs8NlInysZwTdVVSIMLQt3OrW6CQI
EAuNQE4NnIImbPhtPZYY7wTqS17ONzihIW0Ej+zn11omBpcyWSC0TDuRSccDmQnvVRg7hNkCnOsX
r3OF0aLPAcVe2YrhZGuhvE2smo3+s6blzqiLZAcdmXTvPXQkfUn2MdNQRhf5UP8CQa/Q5md9fRLp
07dXpbvjlCNLqAXeXZ4QGkpYY4atrrDcR99olgf5RbvdzwSeLc28wzgULcP+M6cPXYgWHzVpswP3
JjHG6WL/gdYkj+0FmVq7SIpe4UfRNr2b503c2/bCpt2UM6oTb79muO2M8nRTzwxrGv3596fHwUU/
8bHWUcwnGEYwdTZMViwzsz+PjpTvJSdD6xouxloOzOZOPQz5ac9/evN74MyaUptZBtZdba5PLExJ
N2cEicoLTF8p97sIa13n8Xg6wZLNfOt6WqK/NzPHPPELp2goWCkNl2M7Y945cV8O5qYOMn+AJcEC
/0Po3EkoTvcbeOEKUIVP1mmuxnEawz5QVf6Qy/xdwimxFsY3KsUUF1OaF9aZfkBNgc1I16KCkAFh
vF6qwVl92uQQPy8BL2NU770+0OltGRi81zkwP1/4YHmU/wp8gZN1MJYO5qONQn1wbxH4XcZvwCXD
/TOERTmiFlBXFHUm75KW7K9gKoac2MXBKpHBXuSSjPRQ728MQEfIw7C1maFkjQ1/d3aoXSHbQ7E4
EedD3+8vCUnjHty2XX4pcZUI/nGc9diaxK86i/LUXlGfwE5/A7RaGw6GpXIE51VimL+SJZARVRZQ
OXwclsQNzHORfqcCXFdTLupS1uvExq+CNnnMQC0+qlz+tIrXPNkV+vNywM3p9JQRjXJqqysWt1cN
tMlOdZDvDGu58AtCHx1wHCe6zXa3YrcqGgW48Isweby8+OcRCUsQ4sYzWwKfKa3RmOOdzwviDeu4
4hEUwLqAvld6CuBked1J3B+tZG8KPaqnHPlK0Ef1hy3v4aJ5z0Rp9Gj52AgbRs7KhsuOjpPsFmxh
VJccW+NrMhgVHTgFZkzwWdqQDsDO1a8kKi3yPXcoYyA9uHjl9uBfselR7Vy7uho5/O4rs30JScZX
d6H5FWz4QwaMBayyvx3MIYM3GssM5XdPnyJcRJzUaUsCLF70AUUZynQXZijEJ5gt9Azey75F6zYC
V0Nc1OMcBDDzsZfuYr3uG+tyUbQnlFA+1k44D6EehQjVvvL+Q1IEbEbbMIoMGPVJT4Tsm8CkZter
a8KYGrTXmhLt+yavz3SyJdMAwrzh/QJ9SI1srzAo6KK0ItarsNCCCRe2JgGp+4/nHTdElmUphngR
nA6b00iaG8ISLr/2szYUDccSubmJIdIxDl8g4MxCNkXakZaJsNXFJgmJ96pI9C2CGCOM6CHBADWH
DCRGK9rgSjo/+irNIZgOUmb4Z803yGM3kwBr7vqlTeiYtC5FGy7BbCjyqt/cmvYwlaGHJTrVnj+t
8z29qQjwn8Zi7sKfcokpWRIRLojBvo8pIZwK3b3U962KN38e4SG4e1uy0MUOLTczbhcZPJdm+9aP
lb2v/izdgYM5aoucmoir7nYEQdvO/9NvXu2JLGUQNxAuxRx9RmoOR0SuVCH8dkVGMlzH6JtFe7q8
q33B0OlzWKcRbsLzfZzpjRQdi7kBwncdhjcEg+6Uha4LNsrfOjADIZWtyVXwM+Uppfp3gS4tCtVR
RWUacR2jctmmgJf0+uH70YhleuB0gWLHpr9H5HKfaIn1OMVVZiIjrx1+ZV2YPQEjuZs7DiMQKwFe
gZz3vdwg++Y8P3rdxNEOUHK6d4Zvxnrq1KPLJhQH4Hc9VqoHg81PvjlHDmlw1kCssFE2vhRS4a0o
Bkvxpp1I8DjWDjxDBl2Gs2SRSejx0bGXT9YyK2IvJclNbhn7YK4nnRA1FQA/ZDq49tY+lAg0vwXj
02+/t7OjuyztYEz+yJdAsINzlquwAxNu9Jok6pIwd9y22gQGuNcP6bGZVe6UnBOHJnOHjJxK+yfM
v89xxzwnyxeGqehWpvyOkdZlZOhmPCOG2F7QnwR9R/lsfCMgYCiIEjoXxZCie2lcpyTLLL+DOnrI
FyYfmECgSM6Sp/E7rSQmna1pybWD66fCWKHmpfCbOYMuARUYQ/z4wpMdPBDVpOMzy5Bzd/by7Ezf
R/+/470MK0DZEzm/2xWvUDj4rETloVySUFZrcK9UUoy1i7potSyUehOkJF+pl/pDgUZTGJ5gP/nG
NK+gJIjiqgyLs3IuARn6m6lySEPp7jGVGbJSosPK4wg36j7KO3MTVbpwdDdpzdgPHSJpQwMfX6lO
oAlAFPrPRS6iIYRIXZnebp/8rVKrsbH/196Hj6Tz/BBtyeDRyn83URsgGgyo2ulkCnisJ4cYIArM
6pcq+sWA3c9KkD8Vb2CYasv7B3mSP2AAWIi2ZQQfo2bXvdULkjaC5KpX6SAwmJPhInqlDlE+xDkF
TjbvQQCL/LDyFmwbKtk8sUjjcSjpwH7VxVAVGFbER3M4RdpaCstQHMWITEYxbjL3loBhOq7ymiP4
gVe/9qlvOphKvfhwMEMULVbA9870HSdfkfaYg+z+Gv3J58uDzihfn/fRkflM67jHXRCMGeoNGN81
kZuTEjBHOjFKgZJcrVRKoWmAN5Por36ZlgaBWNYTUpQm6isCRfedwe6o9BqNikNOvCvt1yhaN5GQ
+2Wx0Z7ExdsmSszVZCuWjxxEdKAW9fKwQr2ASRGa/EVjLGU3FKzVTVbn0OllShDIHiCFYbX/JU9G
0k2m6yhHBMLevlXf2TSQMMaMfH61BEJ7Woxi59sA3V9Utl176ZPv6/8CIJ815KRFXorC5wufz33b
eBZklPXBrGqWtEktfnpklffvM/BsOoQ6e4e1iKe47g7Ezm19nlOVGsBtKStYaFY23SwQ1ta/5rwX
DIeNv/eSOjI9/gJiE4khqQc2vAlVJvArmHCH1YEr8qxdpOdLmwGgL9orY3hn5yoRK7YNyIpELJav
aA7YEZvrvdMoqi4QCvqcnYWgZZSkWVrPv8Un3MMNPlypG81GNDqPVJblZqZ8UfR9+ddd6oK3JeC7
VlT6kDZ07eL2rH86rKZcrvDSdjBXF5LqJFmJboQ7UisJgscn7OC3lYJYDSmbvPgjcwm8gW7ar2Xl
4lrmajf5vLB2pEbXZ2AoMQa9raM7DSxLv8s5lTJQlr5l5OON58kQiV8XThgbwgcLEyL1Zui018C8
ITsw0Qh0/yY6uAT/qjUsBFsMTqe3bLnRPM6BoWMVIxkkMhV5mTPq878FOU8jLZsuuWRblDUhuDb8
G1lWa2ZH+3qb4hu5F/i/uOFhorId4mDi+lbeDJoALmS4k+gSGtkuwHr4Z2sIQgAceZjl4CY+Lca+
Zfr4g+wNmb+wV2DvJoZ+xBsSfeG97xq9wSYI/vmRZCvCTrcjZh3vv72TiCvXwdFrXfuHiKoFlNFS
u04hPt7lTv7spKYZ7K7YAJQajxeZDYmwM0bf74iZIYyV3b1IDg69x5U/O+CHympP9vMCJzZkBmOQ
Ze6ez9MY9Avu8H7KHp97SCaBnL4r6SLmpYecKcx5x9l0xGmAOXyl2R12b2PjgZPwmFzWGnDSZCPE
cb7AqsRdkd60V/pmDTESCKu8NGiGhQirsdI474ErysmL1vTLzbEdo7gK1e8cwaplIAW/qGUxIDvM
gc0/nVSoP2GddDYZaECmmlXr97flUiWYe9vAMNGvRPwRP4SrkN5YHxLYRCsrorK6CZN9FxYVZAm9
CXNSaybt6p3XBzzw4I93DkyBFLYGgvtzp2r7DSo0i1XzOSqRBcdJPEhAHpuJd+K+v3+mMWjvRBNi
mjQ+dgvg0JNRpRB2vRl/Br1wZ1UDLcoQSH4BGOhiMJUxaDfgNTzSQBplHCcHYHUGOTCqCNpCA6np
LMlqFGLgXMF6oryYXKCnxHOq39eXsmKeVByzsFS1u9lwPv+GggD1neO5QYWwRAlGBHOEvhjQ49Pc
P3+e9I4mAjrj2HWhQDQ0OKvkO9eCMOMzXtKUMl7qP+EASW75vj3dJ0rioyaEuuiqHy8QkNctnGIz
k1LBAd+6I/dhDO1twU8Y18mZ1wKBqiEM5n1l2ntXyqRROW5L3SsL8CICFP4xiPpgGUywWBycn7W4
3CMJ2XgsF1b8LypJSvum9503kq/uAAtG9cSQ6d0O+tOmh/ZUkBuV2h4Ojsu3NGASYD/e0KBghCmX
nsM/hbbKnO5v1sT+aXpkM28G89tXJlGf3txZN9cm51+txLqLWhHcAZRxI2ko7lzEwvHnKLlfUBcb
A5IkEIaFfsySDLjv5OFBHLAqMqlyaF/DNk9Hw8Zkn0NSMi3NcjexDp0ccMbxgQx/N6LncWrNMN7T
xwrpky15Ivpz/s2jP9Kb/YAFgTr8LHEwp9KbFKgU+lu6zxQFjmr7AFwJrKTQ3CYzwfFanBmMitwg
F2jkPCqtw9rBl70MoVqn1afRtldIFxDUmHd5huzHRGdsyhdi6LrzsKCoXQhEyi6oAdC4vuoowhqe
WD9tzwvId49C75ieCMxN4wCgyzIym9ljEF9F7LKIFX+oF3eu2qQ5nHhqXZrpiG3tbmPeO8ndp/YQ
6Wrlua6DJ6+jF0vE9diiykqa7di3DV6bULwW8m62XLLJ90bAUHFUB34aL/i/LcYveS22yknQnEe3
FDZBGJKvSEQPZ9hndzs5rc5XizAWblur2dvowj/VAzKgmJbKyjTbQvKjwh+WzdRl9QzQKhCYhooK
1K0+yLlz9oDln1L8+hAHsvomI4SokmdHu7qqnEzsfr40hGICUayV42vwMa1SJW19SpKeoTW5H5nq
lErsqrohu5cMTC9WNCDjFQkS1Acgvg5iFwrYG3cwKRUK29pHkLAU9jJxeKyJ3/QP7y+h6XhmGlpz
+qamAnF3Mxb7Zv5t6svY3VIJ4g1b9/j7Hp4NsD5ZE5bN3dEuu4Lj4RBLvqUoZR9c5QY9a0OSubcy
w27xYERCrE5qWr9wNGDu8fr+r4zLGKGmBBAw1WOG6/m+qZeptLw8gwacYuwK4kr/qRjVr/eVU1qD
ehcMSN2awraUk9vHofI1xozgZROYkontltmvy8gT3PD31Rpc/aXviBRUgBuahscv9pDQghEcwj0R
/uCGBrmKd6DhbvWt9rzZU2L6WV3rWabZsl4RpbRVfIolVwOSaoW+RgbfOGu3niwaqgHSJpe3nYRn
9qQJgZoyhUADrfoM6zg6sw3GrRtZbn/1yU/soI1mC3axzl/gohLFRdJoIq+ImHrkfUcn4lRSnzVq
VJAAKEr2q0eCgobVXGQ5gEAkRPZyrLrBCz/HgmOmPhWnO08xejEh3/LEwM63UayVU5lI1SDidNjO
3xNN04RosE2f6horCQR7zqF1YN6/Ym+At7E0GQrHMZ0/zcqdCF9i+0kY6qzT3/LEZUhAgR8mUvMk
bVZNnKDxQkEBOmA135DMrQOEtS7DkkXvNFVqeCbmVZ8His6STMkrkHX8FQvd6ir6CdTdCbE0rsWZ
jUi0SbVZEjuxKpfc31j4UiP9ri4zFRknF6IL5Yn8dHHyqBTujWCxJzhHZ1JxombbF/m2AFL3YPLx
SI6bvDu/Q3ZmJ0XVgn4eONf42iGiRHCaGfZ43jzRUby/JgsJut751DFNj7yerAb8BhCz3tagupC4
5cHSb6CWWHys9BvOGcQ+c7ughBlq8qC48px/MX9JwYA1lK87WVSufEAxDLTSoeHp95Xc3DfU0ID4
bSeoZGYB7s+sx+S0+FIEzBmXFkUw9PVEw1J6OZDzHVN+aWhvxJFf47fDt+2g+kt6RweBJKxGNeyz
UprHq4ht7zJIQYxUEqoZhqdNyybVG8aJA1CVwsrIcyk0EobAfDgN1Iu4JBiq1Mc3vAE+MaaaYwUR
dS7QrFBkfr8Pp2rvYLIRxaydswlr/QUiju3F9t5niRxyuBY5fKc2xW9nqNFlSjy87ytiaQXUX8s9
QzN/FoDhV+XC8W/79AKQa5IeuOCZnLfcU5bi3fOB9xfN+x33dcevHGKg+euDAOmkSC6a5RinFidf
aBw7FuS7KKaQz4PA/toxdnaJ611feoe+i0yONZy3M5yFmX76jgt2/Z1Mp9sDNEAjgXKx842FeeQE
4dj8MyUmHT9pDiZkIKxtBq8L6bxOTthegt0aeWVGn4IkCw3jm2Kiu/p8vhDCFIsKXWhmgaxKmPl4
qN4DKva8beAORDjCFz0Uv0t+pifOqCDUiNjq2OIjNYpbR3q0/kExgFazvxVJQqRBcDx1693N0K/D
gSjo1WjMHHDQMsleNajMK5pA/pOfTnV2Ztgt9Xzph9z4zBQLAntGK5UixiiXt1zk0nnmn5lTvjIB
umApUSNzRP+0OGx5FWqga2adpVE5IFyYe+lnCavQdJxlsBuLQDUGvmb+hVZPEtRmqb2ErcIBHDfl
Wjx/SDa4ecBUf3xF40EUxGhBA7gTf+dpvC+VFbnQJLZGgKexu4XuBdu3AoLFeuVO6RGcacMZAG7e
1sGM8V8/KWHkJty9N6J66nrl5fNzmAbvmBRLJr4IXQ2zhFj4APqbwB5e3/XV9OWlqCvPOH8hN63G
bsQD+bRcnRJLcebKhxBc+PZByLbum4oUeKERzD3R/Ue9yc7vt8xFQLTjnTvd/I72urTAIIOPYSQ7
EYs9Pt0RR1dEqNXVsG+6Nq6JLcbvqKJb1hgX6Bvim/kMUP4cJZrb+kP1bawxi2jsgGZ7fb3fxGDS
yXKVrgRi/L2+qKECAX/Pt6qLr7m2fVJZUHmAQm8lEQjmrgqdIPk51E4+fRg5dMmG+hN8Uc3goGdC
t6NYWSv5hrtW1nqEkS82NB9RTIT8Q2YS560u0Q2chDEDXwnpUlJw4pk/GWdXOWrWRglRdsfFi9qT
YeqYNIKqaepm4X7staDK3gP7N1OsgntY11E5jPA0Gx6fFyVhqDzX5FoIVTzekv8My1a0Y1CjQXXz
WYjJlQ/Z36CYkOCKTgqE0sA/kyNc8slS3rHFopWWMeNJ6zCAxLt718fm74CGyckKYK6BPd5wmB5b
MwBzhWI4iXPwatfuqFgEZJ/C/j22l34VIy4pFa9ynIGLRIg1a5IInzS+SGrkSz9tz22dS/Ce/R08
fPNEORi0E+U+u3CnuKIanx9gQBBWeF+RTkCudNhtUESD+w4rtH22tqOo0UKKSgqrvBS4WFY+fOSx
nY6ZgXE1i0F+dEc7zct+cJKk/W+P2mTqby/2VmNjBJsV3zvAZDLjdnc6Q8vS/hsf6xWNcdeUmPAZ
UPBtt/rpy4z546RrDAUhW/2YALIhcywsvFIKc6aji8rV11TubTNZ3hJePLdU5OBSAJCldpW/f2Ug
/IlCCZgj+fUJn7/Quke0FeqzAZQ/1umLKaFwOHwAAURs8pYKlCNiNJfJqpoR3iD7yOZKXtq+Lip0
Pz8Go7YbGmwVtWDO3WOQj0t+AaL7M+e6djWEEKhqRWQ8PgKWsb6Zn672gwfVbKgvdkZDYw0EUlyI
XX/N8sRBIkNlXTtE6uPi9HLwPy6NdJrS/oqUHjjoI4ryvh5ZBCWgPwy9OYTLjmFCq0wmwiYgj0Xr
9StqNII+i+KwF4kv6a1aFElr1VmFv0Ii2Yitljqjn2V4ojN3ajB1jO0CUkQv0S2MOhXsr4QkHhCq
IAQ7XTQ5ZPLO2oRjktP4XThZLbVXxpmfXUucCSnQJ6zFfkzlMj3XUHvoA9OkN98m5yeC2n0kMxrI
SgstQ44raMDs9mlnaGOiMWozItNjmFYytuicJUkxnVHfvguRV/iDFl+y55aRvurWIbu1EDpBdVBG
NNxl0DekaJ21AZ/9vEgatwwwwAfG+rZh9xRfINBz8ymCBgQQW2bDW7jOtYoLI3yOhTMwOYc3TDbJ
Q+A200KZSbgcsUoggWGcyHSzTBgvwabepQwTWIDbPUPrhCbFjnNQxVh7pp/n4lzbRi0OeGleEA/z
xYuAWNxHC9xIQVf7OmCPknbBgz5WcUM0IMYIUR1DP6K1jpb7llm1hcHAuSYFWZ+DzLdm1tg5pZwO
ot/4+IPKEf9IUiTyo34LaiMMOVvL/EWOly8aeD4HwdAuJp/4ZIY8fcGywSJD2001g0HhTqPHAnnV
HK4+8qetlk68m2VFVAlqHaosucPvfPqvNL3idmljL8/YMACl2oeVUDVKh6LSWwXAimt6kzkCfvBN
VRgrUErsg+ylgb1ZECcX+oN+LVx5SzPmhXBYNsXQPzpoRZuAyJ4yTpAg85c2SSy1VR0iIa5TADlN
YZ/p08ARMSu38+EKRshGWyvmwHvmIZgzybLuC99gIxw5zmIU/MXyTj/CyDeVvN66EjC8Bb+k+RGy
Iu0KmgCAkjotoIKFoSJYezmbx3LfONcOml93ZrMfPTXcfl7m3OPn0NgoiU3PMa8Unln329W8tmMa
BE1iN5Dz8itf8V/QprLHlJjUKbSsrp5xGvP74zzefYvhfOYAbF5NiGO/Sz3oRPL0l9tCHIlu8o46
fgRessjYyYfXSBe+SfWczGQAW5nCFFMrA5UvdcXRqkKOjV6Y5DUJW1GK5nPSXhqgqAk/19LOwTHr
cw3C2l3XKn5NEIoVGTPIhrK3N52sAixFisVnglmOdcvGViYzLEcfAV6x4XZ2tjVp9RagYLCQPNfc
urKU8/hLDAmV5jVYZCxr9gM80qzwKP9i6TohwAZS9igS4rn9/YIBcvGPABVws8iqZX9cKbMyFsjy
vhW10r45x+WL6Q1hEj2NUuDmfC8xOW6iGsW9JzqSdWcup44U5CAYsNLxOV4kwgQZ4Iu4F1cYTpdW
AcSxpLgKNRHF3S5koXYv5QG9xJufeEo/1OH+aZw2EEhGPr+dZGxIt8//31Y4TFNOmkVlkI42lVL/
kbk5/NXYgSLYrSCtvOauEZOAhZHDfnM4WoNi1dTMWzHwYp3D/raTz2bkBLZyi97AThd5a5SdwF0p
yPqNUZiVnH8aNCl1uN1KKRLWo7JK1Jf21MrS5IyxKxTFktch1c7fM2wwLF9UrgpyfyjwGXEylNP4
N1hp/p6YsnfpdN3WJ6XBKQYt2T51MpVgp0e3CYjnzGjFiuMgbhB3GPQBFXdkgv3LxbmK+vu06Xkg
q3FY9DTlIe+cOJ2EgjsAOpHADyzjzV7PLhAVszcqh2px8SPHdYJ1ANDgQRg8hLp0LSICMvJNlHA5
wIMSAmMoQLAwT2zHIDzMBqplqcCmQr8gLrxXNt2ZxheaRjz41B7UqqD0GOe/2fIwZ3HPDro6s/NQ
A1nVuQ9uXpXe6y6RzMWkg954mzl/HiNm4LOQf1A2Adtql61N87jkcFRsXIH0SYNVMQSr1htgfUdu
rbS51HI/9VfFA81udacd0kV7fvUWehOoCljYn5vO1FWXQhz0fiXtMobG3KKa6CsLeIIOuXcCc6hi
L+H2aTzOzfVfMGY2PCtrCcqEGwBBrFppRajh2Z7uvNUrvpyJL6yZYhoP6fGOgEWnUDZLzH/O9KUo
T2LZtbpuBrOAwUvi6hQDEjPh67nnCWDcJVUFStniJ7MmI4o0RAVJ+KfTdyn+wPowWYyTeHRGuGM+
Il9i+qQsFl9VdLdqc04wkt+J6ESUdpDbekqTEqCTHD+DLzsWuQ+2jeR+l75ge8Bn/1IQ7bC9GigD
/Hh5ODzrWfV+YRiMgu21dBajvJI6SSaw8/xnhxAG2Fgdg9zVf3QOTHPvR8fPmsnMvSywKkEd+veO
z9+WdQtyaXEuuM1AByjDxN0zvc1Y68Mpn2DJ3IbuPRKkKOoggUW9YM6AoClnWw01EOacGMUR5snW
ea8wmYrEL4MXFEMJgpjKFjR8Z9WLDI04bbF4RFIEUNUQrIZ0k+UKZIB8coBVZZNPFXFeb/wMsu3M
sdNNf7PxO06Ofo5mYwFCWGcxyC/tW6D3c699SpIp3X0xyRVpqnWsJaVs1YPFAzWc71v9RLU7mM4Q
7uNBynmoW0KLk5pDNLChgeHwjXDUdxR9bR3PLtdKi0CMfBKchU7OyAosMTxr/DzAA35V9g6RwE1T
d6oZKs8rot4T8DQPjEA0aeGMIFn9c7uGPgQrL37a3l+21S8iol8PJcuLgiD2lPKo0Cnxs7T7Ivqe
6yoPpve5DcpxcaKMkv6lrQnj1GCQhXxOYZ+PUZINZDGC6NScaD1haD2CzNtUp0bLjLrXPeNH/x1q
R0yCrnJpAaUzDCMaCJgAvDaTLVHeiMXSOEC8gwX96zym8JPn8aKgavhvAKwHDHouKl6ZJhsz3fwS
TrdkbegGxAihBnjpqOoV4qyX8fj8w+ofEc0UqO/ibXq5xrwirrNF6Q0jzx+3juQ3uFVF3OwxX0Oo
uWA/kK6zEQNNcqw65qzj9NbRyibQfJdRGzrgu/kB1R2QyXdGBSpXduo3LEOaZhXpNciHmsMdTcPd
yON5D45aaONn+RLRHb56+Fyd40kBj1tRCnopRVotyGgYiB2S7vh04OUHdJSWEz8kEdu5eVuJyd7D
TDYpYhRh4WqDmDQDYixkVn+6/7iGHvhkNjLabu9Qj6/t4yt1mw+rc6MlPiDEshgSt84sTvu26tCV
iuq1z4p8BLmwsdD/06oPb/a/7LRL9OSAPwr1DiHnqaV3z6BZkkE6EXjh8/zimCf+890sq53Cm2eU
+44a67tSLqNkgcutQISPxtPBx+gP9Kb0en2uTIQXCnd0drbIC5JRGC89wY2QQSClNOHdhETcg4uE
Rqu+1rlSC7ZysTWzw+ZHgIfT2n+NOknDjD/3Ao1bBa8WQyd/kUqN/+y59mt+mkMlB0Sl4jRlKE0U
varuLyaR2TdqX+YuLhRUIAM3Q7mwh82g36PeidfPTh1c08LQJpSc0T2HX7/AwCc4FaeFxSapqw9U
Nh5CqvuDol33SIqokC8BRdBNfAJ0jlluR6kXRMnDBBbnINb0FZ52cPI33YSwjuEskjTJSfU0RPzp
ijAjQJBLTGthULGKnoWvd7yMjd6T02rtUXmzw6hwyiUTxbMKHg3iFA83BVTA4Sq1909g+VW/U4Tv
5odl8+v1Pu9zToVGXnRD46u1p5x1RD9+gIV7SJpztXKaBxELhc8YBjIeEg8RuoZJ7dcy7kb0uZa+
wVgcil/nleIH35lZ1Hz2MZ0KfqLuDMpLjCaZTmTgd6gXobsN5PcsDoLjwpdx1J48S+4gq+wrGm61
p4l9t5JWpm8b6jY0tw2xLHGZi2+g9UzhYuW+EpSCHN/JEydGHKsUMcfC4Y9gIDyadxc3S8QhGEx9
TPd8Ru0HGCvDbhA81XlYc32ywmhRIe7vwEEuAkjLaWn1xZok3GS7JcqlmMIQ24n2p7gd6+CCHMXb
72bwxftQSgpXL3MYqefdySET1Cuhu24eWmKgTktMAKV6c+o6dL/3ZRTMjBfV2Pkff1iYdP626mi4
VaGC3j0w3OiDhMVL+elS9bDw72CF7LdP0H2giNDqq6FuUuahZEdABC2IYXps9W51TH4m+ygJacX2
UA5qO/G38MCSl1QMCVKvnDoo8tTvSlU5S0APrQF8JBCS1c0kPBqQneC0B5oKv73vXowBVU3aPNvS
ZPSqLTF0FLi77qfoeXZ9g8por4Ptoxwuw2+hr9jFkpbnt7bRqMMm91LvQbwTqlaaNxictfxHsuF3
3a1so2nelScYnX0CM4NOLOSrvAqx/KOfDPBMkY+rDK36/JbmZ3B473fx9fgXs+Gt+AtRzBeiQnrE
eWmKKo6/U7klKuI+JVpq/X4xOJXUe4ryvbg8prskH2uIbhea2BhboUk/v275Af1SW7Z+sFXvOAO6
RZHemzixx5RLVOocVzOTarFTKuukppCpBzrjxTdgLyTt67ya7ViEftXBEZE9q3ZKivObQblyBNpD
znDohnYXQfUCAnZ6RxzpDEx4GchQbjV3SsmJxhr9jlOdtCtepP0O/lQRtRHp99RhyrvYyvd52aRn
jB+PsyI23fNJrnuO2GVEj8LNC/vV7cqmg4M7J3LRlCvFLFr/WqNDQT9I1X0Ur0tKpbu2tlzZzsrc
savoG8vRkyGxWoYWZYUPUfVGCOTavZwrSWs9ackC/i+iNJq9prfbMLWeUFKY/CYakuWwM3w8LUD5
Vt0RtYNxnE7WvAEe/e4sOWj0trAjm/qo22R/0nHgjjMRxCH7oopoK5/cLoxHNB+DNBTofi7hdxVo
F8B/gI6n+lo8SDkvE/ol+oFG8Y/tpLehrWzk0+D34I86eaCPKZ5Wt2mo9iA3duSyCXcBBr9o99UB
C23ySdfrTyM/5qJitP0/5UYdvSwNexI3pEuVzAlj1G6IRwgW9rRpeyCUWRwJFqbV9HTa6gR12F2n
7Iaxx3LJca0bvzJrM8AFp+sHwyXMXJvVg1mWPqIEMahbjpgMNTIxMlzoGL1hNbbx/jGkGmQpZgmf
EhB80k1JjP765iXW79Y6DhkUU1o8d4+uTSP3+URo8L99+bqHXnp2V2nd88lj5jO+1q7dlKq08ccs
qBTpBZZ3jcbzZCCcus9M8H4Yetd9mXU4UVvtRdXli33YxrIvhBf+sIrI7Xd5WHQVxxiXfY3jiSzk
PZkZiDXzSuNmDEYm3/FVAOOUCKztU1t1VhScYUd9cbnqlYJiGfCdeyk6c0VdYkLNIk9Sz9Rr3Zgi
8MyzsxIIUzBNRS4rfF7w0X1vevsE8nk69VTcSXbnfdZyY7wWN2pCh6IKowew10zj5psunYhb9ksZ
YhoSdWArxl6us29FRBIwAEDjTQT1oi9wFtAqg7DQcM5AuK5mP2XkrPk65myjnYYzZavOX6MRGyZd
5OK3Rp2E7cYUCtE7ws7aur6MDjEDcQYQUrUlkyjehqezCgG/nyvyTr8trFMEh0hTJSbGPeoRRmb8
Hwg+ptI0PuYe1M/TukysY+6y2AR4vDYgvYbAP505B4sinyZD01NECpYSi00J1QTY58jw+3QoCAyw
sU7RII4P1dJeT1+LnthaT9FhK1CEpunzoAY4d//atnm7axFak3KR6XIZCQn8SS7yXL9oVTNnyF0c
rnReU22rqOGfuZeXWfQ6zb3hTxIts5eMc9A1Q+k3mdOQJ6LuLqGs37yKLks7oZUuWjVNSGz/csRj
7R+O3rJnCxGKosln/eQjES+xulOr2NrVxzgq++0oRn9SSnzEauSIW0/+uj9OE9u72FxvVLP41hch
WsjCY+BXcTDV2x4oUx2jnKakWVJrddMmcGQWexfB2BjTIY6khdEIKILFEiU3M6kcfkOCXz+CKu1r
CHxKl7LuOhrwTrUvzfm2lib8H/vyLFovnJJKdWpnHXXHg0wl8LKcB8c7iYfsoQIhu3orIKLfR5SW
BxAv4KJB0HSiVdGnshpo4uOZFEY/6d+/ZQ+xlfGfGHPLzJ5cYOtXAbbK09zS2f52v7whegyoOJI+
ABAEyGWgj2jexEX5FymhdcGDJJLILgcSy+mRF+5WFom9JhZkJx47crhKg18KzzAXRBXL8tudriHF
VLX4+mV8NEbzqxP10UPE3n5fEbzZLMbzGdcX4byfjps30zIm8BKVYeBAcInaTvEwetx+bp/BNr1V
9RuU1P2nguBB+FgFdymr5lfD95SGAoV3f5DUOidauBUjtS591vTBWIstdA02S4Y4GEh419S+30yJ
vtHz56+msuLwMvoneGj17zfkI6vtjY8oJUTmeqRFosmVdP6rjvn/pYZ3LQD3hfl+BpsZPJu7M1xb
+KWh1goFMrnF+1XiafkoghV5zh0U9KMtHHBtWSYiBnQuWRQ5Z8Uof4qP7gmLl1bPK9oeFkwhWViG
nbiGL5dqOJyg8dV+yg017CUWMtDhdzWzloz5qFzyxhRYvlBOutaHA7K24+2Leu3iHLqa6Wv3rbbR
CarD6lonK7H0JlIJS31/eAq2EpaG0FV1VzPBhrls2sqmJb+Jeqf9vrz7v8/wm6BYZsuXjT6KydJH
bVFxz14zR0WWAjgYchcha2xJVXGNcu7K+CCo7/6NX3OodgeNgpHOLtn9un4LXhtTpgR98/BSkcT8
ySevnsOfjnFHLRmjaD6ySH8eArDPsDPPMTUtnPdV4b/wsWLUrTPRbR8Myxu9KDRzAohS8TVQh6Nd
eOXMAWt3k57YjTcx4mwcTD0wZfSZmmvpsby/QYsJpLqoURBXPKj++OkdXEJjS3IbSik2T4AZznNX
ziS37NMmYaKMxW0c1lwBLsb+cL1pDZIOZ43B99LXbXx8zqlm4qtxE+n3jOUsDClaAODDFkeBl6IH
Gns6JdPlBT8rAr3cW9mcs++y6AgG1zDTL5TfKHBkUdi2IhTd/6HmS6qm/2N+DkGjx78xURn/7hJ4
0l0lLj0QMTTsmR80OtgWBJ5QdgDoNS5KN2H64OAiUEm+Ytlc1204ps5Y2HTJrtunL6bC1PuCBKF8
kdr++keNIvs9aW1LrBo7ZaX+PRbU50TAVg4SjKIBogUgjrfX1KUKUBkMeveAGp71AoVPIA/1xmCY
FcEbuqbDy55A1kDzk6IvCfsXUoPPrqC8VR7bWK+jcRqjaup1OGbG8Sx1X41vP8uIBN5v1234KSei
S5yDQyQwdWAw75Q13ct/cF6AWB+FDGsSI69vuSivfHgUs7/ZgjyNgTzRhn8IgMB+WjDG1W/2mDDf
zVKR7kRjHEoIXVmZL0023jlgDcgnfAd3gnexcIrHHQPYekKhNGfQzAyHaUtNbMYbw/HHMS9hENwi
BqC3HuozVZpdYk7ZCRcSEoaVcq6cWNH70zVib018Ipi63UlGtFkHCKwxGiMpXWlAJj6Z1VhTvGY2
uPmVAX+vTtE+igRWKour0d8H1FOBYXTggPbpw089W26VE81HFtlTQRIRA6sphtgg4pLxsyev23Xp
U1ZsjDz1x1lpj9JFECRvJNiOk0kketIcAKED7HUqy/J7daPKz1Nrpr39JTjlZ6AopdqRLHMxi1hr
EQY9loLmsjNLFmgVIVKoankUPd6ddaK/4NUM5Ghs/KXOJW58UFtQ6rBSeJYx3aJhgtVyDtx/5nD3
OuBjMhKUHHdm6inseWksE86TpWNTS+FVRyd+YFP0/nrteXpO8CeaeaadEEg2KORxCRrcAa3ph7p8
LePHVKaZjjNgpwNu3SG/YCf2WWrWkP+cCGS6NN6f0o4BiceJME2yikUNg5t0mtu4wGqxWOLjHYfW
HPpjlnuAmtvDb2OnYI9ajaIt/M6VIdeWCYX9QJY3IvFxCoF1qvVS+W1UszkiCIaQl1FRAwtvd7uR
okk/vsWza0/fM5UChxasMB69S+yBl+MgGz9ox0vKWuAR0duabZQXj2Jw8XmVeOMzb3NW6QLDQwZ/
ueGlEE5iZv3W3HooOEfe5EcdRYd0+zLTFw+0ZZYwJL4yfXc/wSlPxibSHReCOGMwDS48JQ/yZ3O4
af9/I2ytKrN+tcvjQLpeIk0THHNsqK9mKixvlPMiFLASzWMmuCRRydA7i2B2sbb+jfNjWi2dKTrV
7Aqhv4FIJPQLNWJOhg5TKhO59e8QUnirhkn6nf+atKk95DX/I2oftK6gLiY/6McI07vb8aQDStK9
D8/19HYly+0DCgWPs/iGbFw5A3pdJPtz5V49frmGpBSOBtHjZtdLukuOxAH9l3/zv0POc7UOXkvT
o/iELfi6qJGSJbVCbQ17TbXCQ7txJfr0AZL03lJ/sx0q1/txltSL1eMypz7ob5668ScK2WxAXSLi
l5azQ9n1LBXpeD68cRI4KPn/MQho6LzRNoXSyc2YZsv4VWIgMWUON5DS0Nf/pL4fyOB4B+xUwl1P
QYyw8lFc/rwRv9p2Vf9fH7SOcS99RpgnWXsag1zcs46krzzh1nW8HL6EBpzVOl8rgqarMPDVN0Eb
ZjSBJJYPadYrsuKDNrrzB624LO4E0LvVaG3bZU2ABn03bYW5DBybJIIDh1TSPJnFyRu4DmhpIIAQ
r1oeX1ufSTNU2QIh1CGEru7KhtQrZ3CVelDM23Dn3r7IlE+cLKXEZCJoJ2+nOzA+ZrFI9RuU8RJH
nhlYeGisYdx+bYVgfkcOBgRpDlXdnVDyX3smYOrp7eu8tgWfOmjGO6B1jqwSOkoXiLNwrpf9/n/K
QYZjdl4ogHwAnHUo1gSvyB5oyXm4pueoRCiEqs68PkjusV3PEeE8nJnnvUpUKO7BdOMm4uWx+mkD
2ObjvIk6YXdL6d0dejEz6A5jXXBmx2m4vCQdg7OPcyYFE5gvi457bvtWw2FEj19OQMK1xBPdSAtm
YfbNt4AVEffnQPbjUX1AxjQJuULkmLbu5IJA+1Hmxzd9Mp+DME1GWYlra6jRQEkTGpeXAOEyJUW6
ATCcD9Gp6CWaYJ5slAePHnIaJamveFr8Y6uoWGp+/vJ9DnPGasjNMgBXZndQvu+XWFbttjdUK0cM
YKwSt1Z2NwemgG1KPKb+AQaKz4Juxu5FgHpwpCMn8LfJJfBqB5HzMDwuRbvfD+oYD5hlPJQ6XqGE
BnWmYSNbEvYCtBgOOYoMyPzFCA07Yq58UluziybOvCZ772ZUcIgYv0PCFoKaWIDuBsvjADBE78kH
Ct7ULBL1mD+nP0yAdRQtTOX5nGGAFAGBnBtJzuqDUfdmMXCgqes0V/Do81P6TT7lJiCbFzn7m4ST
DN5RKXy7mx2/ybxsBCMd8uUF6EfVp2AaYZyRnCQIfOTQUBMVpVrzgTBVZgT7dcqv7xQRwxrcC6oF
BhsXDSk4+V+rUOMbNjTy7JrE2cBMJVmKQF1IOXTBU2iqYC7xepX7mboqjqbCTLLKGeihwqbNV9ug
vcyc2qXOHf9BRi5mg7WJGz8vQld/dbbZpF7D3s7C8KwiBEYbFpdl+92+maTmH2nvS6pwffSOkSRP
fLcg5kSX/rNkKYA7iOI9J5QcHZGiJN40o4X1fdjHITu49qgOstpmunCwR8AuDDUk2lrUmT0rVez7
8K7LYNYunz4shXlomODbl1EGy2UIhpOLNOFbt4Lw75P9G9FdYxW05XiKG5Oj9wmHRp/Xci37gAb3
98o1lLS9x3LzAewtJwUFcsUiV17yc5i0RK0cuTmYVr7PjUCHMbM3CRun+GEtiWfpZrxexRmDefGK
K4jZqZF33HgngTxcEJ3ctdk8I0D+Dv+I1TW6AHT1GLtCK3zPZs3TuZK+PjdonQa+tDvWgGjhzc0S
S9NrLWvItUeHFV6VzU6lGc+i16MIymNi+hwZCtc40QilCM6RzRZHNID6aPOPjD80px9H/vCbv5iB
K0zQWqpmVMovqz3llA+D0l+nBLvKUrAWsZU6L2b2DICEUR+rdcAEm7YP9oW7nRFVGZFX2NYPoTZy
H9SpxrpVdfaBkrLWQLec/5rNVe9GY4iYvf3W4CCGnmuolkYrAs9T9itq69cm2sMlumahw8TJh0K0
YWTkPYMDtARtVan+0GyRKuo1pZQxJcgGRJI04iRC9xAerCdX32yBWymA9qp7HOR+Xl/3BNg+KQv9
ygUxR4ec+bHXe3d6vq+PFm6V9bvYZ6957kkj7zEyXbFv2XQopuQfi42EQ7+eJY5KWWAQnz9tbEKd
DcQwMStaVBaK64Dnhn9Kl+A5BsqhxowZ0LtHay+/qsrYO5rgFEsBrdLNYHBFVZk+ytnJ8YdwCTg2
0MpvH574BeAoq5G/O4dXCZBTag9beZEaAEkpC1+Hx2M3Mo0t1CYfvVythojYvY4T9Rk+ay2NMDFG
7r1knPxE0B5Z9bzTHW8bedX7w8QuuE9QqUXjUi81aRxQ3X0Q3eSJkHKolur7zr3l+tY80V2+/MPd
UcRJ556sP97k0VAOLcXR+AXG/VgKDqDm4hxhYuiJR6JR3OMmG4tuIy1Io5olSqTKOgSXm2SbQQ9g
K7mUA2Y77u5qyk3dzoouUTPz4EcpFmr8k6TYkVYE82k7NkkbwcZPsQeryw3NcSyNa7e51rcL65fH
ZvEgpQ9D+4tuuUcaSppj7Siqa3X89Moh6C2r5DDOHgWFb3EH/5tPQajLh01mYyTFoNR2iJliojqY
BVRubuDtRDQSUtpBO66rlWAuDk9cH6ZhhnraYtQ+z7ifIPMA2pH8w2CFOtDnJO7z7C+seXmO8AuA
aAmFbCZrmRDakHXgG9A+Hyq6lDohkXE5eRlBdH2vteJE8SSVmZNUUfMJjCfu6EmwHbJ+66JrzQIG
6uKw/X8mWR+XoRRRMwX1CjofJV4dIMjQcaGDLkdEl8JvIWLVvGYN/YAVMHiyK1HmV8kFxGe83Zjs
yRhnl2YOXn3rF+NQTl9TnCrquA/KW2kMzR9OqA3ACD+gZdEzTL8/f59WpooyTcWwtIsaW7CHznlP
dJ+wZzDH8g9a4TNVKE/8b+paFX4J+HCWfQVjxX2Gzx6DdXqn9fZwfWDELaPQVQO74U4UDh/nkwi9
cJJiyt7ESReSOtNmrW95xPvKp9XxG7okvffDMgt07MuKGcNqi9LFYgLtE8dyNk4G84uLPTd1v+H7
xQ4bjcM+uZwdaInky0rfg7ugRrCRTjqIeKP+Hpgi/AYaL9qVeE+yGGawrWa3+WnQJWg/ykEL+wbZ
R+hce97Hxz0qiwnTKWVXo8CBd2hoLGt8wEQOASCv0Tfpbz5tXUuN7Ov0sdspoIBvUEW66P68b53m
yYCkNZhBw7lbSeU1Q1mv+RVkvz50wWknTAkYkfkAeJPXwtyCCtbT54QII9JMXHCwsTePSiLqXTH6
h7k4Yq205rMSAZ1uNm+9ZAaBCYqgXAzgVsa5hyLdRVV0Dlhm9VKNgg0FFrnGWoPgezubBtizm31y
DgHPSaAhUn32h7fT3FVMNFLh7fL0boFfHNJSMGzf7TWHBTQWdCqEKJfu4sw3mAUU6N7ZCbQpXHca
JBbeEdME4QZsuYNiiiDc5f4jRNE2keYCn//kd1QDbDsg0fOjWBSg7Ax3QGYuM62TFDuTRq7xX9Zf
RMVi0dzQgiiKirhvEfuuN+WGekpPapifunIN/hEcYLkluQOTekYzRUkJUhHO5QgxXw6WSQYqnJ14
6ljecDERVxD+H3XtqfZCRLlrqvnywlhUGFv+ftI+ZftXddWhBSG5Wk3USTRNJZ8x4ZQwvKaTULX4
l+E0UwroJyb4C5VEDOx0PuqUslwicvBOnkKU9uA8N7BbIOwjtadOnnCgWQS1DcrBJMA88zj8zEOC
xJM+PTrqsW1xMBz8FEfVpezTYoOt9t0Z8G4G01DGl94LxmTmyBAaFk5XKdvbD/sUrkoxnbWNNio5
3qkKW7FSSorHst9guM3v1dK3s/dCMJtMr+NsFxvUwMDa3ysvVhxleBqKgAyx1UCi5ZOmdzedoOY0
U03o8TGlCBs9v9UmDBN8yLm8gyzsAF4KRz2BZFyjN6sivz6l2H3zVHX1Ygg96h4s03D3AQYJckfC
rvuEDCQ37zd3jJ72vM8Q3lf5HLwK3aGLAp1bH9Y6JxXje7PbIuAdMV2AkXlVw/cTEG0wSI6OqKy6
8jVAHyUAbOH7cZgnVkFH2ve2mv2Y8ckvQ2cx5PLFWNDSGb+Q00ILIFXxLtwfXjXSAEdP6ow7isEj
yDMncZFyCQCl5Wa43901LuAbC7YkxNpcIu/UDKhk3Sb06y5Sg1fbLd5EVjrofyzmja6qaH4nnihA
9QH7TYRGGMEtJfbifUBipkmoMyQADycmzwcI+WI2Eb7Rer9+3dibDh8tgzJ3OukRopjKys0WbhRI
+q3TsPbPoM1nguM3jFbQ2cNmJRKhHLpUNa2ftj+9p58dWwzmcXKciHw2m1hhPlKTTXf4qPw3mVPO
Aq6MmzcbtVulf6EFmiiA6V0M6IpxYn2WIbAJITy0nnX9l2sdkP55fcL4LcsnDdjikfBjpeMFjETG
fRmLDlSuOQh7NUYF+cv/8VozdystCDKIW/Dj0LjixZ0Dl/zaw4gkJQMRh4flAEM4oyiXe2D+Q8qU
14NdrFrROX5dhEsxkN9DRUBNwLffv9dsrzFairjwAj5oOrNozf8F/GRyyWMXLJscq1GPS1KOmsxn
KgNCl/ddcsad/qbR9vohvCRl4ThAcStI5d8TZZlmFb6gK2K3AwIMBoDMz8JAwL9JTSpdr3PVabQV
+TkDeZBn0dNXaOxIdG5fF+/o6gGb6ukLE0y5NvXNf0r157MrDkzeX7ARclrIPWrMTmbaugtbMlHE
4Ch5qsxh2sE+JY2JNFp2NtpMoBlkKTRZ02b2LFpDeIil1/4vKbu+7KiT6UfuJQDKXUR7kP6nsmR6
6tB7HwOsqYbRlZcv2XOhYv7WxPrtSTVUY1bt94U21Mnl+Uuz5egeE6VI8Eg9NquT4NHvi7oHjlJI
YMcfY+3dg9ZQoqsW7sKh7YOlxoMn4B0aFCvcuqk1o3kslWVCcCAPNIVjit8CZ/C499J92wLKg8PF
Z+rM7wt3DTrGqB/72Gn200dDxyRll8vSCLjAXLhheXteTy+NvpuDaYrJGswzxFP1EgSssU7J9z+Q
/t0prAaRbKf/JfjIMqG/pHAJWjp9CtnaXmiM+O79I7pN4yPu3dDjXeX7H4stMlGuMJdgtcFLyUrI
6PssjJF6xOw3BNd5M0VWf49YBmHS2Cfrvygs2HjwxSl0Rv3a7FP0bMEpPSw6UQgUkfNFzpRMMjGo
ZqAO7K5v4v4JGQXsvBzzEwJU7XMf+IWAEhUqr77xOd4ucIdrC5tEknZEfxCMDs62MQPpB7lCym3p
Qa5RqqJN/U4TjBDzk0sH9BVUC2cqNGw5JxwYPAf3PIBpb4p9wffAAyqYUzz5Q7GxjELiz7U7Sl0p
iitMABBRTcguFtPbGh8zIbjZSYQYbSdnN8muC5z6eAidHrOXQFACVy4Ekb1VMl48OTRy+xTgAyEG
3PDxoVNhoydZSRXCcNm4U3kUiY6rttsoPNrTra8wg+7AEFrSn1kRyk1a+9TuTULwWSR6inpwu2KK
WYuYeag+wRXc6cBpjcpzYX0+TmivNSD6MA/QBSzrxeNqjpPrC9snpvlFmngh/X1zAFPBjHRdPLPl
7p24LpoqXK1kEsfKud8IJaVrP08HqP6ZhTcCsrqFQMZG4MWRvBsEiDx9kjTsm2+4P+6eEVcC5nAD
M6PMj4U5iDGa1xdty4bbHgVvvfRScH/O5RhpsmzSWRTzUP7DZLX/4+aflN1BpV8pNDjIC/1rYDD5
HtJUOb8UltgZNGAEvQ1KHzvHpC5hgePlstRRJVCHj1cs+mgoEr4BAciurXdezlkkgl5puay7rUVL
OLwzfcOOybX4fOeOm5GUZMCMLQpj35C3CWalcGwuYVr3JYJthEck5z4HJDTp+xwmzCirq+k/rls7
1+D4qKpLGpWxYStRZAmfP76VjZuijcM6zYz6WjmGcrdY/oDT+m7j+8ge5DBbBVX2I5dLeeLllbUJ
XdL43Td+IO+nuaZC8pZkI1N18K1yGlmvgg+8IXuWegptx/cpnlgbaMyXAHnzfC2LNqWC9yuGH3iH
exsP2kpbnknpBvV2qqlcMqQtxGq2gaCePy4ts4NuuewZP/zqC5yadZPrOxzqytJzxIzZAVtuoAv8
ZnU78brCWX5ojZBLAPXpPneqiDf7wwtuY0Y0OOAljAQ/T677778gPbDywHJjuDet+ERTsmuu8ik7
5PovIhhmlwc7l722Yw8g6JkwWbnXMpEbRMMVsmSugQFBbL0M54qv3ctnkQ0GNFZStLtnoZMxxAk5
19lfb7/kvbhSAS8mInigDBt1BcSaBTbClpImbPTmt2MbeTzyeDfPvEILmempdiAd5FtSQ3ZEzqp6
pOB1Yve3vs0KhoHEhb6K3y526Xkdja5NBG51nPZruwy+tGemR3k0DLKS4e8t83dwLUmxsYAfk6fS
rN9bJQ4SpCEDdF4pwKEuK2DecOAJCJtbg3cJVyX72LLYv4WwFdMQ1Ling7YAXcoZ+CTTVgr4g4+b
T1NF62B6cSbaAQ7uhSfGCGNEfUNL2NVB/uOjUIhqCx267fdKZSK3GpXBcm++ez3/RFvgquUMyuvv
oGe71CHFl1ok3w9xaMOZXgiYfwYzTC8pmDYViyi//GTfkFrbsBKd/k7vhkiMygTQI8cIk8PbdPIN
Fuu3P57Gz9AHx4hT0yVGZqlHDg/ShcEclYChrwEDQ/K0tvmYuI8rvVDVYzUWG5ieI+KIBGmg5n3x
wB40XT6m+kFAHju6rnWtYnU0j0/7ub25P/i5d+vQ4YlmLrL9YhFiQvXtTAL7DHb7vy7nR6xfKXLt
xtVplsBktPEMzUil9+eXtpfyClZ9E3lpVNZZ6fg2PCgoNj48rzR+zpns7whV02azrOGMgURZojHK
CcrNH29b0C+Zi1WF86U5Uc6BTa5IcqllROMO18AjSzX0on0KrEr+dDZERlykKVSDbQXlzQddtYt5
+7ib8IfB7RLOuU8amcg0MkrIAkU9/fODYKXpts9DLhgUnekT9YCNWWsCg7DoWix8QRopP6OFGLTV
Pr+8Ut9SdXrnO1CmBQKHYJKC4LVAQ5dhGLkDU9WGEjMf1aLxNvTLfX+nGr/DTf/Nv7RaGdrIr01V
JTaMes6NW0KT/IxNglkflHhRZE8hQKJb96UjJePM9/SId63T3qjNbEK1Pe0GPyWldksaqUc8Tb5S
b5WfIR714rV5pWph84ldngJxoocqsd6MeHRGPl8iCfQRRVsa1nJRX7/SddqxqP7IIZQmEymogBZ4
QW8D1DAfi48LILG+pEnLg5mCClgm2uKbPH7bcpquDc+xaGQMh8B72UYjixazpsYINir+SoYYyKji
fYFyn0nAHVP2V/uRy6OgVwRynCVZRN71pxyRnQBHazCKnVFs7QqVYX4meom62oAb+FgIE++qxa9s
cXvsG65j4nc/rw8Ysb0aeM/AaEKVl5DhSNK1CE3vgjtCZEImF64dcoLqFMXBaIUBu3rBTGf1ZNNJ
ijK2tPmZxUxvyKI+DXJxBESMhDsjWF/Pgtky29jjZ7e21gXPUrcBltjkDUoswZdhMNush76e8nZl
QAJKV7a5mbRxFi44kf+rOrsrSRroUTOjkCoDsh1Vii+inrUrD39Zoa4yfENMJnSwk4UZXzbYhpko
vJBDTC7IUbC52wnqNWCRHXqN7vQTilTkBOHFVRtlDY8ne0xVqEWHJYSWXjKIdHiES973zDD/35OB
K+Ulpysyut1ucdQrmYIY/wggoTBf1sVXS4ct2bzwHx92mECDtfZWxbjr22Zbfa4W4b+5PHyJCvar
ZDajjJwHidyaNGO+qu1+b4xWxoxnZKEQcOyinVXNswoju6Br8d63eldwBd0jnYnOVnBnIbyDVbZE
Vte3IWMzR0tNBuHUcRbMy2dA2+nTbqSM0kM+TAjbcAsvg2gQhIV9Ez0lV1f00i/w1U+KohAsU4hQ
kYxKuSjUc9AZ/4fHJQi3VmeECb2umyxtkgTrZfaF2yOjdaUO1p7/HGGqe+YgljnCEEynS28YDpyn
bzSz5mlRk4coAnT+1Urt9r5tWzdHAg5RW97kEMjtYIIzMK3Ggm6zbEUyVsK4MifrKBHuMDPkxa0n
hmtvLrfTlz1YUmehhcIF/bYZIlbeqYkrNyqbmfNv9oFgVf+kpgeW/v7Kj8O7ltyk2rjYqbhxeKbQ
+f3N5fMEs2UbbjzergruiphNgvB5rGtz2JzmKSjXc49oQim+ndpai4MPqcJ5QmCkXibh0E44GRAz
+WfDtgjVlRPvhS0djoQU3lGKGVIKBvGSqqoRfSCOD+gh2os2Tn5vOPJBHtSw4K8rClhBFSHwVC/3
CI4TNIC6n1vlv4r8KzhZGD/7sJgbq6lEM3NZ/3Y3/yZOH5/uJYsDfOD350+AYZkn5I+mgaW4JbqY
5c9N9kaiF1/PJvnLcyQ3QQkDakvr6x/e5PZp0rlGnAlyD2X3oUbQQ1XlfqxVjOkxrGoc3zFSvZzQ
LmzfOM4sD+DcHphOur1qrwWeU8wCd3nb9z3nZbx7rO7CEsN5pjD/ED3zFmO4Do9kcBxXcClH5Woa
t3DTMcS/YaJXINPsvLMEKO9M55s2fwz8lc8MtVBSayTwSJ2RZe9MuFWNGRvA574y/B2IxmzfrxqW
k13UhGfyHjuVvVvUdaOLyoTNcCDVnQPn16EUf9aD/vbdQsBrLDwq0FsuK6VaCgqkXPUZI8b3pgU2
7N3t866x6r3e5YZjvJay4Fy1VH0O91K+6UVhHMVE/Jz5DJWtGRklHx7GQR2iXttb9EVWeXRuP8UP
p8S9LAYiFsuIr2FuTcBCM4F+uqM51E60AUXSBO6gPweSWDGfrwoyvqVRBFsTHf0onrZkrEQ5Q+wH
TFwR2MON8yvwaWRmbE9olnvuxzr7iJ6QZmsJBUSiSQL1D6lR1CirBsey2FjNiGA3hnl2b0Ayz4MM
Yxygdwe7JuPwhvVSt000Jc1PeGc0NyBaIz1vSynpotsv1dSWjRnt54pwsDauESeTlpRLqEuWw8vn
97tVUirGc/sgtp5LzBLJFO9Vv8Lz3nwfiE4aqWbgWSFGua41AoYY6gOBL/H94M/nS45+U40ujv2L
srC3KeCtGdc0tQC+xbmyFDgsVirN+ENroLBN+dHg1/ExlxuWdAAoXP3IkGGx7qaQvt7W0c4KsQF0
2AIn0XQX86y0/Fk01uzuCGV+8gRK3Ldbh1rEilh6iyHLXbLXtKtRokJ7j5t+Q7aLtUfAnbS4unSZ
82YH4Lw0+R7Sy06kD/1V+iFPi1xRXSb0p34A15d4xz5xeNOloA1bZDtwf2/Qz8bXgIWIVExJGlzn
C20Q3WfsRgMhLguu7iprjhcj/5jvX4N48y4fy9nEkuRM7p8n9sHQFGgbIakdK08EboQn9JjM9stG
Oo/Ws1eWVNUNPPdCG6x0hHF1WwmdIOOhpIFerk7SOdNDy7OVGwGKzscMEqP7FildIjoIFp+MQP9l
O5SxibCWowdFUED5evv0GWTQOX31tGFgw3RUsp15FMX9JE+CUivfB3+vTASK1T+KULpCy/wJ8kmB
jiJ861prBiZ5guVI/JfiM4y6GKW+ZR5uSdVeuclkHUn1ytBTEe0JWKQd5aNmb0Es2kvX5jghUIuY
qo8CERexr64o+I0fbdGuLPXR+/HTkBmJ9qsiuctiRI1OE9E7nFvMKZlX872OErNeAgxtTy12umOs
NB7TsHaU3II3nR8A6P8KxyNTXptU3AI2XayxW8iORKskyrz1HgHyFV5ElhWtr72d3AcLHKRLptY+
g1YLymRJxFvhSltGkEd4EynHenj/yiPJYWg7Xkk9OyOR6SxUZ98tH+uAIQs9OuI4izByw+HFyPKO
Rd/YB5Chu5dUcse28kMGJnWr8SbBXzrG6x7aE1t7RbjmCFChy7xlEJQhYZeMsBGGZY1SN7Kj/Nn/
LXEsUiyGlXUhaTlnalYSUNvlR8yQpEoUAIAsFQtMvkf1QGaNUtJkP8b3vlZJ5FAmOXWDdKcMYNXQ
je3irjot/Gtmfc7iszEXF6qRXHFwm7RMRDWjbUTStpTTFKmkM8Ap3/079UiSc7fcT2F/IOiLV5ow
r10SJXirrkA4j0YupF0hYHIpSawu8+WF/ZapR4nHoeTFIoXBWNCvGz8WM+4+RMu9/8Ych0QSKh06
eDIGr48XYKwG97HZFgVfN10mME2Tzttyl3rZ8xCV8P3+HhsBwJ9/OFMHRm8RuD21ic0asNNg+DL6
xa049xUVladKxZIyfmQHKzH02fILQckbnBsmvkndOxU/PUddgiaQLw+HdaWWKtyOpMRRWkVg42ev
R6fqsWuQc28J81U4Dz7Hh+jKJFKyAse7nalzftrxf4kzWLKce2yWtyO+CFjD7OlccFaOwSr8w6Wd
Pm3RciqpPz2RSbjlfLVO/iN2wEx7iWbSr3U6xqTC6YhrSViXYrPI41Cet01cceuqt2fA6Bm9i6o+
/MuGiTjoF138wn37A7/zWR1S5UTBk23py3kw+M34G2lZE5Ug3GrAnDgTTjaCn7CEy+UZvY+kf4aU
oqD8mpvv/E/kHJBNSQne3q5NzJLiQzkGl3uFVWjAP5OsmbaQ5ttWz4yYvj0C6qNo13ry6zQaw0mW
nnnu1ZLoPCQdid/ylz79+CVC3r2FJ3WidqbazQiSRa0hUtJ9hK8sTW3/voDWCv2jbEwh5T1/09nK
cjyNE8OFF5QFMRWYDoeIUvjToL5RqXeUMmNAm2gFHYc/UVbInh9JPFNyGH5tHsYl21ojSfQeJrY4
BBBjwGopgFqvWqdwxY8nSgFrRg7TAeI4xbHCiPunTLtXrXq90HJ4CkbbaIsLWKTs8QIXQwtbQz5P
rKfw/5cp6K13e6Z9e1hUbkFcvARxrD7VaYmuuhONaKXjQ4miu4PQKlNux8N50qBA86uZjlymnatg
GC4+Ap8fgDRj1zkcFI4I750qTvvbKxw8XQ4VtwBRgS7eQdOyUNO92/tW0iV6AhkbpVh/8tYdRYXz
BsPbFB9XSNCE6EofY4RYLcwiyXqwOeZUtgQN2SXemCC/FiFlTZTpVHtxx6mIOmlyapiy4VDtzyPr
Kuqic9fm7Y0xvG3flSrWkO+RqBKj0XjEFqs/l9XX/xiXfCSGPMgHR2eDYao89JeaoVTvQIFEUpxA
A/bIcTvptwaY+5/vO8o+waHj8VSwij2ZkNqaP75IS008JMrR3UnZ1Ll11cBsHHAyse7gBnidc0ZA
F38g/MWvwBtySepnGJ6nc2PT3HBrKI7pORqdVKLblftWJsfezzr4nDFb3Dbj0yKiQIE/HcMk0xqG
EDGb8Djofm6XyG5SHgfXdROkWqCTsvIk2wsdZoRKwLEF/SAifXHurRC7bKRPNwGysfWYmdC39oXk
eIICf3caL5tque0cGUI6a+LgSgFyM+0L5Lo3TUJ7PxMhw7dfIxBSk+WM47+a2qHUr3ORDacrUicQ
VO+URAi7ktxUdw53xGPWus4GnibDBTE3naXIgaaEzh6OupRCx2mFmCCQ9OWsTkI3sS/GvVauUXwu
jo4SMFvUXdpXDeEKAZLFX/x6JVCcwT/k83amMNtuSU3Uc1zf61/UlQTdO8+Ij6aohMo+Nhx3lYBt
Ln9TrHrSWI+a9S6BRYVyiBcZ8++2QNTet8kYI+z4ASYTI11OaEIn0EZpU004XmsXTOXSsX+IfNU8
F5iU8q9wQseErF0fOj2ZVV2waGoe1nj7qiQxFayMJWyJzpIJ2CXgKtCqo6wJtD/FqQiSwrjDW9mK
sPCKlq4G+UZPIN4VDjX34WdAfcrkQwxub/GXyWanL61mrokl36uwXX1A5kxluXeygZeHRnB4gL2u
viXCisfjZyW9kRWr/bV0vWF5ab6XmRVB2tXDTC4pP69+MtcFiCoIA+rg8VJgxzhKbIgu6YcIlgwf
Yn7H7zEdNM2HQaPVnJQv0IbQSSHyaj8Tw9w3WNRPS/qBJXhOPV6MIuxkol0GfaQ/FamWOU+GCLpU
71XiuesvlFncYuyCeQL5AValsdqMwfz3SM0B97gLs7wwoygm6T93SMA3573EJVWNaQDZPJHWedCb
HluD/GAy8L59ifmcB2819vK0S+LUxFrvkg6WCirEMS87JSDHo0EIQ82sxFMP5AysW6P4FpbCKj4h
aD8WtOe6eP53hG/mfsQAwgYdMoBwMzQoZIgm5aXGamUFvjbf8FsYz9hExoUAxs3mYCPAfj6gKlN2
NzFeS0bU9/iutkp3ij4gbXhntBX2PaQd5QOd4aDZyIAYbYby3GKE1WiMnDDB86sHUZ9F/SsBWdW+
rFs0OXkinKU1GJMC3r7Cb7oru6JK3PztUlBul4BUmy4wgX9w8xnPKD7gKne9lSOD85rA2qUboO2G
JHIheU43ddw/qbsovo4zIzGg1RIRceTJhFxlPynODByoHHtDGRTLbSl4oX8sm07ksk9qP8wAmGaY
UtrFEetfS2UXET4FR9KAZ3lvwEnhI6Hb5J/ki37ZziS/tGODziuEN9+gtclRnJTTdUinrD/Oq7jM
f6tUTqyIIquoJtnhrVREzF0emsGPLicFnIoxMbpUtVbm4gxsECS44aPaRLoqrX1HO+aBU+n6r58m
hXBlI63zzulJJbLSuCebiRZOXp0Jex5qNWcDpBxQIv3CX0GYRGwY5e6bSWAyxZaTFQl6GwPMbSqk
oJZQFKrONaxtr8Atnc0Dwn6j/8keneTTdHo0C/rnxHNFlpoCR8qXK5ebdqtwT8JNdt8myo1SEjxL
EX0Y1r/coiuSR8O+bHnP+vrNjWq6ZRrHZGxws/4GAZJPk4L6C50Khuwxc/CRMszp/jREpOgL1EIl
+mSsW2yB5Z17AIZU/n2q9yhu61/XdECpPNNhge3/XStj8CKaL2Q291tIDODn44prheTBlSXOy3uY
bZr5ToF096i5tdOrgp055czr6rEWKZpuoKOttjt8QwyYktUaSHJ6yq5IMWQzkSTIyRTGpbt8zYdP
DcwYLXio/w4DLmDUM+kjxljhl3no5o/4aoJ+i9dEmrrPXQff1kp/22M2H4a3Vs0xzDoYq0cNU3Bl
3uVKP8LaIO+5JF0cQs/c5QbWoMZjt2RrxxpAGmpUFbb8GrsvVDyPvsH1GcM1UMUR+xrpdnOw+OuX
5jiJP622EmIfmDhZfM7+550jjyrz7tLiY4LowiAMQ54nrXEacwN/+zNXla0e32W38qAyKw4T1q9/
hpc34zFmShh1+JiZtM8LZBdUrMJTo/tCSyd4tuXJKw9iXIN4D7f+iYNl2xiMQUWZUXqKYLVo8wuk
BxJpd07STXxSb+iUZAxnaaUOwqepYNsf7Na24kHfV600X/p8ldkusAHCTA04GaqJUZInEEtEkD2Y
J7VUjKbkfbW0LPl8gXmzeh188rrytyCNrzJBppvu4Tn89G47xTLlQkqaKOZJJlVg58NYge/GRQ8A
o2T89AGJ7pjVANH6HQedutGJUZX0/LFqju4yhYHKzxmJwh6akPGsjLY0dZRpLu21WWPmC9ChIPqL
VQhVQRNTuXGsmFYnWHgVFC7MhVMobRoXjgS7DjNngJztFfgnE+11vW2MEds0JKmgyZMYwSx8Ferq
0HJ184+lW1GKHwr9RmUFEmKo+7FSUnc7QaS1GxlyWk8yVlbQ1yy87J7GU0jx1UwQs2/Feqb3Dufj
UsW7GUErBZpm9UaAfcxoisYfCQPxP2I5nxxS6y47HZrOYlCcdjXwP/JMseen87fp5TGTfzdM442/
TNZeB8eJ8gqisPAJwUI3fKk8T+i2jVAAFMMwDaZcb4mAlvvzHWdy/YcVlAK4tCM8gnEsIdVVuQ0r
4Cqk43+8fkxiEXDzGXuaqPfW3sStdvlPf1Wxqve8i+mwdJYtZkJXQHWSmSX2vbWcn+URPPg5OyJ5
4WBKAl4YiNkCYqq2W6VA+YDITZoDTfDpqi1Cvg3NJDwB+Au7BsCG11aWQWxfO55LTr6WPrFWxYCt
1T3yirn4FMwmdyjX3SB8CdhQNDkEhVCK9WI+vsJ5Pl1IffprZhNB3B2TjyNyi+eT5gU8R3301Co7
X6epTqgg3WSytssaVGsAj6WHzqH+VEF2TH0KjyxjG7BeNvy8+5sm6RW2NBT0u2gjIxor8HkhPVy/
ofmc/u/+Xd0HE6CQTTv33gTDLKmdOTHZx3jlmn9pw0bvUYJgtOURwlat4xn85bw0XQX9rHctqRhl
RImwl9zI+i3WShi1uf75z7q+xL/bvRyXIk8QjAnpbOvXZtjlciBoJcqTpgvN47ksRTCP19706S5V
D6k1UElPuqkkU58/JGi5rhIKyk2iyhK7oCrkk54dlFO/SAj2fFloPYJIJymGZ7F2MrgcOM8L7QjC
2voVBnvS68w4GxJCLLlPxtD/SUUUXZRGUqEjcCBqxAFZvP+eN6WLwqIYiFd/onx5jQavTc6f+0ep
zpstqAaXcqbzHafbHTd/v1wEGqzybSesddyDd4DY44nmxGsGPwCzU9h+Mq0dl6xFwzyeAqIeh2tz
Dc0S1jrurXAc9oZCcgz8gS5P0U1gPAA+AonuBfC4xXu0YQwhL00mMomSmubftY1ILQZ6Nr5Fipkd
gXbp6SV+BZjYRPcnkh+Ub2eJcuozkCyZVWyhWbl7Ixo8ETT9O6hXhpRtASxQ7wnFa6aaUrmaDNd7
yvsFKEtOX4Dr2R7RYKDQ5CBCv744TvxnMx6hUIU1hbhjiuPddrw0w6lwXhxUfQeL6/Njhv5K19Xg
JeppA7vrnvGgqepF1twQPu25S4VwhV9Lo/Fz4J7RXOLj8iemLXTF6CVKxnJ7Z5+0SI91IVjX5EuN
46RqGuEEHBGurE/X6gxxSOTacGwQ6XffGuIYo4depi1FHiAUZ8J4M/+PKBEo4fYkSKcCTBbptEWd
L8LSlXGv/n15ALt9nXvO4e5kxEMdpEraWsY+Wcs8sfoE4lBTv6Tvms3jC00Ef1ijbJD4uomWnOxl
wwCL2hA54wGuRJmBZVLxcGVIYCE8gaKWOCvFzuHVzOqi61z7Nw5VmnMDpTKpFunhu3/UhVTLpSs4
SVipbGu7HdbG2dqKLHJSiVsOYpWp/2d1nJcXQlyz/WRSVt/EvlPjDV8JfCKu774OzWGNLlqpjIrS
TZPJk6oZVxmNkImWflNoGfSHstwi30GTfUaufh3HfT7d1FKLypJ4e/xmuMWEz7/2LF/OUHuZnaXI
bYzDqcSBcy4UcmlUarpgNvB/iLa6/KSQWruWe6Efc8tMSrVIRCqrCsHpKZQmEir4uHoQh8jCrZ2c
XbOJHl9jBpxMzEt2iI9h14GXrgFUQKQKNT62A1hRBwtuLlvzInkfil2hxHalHOGKjyL54tYTVMw/
10VjsFQwsg9EEtif8Dewaz9Re1T4qpRezz3JnZB+TovhaVCZ9BRQp/P5cdzmOOdkugn/PFQ7SFW+
2LaGil6Knpsi6da4PQsEo9dsrX1R0xrZTmS8Y2ZKzRz2DldPRhUf1D2EZsevpPrkNsPwyk4kCLkK
1RSJ2/GVERFxHTz6SW/SadzvNvG3uHQrqiYR8IjiSzzqxjcDMdfNtukU6zqGPKYiuGvRtFFa4uhz
n6Cn+SDq0zgH/nT6ENsJ+swgpbt5g4XdF+MoP0+T5u4FL5HjFD24NaTNVQn/ViQ47oRoSb0gvZ/M
t/2hPKbbwWlLRrzOSzDxYVnnQ2SawXHGgaGWZpNhvthEVZI5BTFk15+kRIbXq2TdtyWzOzEL4P/F
PZtbPk7cokx2GbubTyhGXWxyULsZoVvKDgDc+lIDtQPoIUOIVE6tzT4NK60QfnlzKReyOfFPX1Cr
HUpR2xPdvigD7Qa/I0Asrw35iHfC486r3sSVzpqKImobGOm+iqCpf84iz0bCbhSTPoVGvdtEVyWH
XJvogQwkmULdoU4VumZNu3AHT8dNOZ1Ga0eHTGepl3wVbYIs/zlWkX+8HBqlvRh9CaqCY6BwIJUg
yDfJHGZ7KG51GFp+/gHaDJATfopbgYCtAo9bcSHm7MuNbm7zPyqmIoAWX6aoBbEgX95sVIBIDXY1
V81Mm3yEsJHlYfPPzV+rj96TNZIon35SFQAC4XZ3FA/GQXYTMYPo1PRX+Cqe25+aF3ytLe5MbYIE
/K7zDAUHW3IApxoBsPeKJnlkylTlsfQYkZ2OV+yxfkjxozP6577SAuYgNTeWyBZ13UMydK42pfHB
oVOhJ+3CdPy/E815iD0o+EnorlEyqXV0Br583KfmTsVN64OHsWKWDqVQgvtbHCtmZJV9kHKjPwfR
CNpfithazTqENT7IqnuVS7EDXTDjf0TwiiZ7wurDYppC69V+zfhYmt+TC8qTeetoHwql7K+wN9Lw
6e5MS9Xq9Erbbwai2Zu5sTe543iJwqjscgr3PXdedc9XAe6+sfZItbSNnWTcon6156USgr87DLpn
onal+BIMlnXJ2JMOe9jrEyWFfwRBPpgxgd1Ip2w3q3s52b3R1SxdW6NCt8ktdMWV+k+5fDt8o8TD
8MhEEmP/6leQIau3AtSKM2lXY/kiyjTJXX7JJB0ICWLaxVCFc1vP9cFKs8G3lI5JcI+lzFKaWqas
YUFp7qdyTu7OdK3lsLnzCBgC7D4us1gtW9wY4fMrmrcldcfVt2Nh/LKkGaScDdk1VIkCXAYwbNrj
fw5wOB9/q8+xHC2jAUM38vlW1AjIZG0+mf4GvC0frv04Q0ijYjsqmDWUFdVcNyhUGJWobeeAjhOt
8SD6KVeP5uh3yg3DRG+wYkgQftxgpGAKRrjkHlLQ5e7Pi7uPObkV0oBn8jLiv7zMnuF07PBjxZNd
k/iKpp2qRs9Wqf61Z/GMaVrVI3WZ62c3RDM4cp3/KRk4GUAsaRp0qkqOVPUxz8pZOpUowDAS0s+Y
uCc3UjwuvwxsgJMq1aZuz9nLwHQJ122PzRuzjTES9ETC3YrLPcmoWIq8eiq3zA83Uzcrj/XiJ0FR
9jI15ykRf38Y+TvY/K0383CBWkwBkYewg6hoFXUBNxNHcwTAXIeVDHyK6h/fAXE57oyLVPvkkfka
BTALyecbilGTtupiN9ePli0guAV+g8NXxpufCiqQUXcUN4erbwPfzxqjPNe86siHzbAKBy/7jWT8
r8tvOuMiRPEMmXWZRi4Ud/7suehSzK+DL65RdglozmrCULmlTEHeSX2p4KJyO/DxKy4/OE+w4Wu5
4/pTYplnvrD6AbxcSTAhtRQa0y0ql1M309ip6nuI2d9Q/k1z28CLveDwq8S9rQiLXBIV0cRQsHaK
DDU4dJ7kvUao3pjpXjQHV7onKhJWK2x3ONXZtr1g2J6dRzw13vy9JnjTaOX3fQ8GU7U8diROUKgH
xcglebQx0LGS7xVYsuKJseedp4EdTl2o8g99jV9kYSoKgzGfUc+BbCMI/dbVkWJAbQ+dDEEU3IkG
GftURupJNOqn9hG+IOsjBGpCSb7UOrTzaltqvWwE8vk+79i0WXkWVCy8f7NnMAButUb+r+eLT2M2
F75LK4DnuSezqps8rORyRWM/8BHhJ2tU4e8iSCN333VigNdUb1XkXz7PqLr0AZFJUNrVCJH/T1HN
ICJQNmvIGuGG9asKRvhpzspDt0N29qQy3mT032Hy2cYE/2z3T9UWz1GlXJyd6VlPkExc6EIWeiEw
b9LFBwdHrNV45Z/cGsdoBbxM+6StnSO2KVFPxJiEQ1QyitWApV81lThsNu3ICFO/OH8ulUPP3WYS
edMH8UdUK8/u7/5TfOXtRCgLWlu4BB4oG+KaU3D7CQXiSjM77JfoGLoXXs9pL/+wrVpJaCY4EzUo
mlrpcZ6K+x4Ac5N9QGzJDTvhouQWvrNsbRpGafLpE+uC/UgOsaNje1yf8LqnINCCRa7ULc6ro3VJ
BAa+164NDhxy0Bi8yg6q8ApCVwyj3mMyFv4V1Hhxq+fDeiKWJEsq3/MUAhcsAaD1hPCsi5Tu1wQS
XKyBzzebVEFXwTUOcfh/76OwCP420V1T2HCUoA74Ql4mJyE/450/QJjbGpkGsEPLaOFgrpU5Qv9I
ipXmZa5RL8/an6vlKJg3gcT0KFXqzoyY56aP3qyooFw6t7LUp8IM4hj892jLba8DBjLf0ktAxEjX
Od0x39onuWFJNUdj2xsYs5/0UsStXTmQ8A3b1hr7lDH1uChLZzpdksq5JyLXAkrW+JWpsbmzbmKR
nmchNakvE3/nYg7RwntVgcP6GRkkpTL3Yq0ANhp7b+G5HDnhoR8jS+y4w4yypj0Vsc5stZdMim9I
N6Z6KTZcqfRG3fgkn++HN5z8z09wiK847mNlZDWsKEXKzjYi4ZQEbHe3wtX/yZTyIwL9Hi0dwivP
VpLOYHdwg/J9oBv1zVAASc6/xN/4JWvSX2hgPcZCne35eJRvcgZYt+2D7WkyrvEx+jTLlIQ6nZ4s
mOuOTDrzvGSDH0OeMIO1OLmmPear9GwAhoawK+6S0un7mUQYAkDSiGh1/nbO9bn9CNWJFukSRYbb
+1NJprkTPcSMHsjdJAHOf9dJEDbpSkTRJcp+DdnMYDPo4BZmdKR35YzDslbuQAY9A0vFn+iarcM9
8gPE/mW0um0LEqR5yCOaBROMl599zWucKAuD5XQFEYdQZTA4rxmPS1SAXKWUuorHQu+VGvCcyQEx
ZkpHpx+bldwicNzGP+H/WkqWK4PeOSApjx74o/IhsPR+OWULnqxP8DUc7y+ErRux0WF+nb1SP2bh
NCvgUoLBAa/AshPHDeNDZPH6VoIgE7Wjuzg7jISxsIoBGRQviJ+hlt7DhhTz7eIzPU0eRw2UcQHX
kWInZdyQh1DawsbcrzYg/JoBQj6L3xG+SYQr29sieqxM5Fcz7m9Nio8Te4eDi9teCCoNbTm/VWNO
gTmBBAflqf4UCt8rnDLmRgeT7wVT1S8za7U2HSs7NWSgEyZDZg9oflGAvi4nI8J7KKAobBjZS+ni
od4cF8r3g83GnyAGNvuutYYBBhBzBgVb+3HUQZGFBjmAVkCqcBJBJ5EVv0w7Irh8FdKGGD/o3upo
1J00PjKF2Y10pzKtRv/fIzd7VUThg6F934lBjWdXZnXhRUVOZAVXUUex+Tx46PBnAibIDMyG4T1/
+I/BzQ9UhNWyc8y7GzsOKCKjSuabmxuvB5biXr2MUXKky1KhMBQOQ4l91rodCChflOcQEQan4G27
HAKc+LkLevVidcd9rq+6oZXUbBQn5+DbKKWp4aMhzaLD6EUlohTpcMmisrSEcmXn2+aluExsq7EZ
jqvX+WB67DkJyOA9Jh6u6r+0InuEnMg+hDh63Txcl1w3yo+OUWLijSMrw0IQRMCjpYRpluxBAAct
Wcrh3hzQrfrfUIKlD0g7N6TrCWqIDaarLReA8hr5tgF7nBsV8apW8FsLJ8CRBL7HMoSuh14+TIQu
KyfmxxjZV5ErBi4qLaT382h1zBRVjEUHhumFXsI/HL4RgaE6orlZYdjLI08mVFR75zQlyX4klgCT
9t/pXoGgMPAhoSVBNbILUCTlnt3NK9awGI1decMepxQCjwo28zjOTRZNTVWhpH2p0XlogkMbuckv
DpfTVQrzetA8QTbVHQw9jZIoOrw1NcOZecUXVr9ZwrkXhFS9AH4uHSsvn4y1EM65+gtPS5Sc9W1e
aqVKycYF0mnNc3nkZAguwu7Xf5LkdSx4fZAPDLibLfcGtm/sdqBKxH+bf8c0hrptrT9nVjr3Dk5s
0gM5b4Scg3UKV+lVk7MJr4tuI+/zKY6pnq+9EQERx/PUBUmYtHJt+Ho3cFOG6r1KNvjtGjmHQFa7
iutY/R5lxEn5HXf70Vg5agHxWqbUK2YWxBPnO1Cfatp1LmxQUxD3bMafKYpIVZZxQuN0lD+YPOiK
jlorSOpveMQYrzU4elOBvXNewt8YQlDVrIW7e7wRLV5JdwXGQzUg+YJNZI6EFZPUm+qfFZc+W/EH
RzLwsCEuv0QF2z6VSw2rR2yiIjVauM0+42n0whjMvb2QUe7Z6ZoliSQoP/SUXRH2pQFFSkgTskth
+RX2dZvnryN19MISop3BWG3FcQEdrr9nyzoFN2dbl82fOPQ+AIpkH0pdRtOuPcGOju+HdJeeteNN
KV2ohLOE5omez5rBsGzzTh4yD/WcAkRiO0RDvJvD+K02foWgwTTJApWkueRzDEmbqFwHKtI1VVjo
D3RuUE5+EY78TIMy9l2EpfYEgfJ/LdbmA7b1tKOog6JlLj1MUY1eWKLTwD226c2bwvTAhBFCyiVz
TOF2cY+Oh4V009rr5kj6OTj6VeqN1/sDPLZSLLo+LlD6mJJK9ksd3e+QSBDee/vZF8CHs2mI8FaD
rNBLP1cqrd9Toza7IQavXrjCes3NnP+/OyuA8ZIdqFbNguuqZZPn3uMy1CJHBRrpgo/VswPz+Wkx
4J/7nyuBc8b9tgWfXthna+Mpk4dpRjDcUALF8WCVkRlq5LtEtJ2Tbk5YOIVHs83W606AxYfGGjPO
3EFT8QqVPxZLLNPZrd1CGiQypT5B4YDxSYFeiS1kjijxPkEYrbzXpAdQGGmsiBVLzd+c6QTWdt0R
ZsdhX4UhMiJH5J6AxV7B4D+Op08+8oYgyb1zKV9YUAlxHtLgpxwfP4wlD0Pe+ANO0Klu2zpB/DaL
yxGSWp5/qKx/JDHu8+/aBpCL+0vvCZdaVC/POoUD+oiR1G2AGEV+rMCRdUJaM6s4X3QuA8xuXILb
vcN5hszPpIen6fyw6C8ssot2zYQmxXle8e4NOzYAMsPQy74nuYk3eVufW7yIZ6ZxIi2oMqA96p6+
jS4pbgHHRtfGAVOHR0+z3U+7IMZJjMXxkveTnwcWId/IttJSNGPa3mKO7u2xg75AwEQc8s8rf/+U
uX2ebwW1QRBM1lco3q9YSNCoOlhb7NZT4rev/CYSAS+pwXR+IKUo/9oTS7R5/7uFbnH2X+9BBBja
XGO4UyANUyczkAoL+2Nz+O2Jvhl7rTW4zT/C1OdRawOC+v4yVSjvuZK5NxMSypyP4VlfDfzw5/yd
kJl9UfZaBnHnTF5+9kjocFCLo5anHjlMsuoIX04xxymWzXKbCPDZOB7MpL9S0zfhXR8kiHlUi3xn
KJWh44GOm3qVVtJD0Piog2n6HwNA1T4v8gN47vywEWMtsEUOU7i8KdwOf/GA353HO5Nnqtn5g3zs
4U783kjC1X6/Xt2/KfYCK2Ba0o9XXG43O48BtlLsOMMZZ3a/ujXB0ZLmD8dawxDSg4yGKg/r70gs
Gxy1ye+aih+zKeXLoTwU8CLMdFcI9j8HnLT/+gkzZO1FfNRvGfAwYlkQHsCDADXcPPu4MUKcSJeQ
BKG1TcTdELZHpkc8MtJzjJr51Gw8zU1JYR4dblU0KBXarpOh2t5KApzMZ+exSjCktF31XomEKSzP
eIxs0rFhJRhrdckTcqk08gC+8gu6+dT2RehM60yzG3B3CL78VAVdsG4pHUA3SyOfhgNkXqS1tLsU
fbbS6jnrqUBCDD7cQPpOhyBupQHwgLf7OOCC4wSxt7XCELy/fel2kwpqURebb84F/qIPhxyYiSUl
GinB5eAlM6p5vfT/uAgYXbi7n92mJKfbBeSbbfSGikCUJkjl/LnWgNBtdBfEXTkxlNJY34IikRw8
zJ3lRxPGBkfKhKt1tRIOqo1AmsCPOf/Ogiclt/BFIWxhvoeCPsv1BQo4C7kV+chzVzvvAKecl0k0
b46YoOL3bahDtYsZtfzy//rByceYphDBZPYrcrawK9ZAbAW6iKU+hYABPiZVrvx0dKgpcryZ657/
l5Kr/WprDmK29xgbwG/xtUJgG7/cYLZnME1sbkv3+mvWMCTxdvNOYWoqlvasOoEy0CYYgXer69VY
8RHY5CuNl+/eAODb8co70zmMsI0vmqCqgA+/9EDBMoEqgLnwH9rttjbQxcXTaIjVo34xallc6GxN
SuyjmNS5YAtq1R58gfK6tliJNErTdI1smM3hrdYamxSDivHCCHlMCGoXAtWDEaMDvjyG/AaoMwcs
qNKwxpx7yhUqK0hWxffHlXrZKCz8f5Bph33FQdvd5TvqKSKFCzsIPRitxLIk535pYnNtymRsqkbn
op2ZcGQiD6Nk2Mp7aKFfKbg08r39elpr1Q6cNHFDJLO1qjbyZnDII1S8EfhnDT66qodHHfFT2yoE
vpsa8+ZjrA0OWLgXJpmReZUbkVXoIT/9buIclR6cNSc7yQxC6rssyityYahwr4OWuGoIqBnEzK6Z
5uB1ErGu7EW02rbzOrMgo9CJ9+TETHkjObc/y+KGClCaxfWQE4oICdi89/EeZ95WFL+n6ti8QPK9
t0H7w0qRq3bKyvMdVV32t//70LRY6OmRaRbuFQLxOpVhVNe6skR5zTrZsOYYe2lLYNJiXDMxmJ9h
KHXtFEMDFAMB/nNu0LCtxgJ4Dkunu/KWHldG66A0t9IpFWoryWnpgV5S2Ldqz0f2yPRZmouQc4dB
UFmnvmJDbYAMUUv8jP2NdZc1xEv2x3Bbox1Jp8/PILYJbz7c/DSd2adcNFiPJjLSALJmgM29c2Rd
yoOJKYAyx/GAhAJa4LMLr2EbmvBiZZEPZPHI+7QCoSJTB8Vyx14S7mMQnffwe1u1no88cCJwMQrV
TvVZ+kIFhYQMBAK6IleLwV6DRk0ttH6FOCywhj3wgu49xM10sSh9BcUXPtiB+vkdLmmTtzDKOEO1
EwlhbDCrU3rL3iuvtr3lbOUdAH8LQtbtkob3uJdeF9JVvDTeZ2AZr/6T/Os0D2cXlyZK4WQFUVXF
YjInyCk5ziMj4/kqfknQrZXIYFnooWV4tS60jJTZH8YJ0TYUhpxwkJQEFKHNvXdBz+viVSo1eMea
KbYBNoZt+2AOzDk/R0mGhiHmvNSe+kgGofFszZsS61XcilRRjpS0PBaTstWwbERVTGICzOXJmF1S
vg8493aaoEz0dVB5Vsv/Ag8cH9Bx9Lm17w3er96pFTgnsglFQiqiwg1bXkADamBk5WKU2z79gL9m
dYjCmWhMUYtpTgsFiAuPS2PABYj/MVFEkeNI7AXk3T4TewmJU8vMLS8IhZ1Ve8VwltYQW+ftmQ5F
UpjpejkMbZbhU8p6DVKcVf3ZNY5LZW5ReSILHAaSC6cmmeC5Fvwwnne8UWelXzZ85DpOrM1x8kJW
lMOM9Bqdl3O04IF66oDNYybrblGsMekVk05ue9MjT/8UWeErM1AjXQOObtYmZHOUn8MzfmjlhG7U
+PbOa5ZEYnoAHIxhIsr4qX5WK1Rzaz3SLJ1FBbyTC1WJgZDF4Z8nWXIDY0GiAuKQ//2jvMoZVfNP
evuzUDuSaHPu7dvrp9k3FFJTKOUvFSZlwpbZ7YnYPIJZwPqTVsPfUV5kacb0EZIg39HjyhgU3Jtv
LjwhHrtf/LipsH2iUQzu2D67Xa6CY3+a7iqbECeVUfNWbrBZRy8rAMjpneFv/KVd4Mcop1+hHBVb
LWMmWJ5F5sKv3YQfgTDC2fCoAgl7+Hq7j5aCanoM0KeKvf+rW5UMp3gHnXDZ36hNNsvKbiwSyzg/
QvOO0P+AU/ReKin2vCyLi81k1p7j4TfP+X01pDiaTY+B5gjHPi+WL0G/xTI6BCZ/I3+7Hp0UuwO9
SmEURggokl1tVKg5/LuOS9HFW1L2PlZy7oKo9AeOuaX7viiCZz3YaSeV/kRq/ppq7Ja4zP2lbaxI
tzKbsMJYgDsLb8RBu1EzJ2Wi6VaRR9Fhnq16A5H/UNLzxH1vVxGDgPwl9bBBMyyrGqAyIbRwg+Q2
sRFkMueoJS8rB/0LvioM1Z+TXQuNlCDPwQ/6ZCR3neT7X0f02Klk595J9cpenzOXUK7hMi3cLM5D
2UDh0bP77oxaEOdgIZiIcDf95qggrjUTmV3jnqzHsTaot5j80Gn3LO/bSjv6ug057QXYqxXYZMIr
XGcyRf+l5bYTUw48kiAdA3yfuSxm8DUGMoyPQYtGNwec/uAc5T4uJVIsff2xTuZblfNA9J5CvsI8
/+lCWVIxvcP4WbEGwv88GsRkDKSWAaObnG2Wd0En1kRyQCbB9BtfhP68Mg6L/RUOMuyBBizFrvPR
I0bu4dshZ1JvKMglwnhAzzKQwo8VLucnWDsSGInKr8A1XJ8h0pfs9h7hek92pYLwYmETj4dWW3Zk
CSkM0Eh1wkCVn2ay8a0/kVNyvFiB/gsqHdQYWe5C0cMi2gPFOpEbtyKMjdBO+TSWlTfSD64GUowy
eajnyJpnS3QS4ZT/7WpXnGyfKrwvRh5/s0fDKUADpDxTgXj2587VKwYnx8Z1DV4Vd3I6vU1L2j37
0xqxInmYbkP+dNWor2qGtNE7NbSx5G5YTFTY5zsl9+gMiRw+rsDduxkwKmyNJI5tWERKuCvgF4nW
T9eMFOOT7yBRMJbyRgkBLBqeM2+mCGWhxDimFz2G3mIV4iqHfPXqD/aVSWFchiNZXUdvzlDWqQXA
K5tBedg1clzRHUITbOzSTHq2bKyt4QG7kIBsl2HUuS1PQjXN8mjlZNfvTU3/KHRAl3Ig2m1vDuJl
EvxAh3svBrTTIsJ3zX/SpeLICoI3VAKlJWUf6yjTY4qbBu9AuSOO/8LlME6cHtGfbnzwjNuBF1oJ
L9IoEVb1TTxGMd8yu85DEtLrhCq1wMXdNvYfvXX+P8+7pfmOfMlWiAbtVbcHC0hSfTQVzlxq82da
uqonAcXSDBYfwcmRDZxAcskkqm1TmZu+9cBftV79EpwrNAblWqDSQZOVDd3wtwisBEOfXsx5DltT
ECEqt5kg3OvvLpx9IN01GpZKO1V6ZQ8IR9Hb2niZGCaRoqHzVx6kjI6n6JAvxwqoxaU8K5PvkGOv
BjEfZGc2WFKyv0lRUwRulmTUPRuLFZniP2xZqFGO8AmUziJo54RfArW+FIfUitD+u4F21CTdMuSf
8Yz2TXaIyslsnY7h2zUgLmK15WRtbAj3l4kOWGYr0tqYbFJK/oW3eVnJuBkgapCIOae/sx+uCf+9
77DsIgQDLiU2ymLA8gy0johg4md/OACnk2Nv36ZCFz8gZsGHWTas2zYdXAJGM6k8Ya20v6h5dKhT
R55jTVdnyn5bpf9CYviojicUT6oDSr9W8gKpUHsu4P+p0003QKbmAxuyKvSDWcciKi3Px2wsZOom
sAXXYAdgpnQk/eGPiP8LceIIh0/HRx6mIKhjNkx0VGcKxdqo8y1JGIV+2wTr+bMqwGzzFjBfh9NW
aWdJLrozd0ig4HXrDhFUZS/zeDIovbRg/e2MNCFd9PtJDvpS98rU5YcaC/Je07JwKqezXVRogWnr
kdSfLLia8dCkDJnI47sFv+5Dd6dt3p1xH6CaMUaIM91H3UHw07HnkZ5tpzpq39POPCLJduTaNOGr
mIS9asLdf34nKipx88yD7l7tW1kj+AndeTt+7YpKuMX1buP/do+KfbuzxCMFCY2QRm5apgUCmcwZ
+Bl2IJ2ICsWDUfd+strdI7MFkbi1sQdVm8VzJT6nLqyhEHP3KfB2Gp4kXitMSieOMt+mThB6Xj+Y
ni4HlxGvuxu8ImdoRrGNww1B/UXzcpO9fb0zoFU3xCJPg0vX75Nm1EQk3f5HAhJIwTTqipBhpyaZ
Hpa8130DVg7HpGRDtOYEn6STwU9BH3lLHueDqpkGuIevm0RK6yTAzgle6jm7abP5BOwbSPuXXo1P
wjomJe0xu0ZMohTmoXac1xjPyJJAV5lJA1nvJK6QyQ+cNjoKu1/v1PSIT5sb0cciA7XcoVe9gki9
SPeYC43/uVFZAn/VnEnsUZcPWwkmPvkpYJ90JkdIH9a73n94IAdRSoMfrla6sOL731UHwz7v5mJ7
nqZ0Ci8Yk3rO1KaJfgB5cRZjpg6Ef0Q0WvSnctcuio5tjnibGRg83DjMquu4xORvtCbbWKBYggTD
kzQsBziPdcwgwVyvs84wwQNopcQhCA3WPncQqUx8EvfctZ144jcm87sa2V+IsAxPpFfQM/3i+FtN
9lkldhO/3Fja5nlOzVsMU9Es8IpOys7Mh3syD5SYjqvHIdAalGtOLJcIJ/w9iWvRRNexcmBMLuxi
86cKWC4v5SmUIylcBX8C26NysiHxnnaOAD1QbX375p5uFKaw6bTGb3CK9xsPjuR0ZK/rt8IYBUIo
hmr4vvQLJKbaT1GxtWqKWIZhSiUsXbVIZRNHVkgntSpli6GH6euZaqbqyYZiGcpra690wPsYfwvJ
ZmBUAmy+1HVJ96t2vMr4OimsJQRtmy9i3t8Ll2xPiv7rDZzA4xsv/CiNv5IW62jtp/SRhIiQyJ0a
02gqJoItWADCi5SvRai94x3DOE3bZv7wwK1hmcUofqiEmIz8lD+q4/GkEOr5pcZc3Abixa8ku+SS
r75+5MHGjvoD2Zh8X0HJDYFw79rJvuA5MSjtkjKse+VqtdA98ZlAeiHIBhsIkA9m9EZr0cY/hYis
Ih1CyV5sO4brxN7ohq+FuWollcOdVRNKtNvaROTVwMNE4v8d4DyTzuNZUqhiiUDJDJwpWKWL0MjH
4Jz7awyGUQbVq9WSEn1BeC1cRaVGvU/kHwmgFIMbmAau6qXfLjIb2n0B5gcOA4dbeUR6SV+OPcCh
QhS8XxMBJBxYuTz8aWg346O5L/x3JFaE+uBCp8vMiCGCAn8OuKp9FhM6OMMq/8b8t7Pa2vVI0E1y
xdVN2LYr4iMm9sJvck6Ei24aTEOBVr2QAeYwwjS1v9Qp/XZ6eO/sYd1k14XayzjTnZNd+CrYTX15
Oe7x7T+iV+gdGVLW5ASMvOXBHO6OXrIYA0OlpuetwEX+k3V/u5N7C0ebrlv0HHOuG57EVZ8k0trM
E74VASxKM66w2u/N8wp8vDziR5oi3pLe0Q70oa8QhCyMb47Agdsl78haLeqZZ7638kYBo0Fi6jyp
e8f4fLY5/TVdiMDz/hs1ZmXWEFSyI7r3JlOYfwpz02g6byyNQ/jsERHeboNhjKiLIEniKvfmnj+t
ZIw0sp0AoLFtg7m4bG7rXFoLKmaZPKFWjIG+mS7kEGmMVFUhTZ9tsnXw8gj8whJQ4jNnGqe+ETd3
9Lqfjhzq57juS+uv9AegEQYtvMMKRs0QexN7QoZGeQ96Ln0HCxpC2OyCNF3lIaTrrf013o2RzHsB
WXRnCAmW5XmXp4ctJsnXK1MtnHsce2HzYwWCzQ4MU/zajf+AaohzAevGTe1UfYYAUQRjM5c90UIp
5VrlfqWtZSIR5Y18yi4L6p8eHsqo7/tmnGcY65oMU/bXotSPN5mQtmiBPy/tMUbSopXaJYhAcXKc
gcSaQcw4WVhjOg2fFtyyUdqaXwtvm9+C/wmutvd7EFOT0nKwLz5fANB0B1/54WIWgf1bIaFxXW4g
ZNgSLwAqHh0zz0Gnwks14g29eRZKXSkdcy4tie64LAx2lAVu10I/3dLFbw1PPaDyWwQ6SgxeDiNG
LYCLVDTJTHJ5qibgjiLKpJDA+9dUc4n0n5UHlddoT2Rndum5wqHIiUJSf+YhmmBdzzY7wBPKywj9
8rdJW3wALBrfSZp6zYdMKUeS15hboAsMVqGgyycVcVfwldYY7Z9dB+u26gIrItqMQF5XpGLLnvIO
NqHDf8svFlAegCCZ+Rz2CTC6GOt88FI6wA79oUlr+ZVrNENASSsQ6FOSOz4YiiPa303+N/EopYmD
2dxGYZoXEY8+yQlvXnlcHzofPbEoh51ZXdC+1qEFptVNS8e/RLgmS7Ojtw7378OXn96GLNrIiihP
KYRaQiRrRw5WqORtxiSolTC7nD8maWIsHff1Nq5oQTGPsA/OzSJn2YbijzB8tnwNKtxGpAZV0qms
aj6qNVQhFmwnTc2zUFW36pwlacZ99eTkiBGICqGA5FOmFVkFoYYqGcISoUB5SWAIgRwkyrrM42qU
6Lh4r8TtDSji99/jkCXT0xmK3AIV/tUWHKa8HIAzz4DIbXpf/xU+KhwrWUgHKz6XIHbIxucL+T3m
YHeYjkQOjVY0/qS4x0jF5qlLR5PjRMpWxmCLfDZnxcSAquD8fjvd9ZgQbiQlQaVlFHcB8N7vg7ig
SGQDm3iwPmDZqCf6ITXHOpzzWCkNcf5qSd7dVSzD0e/EcVUW4ioGKGHyVhKR2Wjmz6QSvxjxjFdg
qkcpVXytdv90uwE8pB8v8MGC88RlywNrfNiamSRsC95MmlCdRCw219/0Ol2CQ5LX862ZQpDOfloH
WnGWK33QzO6UvvKXy3atEKa/56y5V0NG5VG1F1zMGBGfERkOhl/S3jtiYyFf/YoidwV3rEqUmwBc
VT8cE2uF9Un2uR+dDqcd8bjDj7Trq3VzTMCDhcL7Krpd+LGC2PwesXmIJ+HARVQLqTUTiMHUHwXl
VIXdvZsUzc2sjkq9O2Z0eU0McdiokW2jn0BSwqny+qxGAm/zMzauIu0M7wJLasnjFFYmyCpjVcZx
GIsbAwak27afr5og4tDyFjLyRlAiptqj84NI14kx4sLlecHJ/CZmP0+um9vtrAIitrHZnNBEUjtH
0qONlE0arYUTRUKDDAmx943dkZhJRhqcppeXRVhdILa2QsnIfb1/vV9zhFHBzGM5miDgvxgxifAz
7+tiGeq9GGLJONVj+01cp+E0wKwnhLfAM4EU6QuTe7/cVx/CxVYDhwRVLwUQ69tbBCBmMnU8JCNO
mNKNznRyw3DE7Atn3AANffvVfGek7SJRR78PSwX49IP1L9wsPBjpTNqVQqIlBrS3j8tHSx7vn+Cv
mnRmirnWI0KZ0Bo+9NfoFK9Wy3dZ0Vc4ii6HupiDiZWMFZ9OK3ziYflcm7u0dmz5868MA9tJnMPH
f/vdQjRgnUIXs6BnOYHvZzxfelRVLkmEaTmZDk8wdewV9Z1iBrf6aqTf/g0koinnLrVjyErW91mX
SjQC39tDsbUWH9P96T7jH36e60jnmlJcg//tcnDdclZMp5xGpx6kJUr3CvXqwYurIS6bw3TE18mL
BUkws8TY9K8z0i9/6UqxuGGoiRYk/WINauDHI8ZEpHR/OBvzoSMnEZzO197uTIqLP4a7zxtPnyhT
0Td4hvshWPUS7V2YFLy02mOQAHKo+jUrXpzbupkMysQy93ZtmJxrTQo6H95+/rgzoEMC8VUt6SGG
pbVMYhuamiNfbdmJLiaRq8Ms0tH5UV/9SKvFpzDz2+DQS83whOUznU4flznX6JkWxVIBQKnlDRla
FfgDCrprIdQjudW3SDo0MiomJOtgNoO9an+gsJbllofT2GJEFJ+bo4kaP83vmWnLJvCm9e6NTmYd
WPmUWgZ6Z89TrIIrsihxlZ1qeD9fmxa0oaTfZmE30TfiNFHgMLxct2nFnyLWCzcxIsRb5m6im5Dn
0DJpq6Ast3Apn5EpKyC7ppWME4cUfzC7dU2vInj5l3NbM9SxOrwW6WeG/8DTCpXKhyE1NIcQNF1T
k+nbDU4fKZeTj3Y95F6rA8KDgauRxCvbtPaX5MMO01sJv//lKR8brBxVxbjdh+1c1spz+kJJ3ys3
C4ArkUYZtuGkRkHOeNPpPW+cXfVGpWacxaLzrr0Th9IqcVcyxQsB+17uqyaXCuzn1aNG3JHMFWh4
Fd/dT+8HRT/jvkr/JUX/iPD3n+YmJdo8gmZkr2K9ZcFTjQLQfRDRAHmhFWu8Mtf5lB8wz/W1OOKR
us0PLAX61eMRqhV7GSf3Sw+GmhR56WAxJAZnhvLDqTtG+oZcEibxVO5eKTlD+2l9XDlW8kP78F+K
bePtgHKBaQFdbPfcLjRxBUmzOBUSGR5V2BWlJjGx35SGMDmw6LwLG+qJAhFTQsrbA4HCGoe7GxiV
+wL582XIqw0nqA5yOry2LSrqhZGOWGgu3LqNUpqXz4yNq8G+Ws3WyIxhtA40sJi4IG/yQ1WDOgrp
oTUvVhkEv5gosGYo3dVDWUU6OnnhMNUP3WUf6EEBeyaiOosb34EvKlr27B9KW7cvd1zViYT+ZafP
+JF7tdkH8k/CeNZhmKTkLlgWWr2mpPaVeAYResXr0HUk9bTw+M9l/Mona3TaBcwTixn08WmaKT32
WFtIWpGM2T0ccbdjs1qtbrWQUdxXAndexU/f51NSUNuc9wplKnEvUCJ51vDDeclWMEpr8G4GnHwq
KHLXR3truqClHi+nL1AZmBWfGoLz2AkLLSZTXhItrAPmW/TF1/Zsw5raaY3/RSWEJ9bmSp2M6utk
TrieFFfXtCV2VANWdr1Wk338IqMyDxZP6gynd6M0pHb5lYxyy1XU2yuKa2KsLxGM1lcOec7beEYP
CaTwLJ69N72FHKG58vFMu58m5qOBfG6MXfciKuuYIluylxv5PV1iLMzNJVNh/x4QeEJ1ealeaaLC
Upw2mXg2CEuB/kC/Jr2WXmn6gG3kFFvQh3UYbLr6+eMhL9nBEdcJ90T71yx33g1m6S6LXFruoNDo
qOlMI9R69zG/cWfC1BfvkCX5r4udlhXy3r0MTh7b1UuB0I+0TofUGinPpcyQhycmhjnTJn1eS7c0
0RZtR0CvCEf/bMnRYUx6YWFgish96bhVKs6EtZMpWaf30m4OVzB6tzfoT79wJ92pFc7IyJedeJ3A
+rnvDxgkUaTfSzOMTJ6neoQyVfHFOblyjV9zhVVww6dFFqJ9iWScSDcxAynlHJGVEoGO2ep6bvIa
zevXJzzJrhuV/9Gi0x5bF9xEfAsk4Kt0/8weXmHf+38/kvauBUnnpB7cJj7K6fPjwnO73lpQ7REn
4UokUfIyiTpVFlAWfYwQE6Ie55v1xm939Pu7h3rUUaFnex1R9KIiLizA1x7KFHhAmfEE1jNgcAIf
FL5PHOem/L7Um3ZKPmww3YRKKKEkByXrP3MololfG/it5INj+PRkHceuc+TIwvVYlb4WQNotkbDB
dBsMQfjECLq3QmZQkHe8cghC9D64anc4SccT2XR5K4o05tDXokpbIrU8syS/mRg/M/uTpPLL7Xs+
cPvhoXilH55YpN2mIE+IXLuvMjouuMtY9SSK4F4KNqa8+3IsbAs410n+F1AwLtjg33F2MIHuKAq5
TAQcHVmMn6Ok679shYZuq6u8/66Ejon8LNYVLxdxk5WbGyZTIjosqxhxWlw+OaHMej8jsDhk2wIc
cz+JedFWaNFGkRfKQOFdCREz6B1Qt5/kQDSa+LT4zfk6FeF4NEMFzNKa6aZEdsH4Km81WMY25hMw
2stJOiaFe4mlC9SfDb31cPIRmYSbD0dVPrvZ/TZHWb3N78671qq/wQMysJlEE/QveKYwdT1F8ErY
RTQyx2YO3E6GWHaWB9pHO4ZuyOEEr7gEvsIe1eDZuIA/ULAhEyZrn0nyC3NcV/upX6fS/XKHCqqo
OJsiUviOgVE6b9O7WkGc5NRZtCDrBvkIXl2Ct62H/xbqe18F/FRsISz73e1guH61Q93yrMxDMx2O
hCVsHZcyEMts0hmuLYHocupSpQEflFMfFqxjy9cPrS0O2sULyDgLBdOMoevnAT6rTHfD/OXmWBg8
QbtFdz7hKq7BLdhOmpasmyIOEgywFLKf0MQf6qn5eriQWfpKwfUmpiLQC29cPeecwMRopki2/sO1
VTnkDnypIMwS+Hd/aR1q+t/gfYfCMEJKxX1lqaXXVA1YC1yLCcrQ1n3ENX+jwIaixFajx0H5FuGX
BcbmFrnQe4OoVALeVukvloqNdZ9XtN9hsKUKtZvBLaWGrih+0aamOgkisUmJaTdIFsRTdqRphr8N
Hpz+vCsh8C4zf2gTZcA86Y2UeyvuJFYeBrwx2mvOVJMFgXM2GzlBtnI9fA2SxM5tcXAQXBHZKbKY
QrcoAHRmqihdjZcxTeZgthCRRRyZV9hJma16TRgCTcSdQqVyiXsjWVQFIwWvjks3AIUW2TKkJVOi
ei2ffbCN/kUQ7M7iMd3ZHnedhR7eS6GG5GJUfwQkbC7WyIHbqAu6NIyE2P1CLkqUfO0eKTE7iONv
MFCUBGvnJFJokWKQGB8kwnjt80iLQQ5SCMNCt5XSfTmFZbtNAA8atgTrRn8m3OTwP5CdY8Vugi6F
XTiJ+pOPgZLY2xB/57LTC5BhgHRcCsf7SBFd9cmnlYaC9+avCL2Swyz3DZpTRD0mFlQTrfUihTQF
/Y2OL7iBJsGkqYVc/bJ+pgwhOhLHCNUOdYSYLADq7G25+oBDfBSNbnYCAxasbAG+eUXeCEVsnoTz
MWBihc6/NjHF2k6QvqCcnuekDt46v7HHhQVRpbs3aiCJsVvU1ccy4IWVWYU4GEwSlg9zsW2YGupj
IuVnLdhaWUeaNkK+VYlOkjrtT+szd7rK0+ouX9pYY+SODXMJusYCcvf0/vQq+eNF6yC71E1G8b1d
ymavN1/UJ9jSJjFJ1+R6SfDT1BUiaC4G3nydP+T4InhV59ztyp0ywobZI+TQc57xUUaixo3YSzvK
rUCHM8K2UhyGfubMwgsfh/41IyMmD7ZNsZcCGsAN9i+6t5Swx3mgGQfxYcyKzk5NPvJX84rI/+Sn
nuv4Q+PyBdNzrPpW0g/Lq1gkP7MIskkm482YDvgbL7jFBNwQuQcVUZgxhs61tO26DavNUB153bhP
NiQAeTSpbjsWtnNkdWTQ3l1EfMTgpJkek4ikAcfJC7IsjmW0H+ExPKX86tyWvszdsMjeoXAlHoag
NLGdq3G7uCxuvBrUfcQRuRQRSZl73HXUSHMQD4AVIyKfRtSfiIfLliOLNq+ncn9BAe4kZb5/SCWp
V0+m5f7CC4AYpkPlIVFGWTEHHJitp/COpkOs+vCGq+e4krIhZwSdU6+H9KEv7VBCUTCF2L4tI7GB
O/kWXOqFXBI/M10BGGQYRqHnh+alCNMFKwF47r4SeELbaJsw2S1tVTy8IgrNFd7/tgY4aqPmuUkY
G5PFL4VtvpuR06FeMfPLTtM+xyo8Uw+0LVrYixkN9+RQQ3hBFwkTAnMkRClZAUxawATlu0hdHnM1
ru4ivfgfLABM578bP/mAd60nnWjW1iSNwSpxKQ+hgObWLx1i4lDq7pJaLY0IE3CpbywtzVhuxe5I
pP9PZpf1fwDO5n/nF8Pg0iql0bj2f3QE7OFWvZ4IUXQdCdR24z4HSnaubeGISWeayKUG7wVLrLYo
Pumi8sVQ2xG5q2jZSCM+NaLM42K2IgthH3S1TftK+zp1RkQ/M2XAG3i3SEAou43aM90b19Suhd1O
nXLqjmm63V4daMA3bBTkzvq1960u3DwIMDMYhwZxFxMJc+ceNBqwgI7GZDENM2s0GMnzW0oRPZ5j
McehJH0tjwNoPWLn2NRTI01eejFDD2YzjimdlbgSkfJ6R/N7WGUKVl9T2hSRJm+q8NpS9RjaAtLE
yZHA47KQr0WBBeHGbiBKWnye9eqOrMvUqrK1GVGaLsgaV+6TkNyrZxZzJY7BHtaa192IDX70z/26
H5h9DjFoofFeqeAnfk8jlzv6utmb7QFi24dCCebH2K6otB3TzQFHPMVrBV19UGiL11eimznWHRwZ
SiDfgzDj8XjPJnkOaS4KDajPCT2EnGvDIeB4GgzhaXPX6n509ja9mvqmU34uWOoHzLSsCEcpt8aB
muGAxS4Afvc0gsiHtrfmHPuMyF0MdmIDpR09WHXHt2d0f5DzJDf9Yeuxuid/syrlX+YOrk7Q5FxA
GVh0b5MK2/LCfjfpEC3/C2klRDHoTnfmeOT/WXJn8S7/AWeFdSICMtfjyv7r7U52tk2xAKm4t3k/
jvsObd2E8REepN+vhwQXQLhh0YSCsKSbMATMbADB2WZvr+tkytSaRntKGGcWzktCsyv/HXhJvqOG
Zd54hS8c/WhmixuwPAcgBH3CIsJemoDZL34e27116+P2QJ1quFquwu7V3yDCkwGV3GG9cZBiNqia
fAx0ONAMgDxVi9hevWvh2q5kSsLH2lnc+tCcPOrMrkqOxROMGABEUMprWFS6dbFKOygQdoBOZ9Il
65Vb9IIhKBzg7ROQ6fxy6TyEfIA4bj1Yiq8FCpQY1Uxc4hZGiAkmRzDywZDz4c2rNJxYo2m57QRt
osgWd7h44cTeXPstEzIyXvxw4UW/AcU5RUaPMxC2hPgEFl7yQvX7H30p5WdTZ6Z3an1x3DciS60f
gzICeUieussA4xJhfzLm7getWbh4bWoQYZDSyh+5dDcEfMdEtjyGeXHuFPXnx3DWevd+Yld2+hg3
mjEUp3vSnVXZyeLBvZro5ZCctgWtyDHkqiwe28aOafYQv55/sp+DVUZ1omSH2g5MREQT7ly+RKGv
suPiexl2DHNTGaSqaZGggj8d4ML5DG27Xf62yRP1WkrDwX+zefgrxEHdzXo/iuxVNZ1U1roIDkGi
PihudAS3YnyMa4VDItcgxGWDYaQXlO+X5MLsRa4B503EqJOB30J7/1EY+7+6kYqQdc/SsVFVuPcS
zR1s9k1eSOe7YQjLgyazp548+G/XKA+FajAcGaZdOfm2cTt3H+2MivKoe8bvKveEBSudEHqi+cjf
H3OOi3LFHY/AacKxNPedEZAlnIuhNZ31M/VXq24lVdndmJkroplBKDxgb0WILUpnfSnnwTApiutH
22hdYvVCKxuJxy2NNj7VXresy6z+jE0KUZqGWNAhOIQyKasL5S3qn+vm6+i7k+QdZUQYZCp9LLUM
X6lQvwrLkT+Sh1AF4H470aEplfIZCcai2zwSl2vliM7a3F5CYZaXg5mnEpdtOpsFyQFXbXb1mFDq
qfO2hxv7mrUnK2Zlpw1srUPXv6vnR894IwB1ow+n4TWMBMe967Io4BCvptUeXXntFWRThHAMxTRh
MFIwmRgPsBuegsAPYy9gOKs0S1Tl6p+a7lT6Aqqas+e99tyHtskr4SGgGEe45RY1G3aKFmxhJ+K0
3bvO3D0AG5wGaWuJ3RoNDUUSX9rpBEU0/zLKEgn87bIqGQDKGtpgIDzWviVrGXs6PJI4kdi2G4+R
tus/gQqW4JT+MuzYt+uAiiJwQ9JCgrEO1f/lGp6uug2aW1ANDGFiJCEMASFyk+ZE4gcKAZPQbL6f
d3qhkRPqj+aqUq+xV6eBVO52G/No/Qzi6GwGrIn7EqzHALHkoywiv90QSZ+8165BzPKOnUYJFFZn
m64YdeXGSIxAVwJdjKG/GaaymSPIAyceOqdoiLR40iS0mu9INSz5GguWxa+w1uZX1ItA8FhPkfJn
O4vPG7Xi/iaqaTEiaHi/WfUD06dJEZR3ou2UyqoLkBAzYX8bQfRc1s28TV2Uea2Rru25Ffp6HL1G
jqd14w0B5cWS3Cznq/D8IOeLw7EYRw8C0YUWWlVQl53ztirBRIdzObf4cC2kVmn+Xi+IFkZ3JawY
hsOtjD0KrfeIP6lQl2zcYbNNf6wVBZnbQ28/t+XL9FKC/CNs41qXbddW1JNFRR8FTYfiSsPBcHQZ
CxeoBMwxscbr6AghQyypiqDEonnYO7Vap41mwBH2KdWtUCs4bQO53Bte5HECmBF9sK/bfQUxxxAT
v5hryMU6Y3UBXLII6L93aL6KHDUyE7wwD25CDbPT8YLsTiNjS/Y06x7kEhxnPVea7CSG3fweEVkq
CNMok4PSnwxfiAGtULOWnMhP556Al/9UpFxFykb4hSlfUpnOPHcH00ZBEUFX2e3TE8Cyufi9Xdr4
z8Hp7PxKGLWQ7BM4GUXicKMqgoGFuDAXdHEsBZ5xzqmO4knl2/BvrK8NwKSrpbIzP+W13Df4L3ro
5bsVR4Q7tuKWsVoSQsaQYEEUGmDUss+x1MdjOuUSbaW4vEJVFKwH9OA5SjLdqgbJM+MkRPCB50fN
DSTUMNuZH4207/kIkmIOymXEoJj4TlRi3xDgcU+2CZUAql5+kM6j/tjSxjvRVA5xFIwEuhhU3m5I
zhMZDlpkQ6sz+2+wn8fuOw5VKlNAvfUkzaZ2RJKAO30uAtX8jRq6GOq9FeFanWPevuDC/VSCrvrK
SNx4ybZwWuhwq5sPFarnzJ0sVKC3YHzyb7Y/on9ZKNAQwijJkNeiMbPWVwIvVKZQtPyXkS3Q4B1M
wCPw+9/va7iBKjitdhJOKv9oxZJ5biu6uIwYfzpF6FYqJB2DwBsUhDFlVbLvoYSLNGjoZXTShrr9
dTWPhfeONIKu8r1ZcLS9jpjjx17Iaxp1K+ukH74vaPjRJ/LVbsHUSg3FMRGzZE2q3mxkjamtt+8R
4Y8Coo36arJBWzhVfhrfj7lIGo+9oZL8DNYIiZU15EjKXyy1FX7kqrO/KN1mIuetgdZpOXHQ6PiP
4EwsddoLMUlV8SRbiM73e+ns/Tp9eM+19TUTtDTy6rWD3c6qUg034z0b8/fnI1UWdrCGG5XMvW4t
RYda4IJHyHOR9q5Q5/zoTS0gAfhH2b0pcreZfapP5qCFQkwTVQWdV6KxAfOi7ySKkJzmFdXvS0Lm
/rLgkKmU+850KitWtEJ4VKY4devKmdWcNn6VYlQuBi7O9KhZSVYzA0z3wkvaJ91hcEyu9uGWej4P
T426/egwakaKUrKOthMELDISk036t9rIfotqlHrizbPq3RfMCOJjxBFIbHoJPK6EJ8eWiQMrL1Rm
Wk7hZ6F5Mb9be9BpS/e+AyCu7Sbm3NY8gZDYIKVIMmH7gSLmcJSQY4/Q9OOjxQ1x6GSTZzWuN3K0
V9i6fKZmndhxo42zhjF8sntuZQK0WaNw3PrrTF2LapB2303kcOKl6m3ph3UI4ALb7Q8GfUhD6xdp
O80bygXBpiQv2bUZ08QiZhZRCXtpxkcUSQpIEs86U+OIV6J+xL9QKbv//JrzS9xBxOa8PNPfC/+b
L7Jt2timoQ4SeGgI/YH3DryQIQmAy1dIiEQ9vWAoRccHUC71Yw9DjR7DxjJGgFJcjxWoPyxhtwVT
kXYLDYJ+KJ60Ubm5MwDWAONJFsw9na0ImHmfNY2ukqU+p/M52IIkREaytJq4gGE19XsbBpBhTHeL
TvPo66NaO2jzAy2HZDu2GW/f+IFBRjgrJ7SWSQ4vm7SlT4DsTkaIdWvcNjetMvj3uw0x12xCJUe3
f6x3QS3PhqRsoxLgpWRY2Qdawdk6VdYWK0ifJszAgk3dAgC3Bb7EcQAUQTZGio4rNsWEKBeiE0Gy
2mQYB0GfGx/kdagaeWgwVpvM7244i5JM8pYIRm4vIVZ2ORHcUgGKz2S3VeYQa66mPpBR+paj2AB8
kfdd2Ewob+/zfC0yG0zpfs1KAlaGmdaQAc3N71ZBxvTrgo3QDlCIrBsee6KaKiAwWMGWDuD+gTVU
G383q2Lih4XLG0qZ+jFVD6nWVCmSDVFTvv5NtWwqdfJ1qDz6XBR5WZ5SgJBZ1/cLj92m1E+5FMKQ
dUivBVBWv+u3RFgZkk9xGtdilKu4i7gIMbVF2Xmg8jo2HHEEN+0e1P13AcbX3DUQB/Q8Ejo/pnTv
xRDQXTJH1A1X67U8FhWKGCkeD/b0GAN7rNHeSmtoeNpWKyKOFJjr7v+qsPOz0OKYRfAYAflWM//K
Ucg3t6B2/rVeYjb06rSE0GbilHGhco2hlu9jOYT37w6AW9zFUdZYdT80F5+xnznyBpF3lTzvDxRd
em+pqZW4Jeqfl+U7ZVcgmK9CzN7EB5ScxjrGNyyXv3RGDFAnV5f5TknbR9MI2AA/hm+dy1F18Ird
7aUQHR/f64Ksp3md+9tnD6V16uVMSTil1ECya8ycRIAnSpYGIb4xScwJeaSWVTP08+of99IoHRmr
h1Dpmb4T1G0fT1ciI0ib2CUdpzgejU5M2DlQAylTxxm7XJ/xebcSYPY5OcCtV/E5VTLH1bgkBBcG
YQvT2mdEm+zn9BibX90I8ugFHTFUIEGMyf+GHwQNoOFGjIJk22F8wVF5VYBFTx1Do1EhDR8laMJt
a4D+z+JJmYewvHWIiJ/pQGZmc5+riYwBN3JRzzv5wiCSpsK8Td1OD+2SNRb+vEtKpKTkDGZAj+Bj
jyU9ZrKk7GMCWZN5Vgiph3zhwYuoXYFC2yuvGjw1bX7JRUCo44jlSWxKW98XKtdlialWJfhtER0l
ftgZwxkzJx4lfJMMFWsShO26zBu5L+OGCDO+NjlA70fA5uB+LRv2P1Zx1KCwv1OJ9d1qnRqWCYOJ
ySBaL/WKCPhDPKTvTHR1GaSTbmFC7uMYLZYq/jArz77KcOVxIPICVN1oix2bDKQi8HprR/O/dLcg
DbPKg/heV8yuTAQsLkx0VskIeizvpo6FvsUT0UYqdVQT0MV8IbIUW0Z2Y7D/GrNS9G7gCm6kSdiR
zKbOeb2/aTXVqwdroHzJ1Z9yFqgU7wWX0/WVODR87OwbQVMJ6k2krH+cyHQv449mykdm/931jXfn
SUA6UEBnI+YOOIsuan0c2oaRwHop7F9PiMfjVLAo1X3EllXytf7hBE9dDfw5OT/lPH2pSJL1mjw7
xRrM6E/8aK6/utGfoJxFIM77KM7jtWjyfStvoa/51/XAG0UHQFfmR4EKS5aZL8wS4WWXJA+CoNQu
VylTYeag2yafn2X3ExrXJrI/NdPVLP9FJiAZvPgkpwxyCsyzOmkjJ00xfp3BTDcOc/cxnoXLZNpH
mwTDxH1G0LCHkKzlH0UxB/gtYI7Tt0h05mJtYlk3ydEuOTXwguUEpX/n8rKd/ChjNiJDAoU+arhX
8eCtjekqOUXYqWWe9di8t589b1VEY5idbvpH2qOwVD8J9ZVvwFR69jFUOhNs6wTbtB9Qejcjdxix
KBu5K/40/D4cD1ruOvYhPFEB/3YB3T6MCDVBsYne9RB2TY57xun876/hQ400VRWqlPiREd/JWs/r
8M/pNSyrFhXFyN75hnnk3RYqWkvHvLm/16iCzF04+Xy1P0U+bu0JKRRkmDtlCaIQ4V4YE8EPuKOt
LJNBALk8aCqMqZQnYOJ5Tm/w3SgToVGQchdIUvoxo2U2rI+WsQSQzQnKHpODdcwpapeff4bEtC3x
+L6lu6vtbuu+AgaiG6dX/s/vCs3J78Ow8AKDR4jyJxJHEfcukZZaMeHH66JrQwq3lI276LBGOe0Z
UJw4Vkq/J0nFyE2nuW1WmspXmyUlqz/vlz2TlYBMCXE5/QFLd+9p2v2Cm0bWGvoCFchBoF2FGJRh
IDnuR1DeW+TeXflDoLGlh4dpo7VVBXLPTpkvNqfCTU1plxQFr4XFH8bT0Di6docJC+Bnfz5j+WQ0
Ihs/aW3p3wclRyWLWs0FH2UQ/9YdmOymxof9MpoNlytXRL7uCtsfApw7b5vDaBp9sh9DY3ONihTo
n6eG0WeDq6umaB07T/zf0jgBGxfVZ8UzgdhFENeeG3BnP7b3tQ/5M/+mA1w4bz15nFsS3usHFRJ9
0JXf/E3HWpyXGOiJwBNeRwa3S4c0TznT1rqYPY0RAFnLDoHa46d3DBWxgxkRo4BhFEBPEAVG5XQD
RkI7r5vN92Eru7b4h4Ir7uclrRTZcEJGFYs+1n1gu/nHhom3CkWWTNM3l9GB+KpRy6gClkvFsnDz
JFyCZLjvMHdw0AqaoSLeRekn4v4onpsmTz3csCMKzKd7qZQNbG8yYC7RCueM9BMVGIWSLFDs+WhL
+4ptmTa3c4GnzuysD/8ERqmjtofZJMRm+ff7wHDJk3/uMgyJ2IuF+VUgJSYdttFwYM3EyR89AQke
YIzIBWfus2RqF7GL98qSB9gxlIQ31xp7i7l7n2mxrgRVv8m/YDtnTDFQxLnpsP0fQgpNM9TXGJiL
pFBVie0QUU3VanceBwVKbixYBN8KanMh4IlXjHTtmo5wVzonrqcjs10jzctuRSaC36ehkM6yTH6y
tiEtgH/j3RNqs7Yk9XJTn9VNXIy8PyDFJJLTqIrYGMhv9e1SbHJcXEssDNJqm8WSusiP/ueMjltk
DhNO3vZHDvElco3NoBI+D85m5b8JzzYPhQTUwHOKD1gWK/qVv0D+bMDjuBFZV469/tTbKTrBvpnb
W65M0bThN7VIvIQiq/4UzqXfSySuGQEWIGWZa6XyNjUl1apbROFu09bQ5lp/pInNA1WtGApU5k0u
/xbvBhYTPTqZiAwfQOOxS1P6H9US5r9vxQXw6sBqTTsEyz9DEwWWq1ZiDlJWBzS6I3RICavxX3tS
fIMIizN/QbtuWVj6k1cwCb4bwb9uF8WM0jUiQPOFyCmBEUMseF0gfU0MtdzLer23/q0AGnHd7O3T
1kRusj7wakeC0k2s184IpDKX3Li6A2XqFc5sd1ULUHjJ48dODsiM7xHcMWa9R/YtdhRYYK0NDUMJ
as2+1OzAi4UpFpdZrI7ctK72VEyvJBrjS6B2Vr+N+uvEXPeYEXBp7euVmms8tR8br3/Te6QQyZvz
QQqGvblkAANICuK/yBX0x8iIFhassqSl8Ghnv/m7lFJdrhlIn9nP2zQBgE4wtBSRV+JBYEcVpA6L
kvGPbn3jyaXbznyzLkpZPQAMorSz5roUna6KHDOdJ8fgJgByizSUW52lxGXil5vkKc83PQ24R5wP
PIxURt7Zm2K8sLwxnhSea7ZOyenWgZc4ra0XfFrQSalrXLImTi8rKkMpGRxB/Zk7Jh7xrZjdi6FM
nI1elTlejrzzVLJQSab+A0DU7GUvWovMHYLSMoyw4435EHzzdm21tRBHq2We0qbNl7tbc2SpYf98
A2VvY4Sjrzb4zbkN3F5SdsQAxfiFH9EDqFGc2jPNQWSmXlDQs652Qx+T2K71nNbAv4PAIzkmZ6RS
61nlds78Q6xyJMQY8P5Rs3JGmbsHKZVGYRIXH27k6i02Kc/OPmM4g+PA2tNQiO33amqeASx0AscF
/QBbPNUBF5j41PfB4T0w5ezdR4XA/AaCe/wFGIBDeZqCKcWBxqUEtf3bfydqsFVctw1gcf/CxFTu
P5ZTAS/gfyy6vVAVd0LQL3N4ZWChCNOvEmf2hkGIkul0y06UNUkCGGktM5yzOCEyFzeqpCRchU3d
JBZppyJGJcjxbSncvAP0Ch3NMXEvOldeAElkVlRl5LPB/v20ozix2rDnXVpOlNuzkn0ikUSQfUSq
p6RkGtfUhZt2Hco5l8rhX1pZiSpw78AXZxsX4B85WvUQjkoq23wRh9XZ1A9vuPzl597fVjPoow4+
h6HVrtaX88lSyphbFTMCgjDv7omlqb9h/85q/l2fBVKUVZQl/KGmxymqWfWCXzqKKd8JL8cJ0+YK
fhMOoLs/eb9JkL0o4nVuJuiH2qc5fcil58UGbvvKz11R9BkbXAT3nJul6t7ie1vJcN96eT5sQTBC
xNal/xePS5FTRVzBEt38usbCK7O0FbLGP18+8b+7AvdXsEkUcQ3djfbWSheQPcEcYrWgFHZych7I
73nAEYjYzbcPiQvRhSx1nhs6DH5lCJkXi7b7CAWP52vSR1tIcwxzRofM7H9OUdYIDDwFT3DMvU6p
aXxtOhoa/EDzuXziKWKtLw31s8Rs/W91+kbMv+Gq1sna6xLMsCkR6iqsvddiqkc9QlVv4D0gH10A
dNHlNpLbPmSHM7/jF55l7gUw+AEpddasRDONgaX27hZM6k4pe9fV0A5iSCb6SYt0izL7zGYjbdN7
YZp1uJ8iCAQojqQjkpXxT2By9mnEOnhJ9xniP6YNPjSCzsVzAahbAbEgNJTJBSFabn4uT/Pr1gQo
Sv1d1iLI87/lYaxf7mNO9ufXZ+/wLy5WqoI6YclgpQPGYG0FrgTBStLMzAAvEtuKjAnFSMYjf93x
dz5daeUGTlL9T1+Tu641mjAgPwpkfMenTQm94VOcVeB2owshkSfh2HB7PyIEO72ADGHR7dJ6ZSzT
5IJRl2+IRFUjHZXQC2LU+JHF/BGVY9+Sh4MjRd98vSXt02Zgh+7GHxPqHpo6MfxoTC0s3mCV+kFr
8GYGaoR7+UphZlbZOb1ad/+U9iY37jkmJkPjee+fgK5OAeFJuBbFrTNiW6W5mOx9LzPfH5vtGpQP
YBZL8k54rIUAUn8aEw5WdVkIxA9vRs37AUb5DKWbCsUBTlcpOnACsDHCWLQ42ZH1gslt1zotiS3E
JQjSMM7FF7yO4WiNGCmRNPauoeIVED8b716LLuX3lNOvajcjSRLrIwVLdPBu3VZR1FXtuCrBSg+E
dAB+8DlnBfb0ZKZPY/U89S4Nr80GECvcdErBoEHIvRiC52jbkOmvwn0BEGwg17q5D1SQbdZE0E50
gX1Iby6OKjksVMDPSOHz6WQhgfK4kSkoFxqs5LPYXYwxb46sMorpaEQM0uWClC4YDnEJYc8UmGS7
gok5a+iSWIfn8budObglnQ4zt5WASfqlz9PcrrDP1fByw80H9C2MJrhe9wo0IKwoe+5Vcc45XLtN
wlvpuGeeRCI6zQWxZ4aSZAPTkJavTaeK5JbFCinQsRoLZKVz+1r6qyEB3fR0JL7N6jR9jW4TpW1t
2QJ6hE0C4GT7uYWGXgYzUtubJpebxWbFrUCyN3k9H3UkyxO9tsqj5EG4+suX25f/mFWg1U6Il5Af
muZ19RdGBBPhF/EgdWadVcJhSuhwxapDasm3gesdLaq8445mzbkZrgAHk+iECdYfiS9fhxGVC6Br
PISKX6osiufr6tKdZ//05ZV8tOrnPyIn+svw4pL9yxuiLYLeGE3NAVZGKwifMYrCetRB+QCATJ89
3MGFWh2xSTxXVMLkrgocBpfcZWkhIpyN6Tqgwo+1t5PX3tYn88RWOrq6YOrGDBaoUDTXBylJFEeV
TWceHpEbey9v7Yz8dOks3jw/uo4EwigaRmYFnLQ6Uv7yh1Za7+GyB8lfnQYHmPb5UH3XjfFOq2nH
QjnHQnAFISfSGva6ye7s9bPSw357xWv52KnEMXnyPoRayKZ0nTJ7h5Pzc0KWHIEWdj8wLPxeMbq3
sMpPp72cNfrFFk6ND2UU4AnCkY6YjRSq0pkLcXPtu52STp263X3SU4DccYav6/v0syCuuWZyEP5s
O/dXtq/j7d8JXGn1ITaFwhWOC4booHM0OapQClg1VyfbqnHqXPapLg0UQRIv4iwuk8D0y0R5UjJk
FQyw3o+oiLXnso2BKq0GOEAZZv6yYWNJKcILpnxqLR3x+38keW8vtAbRXr+FVL/Q64wUVPN7mBQ7
UgBpY4rvUJNDgHuMc7SUcael0CoqCOifoQucnpqdQU6qun8tiVGqqr5HZdkPqTn1IIWzylMEM/Tq
qrj+rFOlRtT8NhnmKH7UFi53vq83z9owBWJht5SML4cusy5VlRpZpJi+1GLmqH9jGe1yK43TG3ma
tyW6g1hwba9qIfGlD57r6C8RNf4o7yn/aq9K9nq/6DqZuv+7JD93ATQTnRp0tJFmD5jlSeN37M79
MTLABTSAP2uP2ODxUo40nvxNqX9kpnITZcQRiQom7BdSNYYykTt57/tQaw/cy5e9KT2RQt9ODIZx
Dg1C4koYQp1rh3SREOXv85EqWBYtxqxtDnO9gXlf84WR4M/73H7WVeyy2zjp5ju/gWjy2ByMrPgV
hs89/kE0Sg9aKfpQmSCxUdC8cCq1d8RgE3ak60zwLjUk8RzpaottRfA3xBPqld2hlkFZZL5SYqyn
b1519xUuR27crFW30TMscw03ubKJhcG48atxQ8ZBQyaZCf7rVqP6yjB5qPGDi9cvr88vOgG+eDcO
Fa9ZiaGMF6NKwwwpZvTWeoN9rmG2JCKRqhYPDnUNyHr0LauzCKbTttHlyt9sCSidw3zqe/xbMTCH
ruHqR2gUpqpimpJbQ2hX7e+x/+i408dISO60Gf5z/BvfhqvyHNGd7bx+DCDbSELDi0g4gHXYmAvW
jsCnNFeYtTn5r4cEZ9A08IcJiJ3cgQzWQo6PioCafblLv58PYz8ASgJ/LW8FevdLY6twIr/0YO9e
CcmoDkbOQVDDw6Ah9AozcbwmPfWKxZqXDmflTdm8dK1oH9w3dl+hb6fnC5GHRYv4KKq9Ic/uQ8zg
8iC18WBjNwzQzJsONOUo9UW35QCs0U4nr/T+mhWemrRk3knPK1yQFReeUcKrUfGVWBUxnA15bNyL
oaPnMbwu6oQpe/gg5NlDfdZLiu2t5QTOakvegymqM+RoYjf5r+us5J9W2pOftve27I1KNCahbNZ1
RHNiI7vk7TcdlMwypR85NIG1LgeE7if3ZMOP8QmZG/Bl1mQBDydyKCZKBDp0XOf7mgcP7msmvqz3
+6MPE2mKwEFCcvH+ebP7a+vlrELiSq3cfZCTYZgShzNHyyvfe34Ty7pmFC0nM7TPYxwN6EbLnEja
11GE3/Ig7OL/rVJATcO4jy7NDZ7m+zbWDNV1c//qzAjOG64m7klJEIVaqAhi/31FN69kSayJe8vH
0CTFNiY3p0zVfoGRapYR8l2s0zcAXqeSApn/q3oYt4qcN0EmtXgKqLtZ2ApGM8J1HXMIlpF4Y1ez
v3iK+FrX8Kh3O7xCvwnysg/L+31BJwtvVJUL2hQIPbNSNitdz5QbscDMoo2vq0TDoUBTEXCu6f3k
qiCe+Kv7a+1utA4gpk1lFg3MGEUBdIMY34leCrzOmuQzVeKeO5B+FqgSkTBKntrN77xBT373DpPI
jKrVqB1+1qSynUwWA8+AFvScF/5CNlHxp/0jb+r7ndgQB9EGxvPIItLWdGzlR/LpaRlJgZ3XYRjR
2Qom6tz1DktjiBSvBokuDDKAxcCPyP6uBZlItKREz2IVDXZZ/jbqwa5t83cMQ3UEFkrbJYGAGHFB
XBdeMe+6MFhRrR/1nvRABpeIa4jU2cINVivggdIxRObQsJRrkcy4o8Ftnluaar3kh9RMHyMpfPsu
kAb17Zj5cRQnzwTqqW29BVmZZsB1QE4jBQEkmCVykJpGIlfaTFaDTyl+zMUCjktvVOGlIxXlYKpK
0sy9vzsVAlHgwl3VEBEw1fmAYHuLg32LoOXTs8hE9pIMg5tBYszYaidpC/+sChamnJ35Ohg6P5sY
3+dNYrJrrPQGJtT8oTNoCBd4di4sk89WhIp2aOd2xZDKH3UfQ+i2+YfC8wzeyaz/p4NDc/59ZjxW
77uWohtZXlIQswoxsNcnQwTDodZqEcp1PRlZX/Z7c1ITYae+nRYdLsU9PZM9N9eDaY2XXI2E2SdX
tuHQgrtAoiMGip+a2brWNaAN2GkheFPkERX+0v2RHsnRGxhIDLeB4mW9yEnXRwAonDf8f3/CRH2l
yvdoFpyvx3O862c2+1wsCWj3XodjIfbsBlGF29syvBqSMSXowGPuKiYO/Nu8qehZ2jhMuZRbpNFw
pp7GnBfh65IDm6bLZeJgHC/Qnwp5bym6zB1h+FADT56tQ1Pk48r0HL5271YQWtQvlq7rymEuQfHN
5u2aQa8jIUGRCq0aeBEI5pqVhi6EnXMKkfo6OjmMn5yOOtEusakkW0+KCSkDXMjjxHGTSqoItI+5
Uc/o2ipIcwFAqyW4QRN+kqmaKU+B6yF74o4O6zp4EwOVeqQ79GUDylhX5+5xReBP1uHS7Z6NaoHY
Kbl9yzmGjtOza/mjkEva6oGUvLcRpAWLONmYgH9ccjijxmgX71JKTE/g70IMB6WSks4AoCNxICWI
j9IZpZLbPD6CjV4hWY7W2Fsksm0yqeDalSOSNqXSfjm/G7hD8S36Ox01a7sS97dc8I2Sv5RYV9aX
TJQMEz0cYLKlo/l4EgK+TfCF5dnohiYYic6IFN1LzFW5HpgtdX/GP62WRnA1SwwtDpwiJagyd0kr
xuQPFExqJMtseAaIKPN6LqmGoXbQrCRMMzHFrnEVNYEO+0KWtFn3UTQI3O4DSdK6eddhwFTgLmlX
fy2sULWNQzWCAdtqMlZhw81uZ0qeTSvUj8tc6d6n6vmuF1NP6GOtGq5wjdr0MYmaVz+uH2ELg+uV
KSbV53Kx7a8kYWBkpvO+CfDmNolWew7PusCA08Hzr9vG1TufoFfyhex5tq83nhdyIWi0w141U6gR
sTC7xy3cAJJ2jrk0k+MCuUMx6xkmedssh4BFcVPDrgHqiDy+Bal7Zjg9LB/0/xGhhiCIf1TEUakv
qAKjx4PDv3xKnyQPFk0Uuq5vDFmxp8LO3P5I67eYi/xEcchqfqes+YblujTvpKNZ31pBQDaNaGqQ
9Obez7V6L86tTJ7KCvWp2SxaWxK6jpf+X5BwuJv68FqKO+N+ZV408hGNX+iBqOquVcPZYE9PjIUK
62lbXmRi6Lxr6Y+KoA/BJivaPvvkm7IZ0pzXqodFDte7JpqngfOebpgbizA5mB6dxjXzFq8ysoIS
TPeqhuiP8+rdjRA9iUEKDUQ3jB01FO94+xCQJW1Hy7uFiM3OyWh9KDLSAHQmCKPCHVyXb3InmHjx
htpz9LiZee7emvvc3w0FEPCrLz1cBH/TL19EpmQvT/R/6XDxOSg+9t2uO29/Qa9sEip81pEHj4tg
remiPTUniEKtyCpWBjfobecIljxuT2oh7inmR9t+Af9w75301Sg5v4lq4B0g3GpLHWfIPYAHxGbe
lXuZf3I1JNWJfbC0E8nrPCKB4H1OyUpgZCZCcFIxnY/OVxZnVZdupHAFvNQCgKdeCF2adR7TJfuP
7+pQLbbhWSzgewlrSRDdyUIP3i5iAOcNda6VDjGlGNDIXwngMfpRRW26ODfWp4zm50f7G+6hIHHh
ENU2G++K55LTS8tXsALXRdeGnIeBrfW/gMEcCeSfoT8Awyyh7jf4v4zWhOLzTpxtOnXa4f7o0od3
hO6rhleXHjko99QpYWN1eGgJb4wPTVbnBoHAVBwUXDrzuZCa8TqOd+iOlbLqVtsuVUfx5QTxhec1
uQAjknJDmZwSoEUB4BJa6YGAZTVNoPVQoa+B0ewREmXvFzGGfyg1+6FiNH0KAEv0WUMgiRLEGMBQ
qqt7/BQPARCVHWEdJWzNL2CKomnZBFN1XZGjPRH9iZoF/VWoCo2h8VKWe5AdOIuux5Jec5jxCW4x
Q6oAjBs19DPTx7TjNpwKVebPNRV9oRbzHKGnXzDNHuyI+GYlsJHLA/Je0InHAzlCcVia8dYYh/ZL
Zvt9bJoIFz5FjvnN+Yw8uJrhVh1ao94K/BfLnCFsm8+sK8aQPA3VVXtF/jBOJcYCGgYTPzKlkTap
O1EF1YC2UQoCPQ4ko8M3Pn77/9QajFYLayBxGFD2yWjXZQPCJJoTRJPlCohRUhzaxwI3nKnsEssX
JVMUwc+Ox6shB0hAU4643igGQ7lwhDQ47pxFZKZ9Jsr8jGU/XORFk8zFZMMZz8CWrrAkiwMr6aUp
UlR0WUQ4QI8uijsJFjaC2PdN5cthXFhrlsayi9DYginV73FQ66i//Sedro162RYvLKY1WkO/pNsO
IiHntbADUIIQMOG8/4/JIAFDVjaNt1/lCyTjLFMtNqaGRegEiV45AYY2ekBRcSM06QXstUO2MnHe
ogKo9YNm7z7c6fgphOBshRWxuh8aozfG4mq2Gioe1F8fOqe39MnT49gJNnc15akDO3RPNzSF7Ij0
L6PTFWzxZlDErj011PS5U21lh3mZ+dRtBufwm6X9yul7nnpNexXeD0+hxjrma9mlKo1GVk6XpK4F
+IbTarh5guYYlaz6nCE5FaSX/zP2BxIufH5EXNZQ8P/Vgfr9kZl8T6Zr59zi4WBaQ5fiG7muCBva
IlZfNa3yhW+hQDJ45/HX5sUsT6mSOxOr6VG9clyFRtiqcQAdBBFvP7VezqSC/EcX05dAkQEWm9ek
qRDARiYmNTqHfQ9v4+Bt4nRUPsaxhi91AOXiy+qrbWge5r+tsudLfDHAlhxwiFz7nrndlvNS/Osd
TYmfLHL5geuL7jTkbD/TDh6lJ0YM7ydZ9lEBDl71X9pS8PlFLcpUSUVm6M6fOiFigA1f0FCWlG+k
RiB7KYQJUXAvxXiC0aFnI/I6lOY9B2T1w7/F5rI4daXLDSdNLTJKR2tprDPld245qMtr7ySiKVj+
jdmdhRWFeIgUHNZfODSUf847OaOXDxRKMa6Yr/cRMu+07YX6lXXBW9iBpwBsQ8b5bUqIoTV9TZcC
+05W9DfMY7uy4dhRbhnL7NYmhbhrHl+/p7v/Pm0q97ZP47buxtH0D4ydDxrhVtsbE3cyDDZtZgLh
XO++cupCKzkOyOpD8VtyxgsBnVMXR1PPISUIJXXqWJYLxgwG5Yx6s1KPJXDtF4pdaNlOAFXUOvKq
Iwd/UNt3P66cXdMhqB5vu3kKWd5wnGJsX46RrrZ98ptfCsz7Mthml5Ali8s3u7IZlguRMiVOafpH
0sE1kLtmoZ988oeVSs7bq96L8pTyu+AYY57zEdZew4tfdZIR1xW/16I8bSz4rG22nP2ndB1id7rr
8XsTQp4emJcq5GxdINuyzHhFtIgdBjvitWNU4crCcs95HMZN8FfJjnLNU/8H4JxVeP54El6+x4qV
xqE/Iza5mbQdXhizftftUrzGrXtbca2VHyQrqXJY8H13r+OtZRqwDHKWuir19XJZBjXYm2tmKZoC
PR2ibaRA4OFYk7Z/kr3aea60a7Z+4Rl1XAgKyN/4xluFRDei8mbmDp0RSvNwL2s65PGOyyjLLouG
svD1ILNlBJuQQmX0xOaeaRE1ByDvc6RFbfbhwhWyjmZk2/pfFqAp/3E3rMknw1rASu+g2+mcKEhd
zpEHTGwaMidgh5vcWit2Usj1HPGnYn6nbmeE7+4lhK2SvpMB7cdjSWDpUu9qqgz9prN4Gis5m+nZ
3chh2mrZi4uKqpGAzCyNNxhX96llCi7Xz0lYw5rYfOIHeUowjioSaj15WlPaeutOweJWr0SNj0tg
z5fBxgua+s1plyH9SyQmw34wYX2THnY8A/Q2AHPdY5rJDbZS/qWreRfJoRnAcwtcIs7VC33uQlHB
DTKw3gT069vOf3lZbhhY0lqReVuYJawhFqAfj2lDc3/uPBusBMIkiMcvNM6XiJ7yM98OqxfH2zX1
wKfoYk4E/kNizLRBZpj5kiv4Il6K7Dm8Mw/cZbF8l5evyhwDCx1JF/BJlLVZH4jDKLDjcOhG4I7h
4C202r0QFrOKKmyDCMP97bvQKyomYdo7oIzGotpf0uArUuvjX4YqU+r6NZ/3A96jVisCD36ITrIs
GO+VJ4iZwONPluFjmCqbsyov6qsmiJpXOPujOtUzGCUT4tzA4515ywqT9bI5SFq0Pyqla/1BuMl+
Z5xTiLESoL9YmiTn0BNQR/NHRve3wpCD1gx33pg2kMrQPqWD5M5ksigPLo/wm1t4+uM2GMDlbGmm
CZ+QBZAK6x8v+0Zd1F/CbiUZpHlJRJMAB9unHG6nmzKLNc1NRrbjzrRsQkEYzOrvUqkeYE5TvVc0
Yeq08Utmv8qY93/Gi9Bg5/3BuCkAhO3Ufe10/kc+/o5jRfEr3iUgk1R/b2iy+5PgvgpJqEBgCOZe
R4uN/UR01Y1wlizbyHz9xUlTZCXizIpO2nrMdPjycI2q1krZyDqIb3Dhdu0HC9o54fKv8xMlJ3YP
dkRIkxdpCzI4VLioPbpbj4P5J88L3mwZstLh9Dw2biOmz8IN+RlCSUTC537ik9zTGcPDDfqAvatN
BUKn8vxldH4DB4MbeTRuApN1BnbO+oV/UmDnFwWryWbnt+u6lMmpZt5I4iK7gnycBhnAMhotCBD5
VwXUYN1/n9ysTGE4/gLn+RggOdX1FOKaWmhXwYXDCI3XLgcMLvnQdYL2x0jvJhcM1B+Q/aYqGZLd
0S6X543dR3K9kKtb4A1mbPlvqSijNJEFbz/WRzzH4f8VRR1s8MgC6ZRWQL9j/TjqsdWwO7TGGHww
PBhElODSzyeqH7zpsDYYb8ZDR5L5FO+tufllFDJ+g51YDXgygjavG+7hRNmFiOk722LDDA6aXca/
ekdH6L7CnduvH5k9cZ3qAxxtW+eEDk4vXJ8CqcCPm8pDoBJCi5nRGK/Jk6565Z1oNNuc2CUe8lTR
vO624HF5oypKTMe8PkdZC/H7wMNPCQ0IsbbmuDC+Y3WtUPzbDOi9YfG/1pGaZ8OkzvyYhQjZb4OZ
dKbLygFvORX/zCz9rbY5miF0yNorkT+8ciwq4WUEk104XyUkgdGW7nIyqPF8gJLJSW1/hFGrF1nG
MSWOl6kmvLvJVOEJkTNCdy1F1rRP82LPRi8qRkcCGF7/a0cHLczTH18dhZYg8HMLxXo9fqa10wuu
xzSb3548BM9sM2oalGXj1XYmF0sFTF6Ci0uPCI5s4ai9ycJ7LZbEEX+mdP5d+btVeTiSlDL41kFn
0A9Clf3mEMEqucRE+TNaw5baQwo5PHWffkoU1yU0OHL4dhsXhNWrGBekP1om6RxIdhPkmqejyFqL
xMXdw4AJ/e98lF4anABSu22fiu6dc5d+1ee0snWaMQQgM9b1ckkAVCzhtoS4ngkTWN7cKQo5DklD
XtP5UQ3UfUk0TJWOYGkANet5TH57X4X+BtLyoi99uVsO2ded1ZqNE6RwaypTSey7TritQ1yE5kRi
o1+a5CYgy09Sc5MxQZwIMiCxIbyv+zhon8sK0jRUmOeJH7z5ImiUZgShmNCtFWQ5HM5y1pIAClAT
SzI5yReO30udzIfEW+Ia/sN7s15nIcVjs4ifQ5wVbIazVDPt09ytroySU/040Iwt98d4IAv0KvbD
eL4ESBF7X27TmHDBYc0wEuqCk/lZuVZcBwzEU5wULQxiVr0R1dmcdwgVAto/Gjv8FjcPz7rlQpW8
+Ijj2WdDYKG0olXLAt5h/puwsV+SSM5MejBazZqWrYhauKIULH6Xs2JOoRv9VVNOg7gQGlpDBEQj
knNHU4lTajXO7Ue1l7Q1hATsgoF84oTjYjJTBO+WRo4gfs/oCT3FgwBvpIGr83mKwg5+4cADH8/I
+W/zwZtFSIIyd5mJPFAbF4KSkbS/q/Z+q/QMRH70B7/fCygrlFxyRrKLd7U8nkHYpxxvEHtTyIrg
gSAYl+WhLpCVseqrbMVI6SDnRI72Ge9a4/ahC62HgheiKyGhxZg7EH5jsqVr7pCePyvryrg3aOol
3axo/oyAs+Lft8XrvRoEi4O10Ul8D7O7RAs9Xh/852knevUFnBk7oSqjtBgUtVmNGRxvYiUD1ahh
Dem/nbhxM2xctKcfFAUQ8Y/ENZvOGFFDVgRVoM1uvPf0365cBxcQ5/fzgu7YbIvciyPmW5rzu8HA
5LwBxiHnLqy5OCjd0TbfbHWgxcmw35fc6srofH2+aNBv7wXUDbA0gJb9GuvPi5kCMTdvenIFWUQJ
GWHSu+1ax869J4JlXwAqoabUUkAHYS4zswATDDGZPML9xisXrUA/46yq8wzzIWmJg/e+jy1OOFxh
6PqkYELCSvvtJlHQZ8p1mjcAg96ZvnRrzKKRmlAH2CnPfv07qVoYJnZecgx0MuU1fs1GvBCuqxPH
9Ba9lw1zaBmHqwScqBagbHPUmWBuipCQWwBCnxXZjj4lzpxOQEAZYMQt7hxw55rY2LJAlfrodtSN
8+YHuZ8zv17A+dIWUwibem68wHspXFY/h+sY1iiY1EF54UDNJpFTExJGrf5pHl3/jne0j5r2nL8J
jdj5IttHo8qGiHntnATdVGEo+evPV1CZo5ck5C1RtJ0pTNB8hjkCcIhpJDVXqw5kilpewrmiai8t
BY73DtC/yKzdqqsKLG7m7SwHu/mA2gDbCE+z8Q9kqGcaizjRCYBEB4c91vd7pUPbwFkHtN2XQ9zg
qudcczJi/qf/0vDwE3tZWvO+C3L3VjV1hf3uuvkdfowaGu40NYNzkwLK/I13vGDJ1hGlEqhxWJXX
2bj3wnjD2VwQ+QK8P+M3OAENAtMNj5VhPYhOtdOOtXnMZMvpA0DiMQFQ+gV5nvRN3DoMQ4ogTDUS
5C1cJNcwbIwA9T0MOTOqsZezU7T5BUoQB8vda81D68+x2SC+9BzrhsXpoX3pGdxTwDiQhGpCeieT
UizADjZ+N6tdSeA04KbI9O1KeKO0Op6OfL1q+YzovLJ+FVI1J2JZWvCo9rTzbqWeMp1VjJ4oO6dq
vGN46obmW9ALE0iWQ+M9y88xIqL9ScTxh2Bvi8WK6VERYzdy/r0+wWY8Uo7NKfSH6i5TGtlKpcbK
G+eZ3WF8ENSt/7dfLro53L0UwK6uaenrA/T3oEfW9WCpkhdZBVi3/dfkpaqvB+8sjS22UIsPvskJ
S4gqvgm+sHV0+s417yjDRRwTAscjBoo8c8RfXWgCW9tyhgR4YoTqp/G2sHtz9kRX5AhPFVWrXGoK
niToCWyIXurEoChSKvIWg8KE4IkSCZQ2+ZkUr81+PxDdEcJc5zjc5xMS5CWEtqFz6Gks/PSid1NC
cQUldlwCpWBGWZTDC1JmD+lzyRsMaazTQfI9IDZWkdks9is4sG97HmhnvPzxS07wSofBIngCwN+2
ARlsHt4adSkWwhqBfCUwVrQG4O1rRlWFGq2ExN4T8yVzEzYfMDTHKSKsdqR4tjdrwZoWhS9k0WxL
9Kh+irbWXIK0YwCojIyrseME1eOerCuZIYXiwqu5figUsewWLj0lpnQ3tP7QJ5mjRZ3pLwNWSJR6
K/RL17aDzPS9Ldg5UEdqEbxYdKTBkt6uzSkyvZKxekjFKI+AGaWr60kloC3qYNoILiQf3wYTm9D/
hHXi729rXFItwfcTRA/zOXBRgn1Zsj3BBefBrnBgS71rxUcC4cbRhr+PPOTtGanDCNqLvw6eV37Y
oeGMtfjwBwTL/MSabJ7d2pCMz1OIxp0L0USadFGuM3p4YIw5Af5sV6NchnGbRFdhHAxLEfWgySRL
ede+kQJeAagXr6Ch6CXjJ7p5Pc3uTcG79NKUZXgk4pyBe5x6eEhcgkrmOHRUpx6eERhWzemEYpiX
gXb7YA2hWM7XvgTFo5Bd8swKuy6V9Mz88LRDYZY4qntWgiSDHG9OLx8AbIMswLC3PiniY4WOifCc
BpLJY5WTtBQkNnFPPPHtleJ50xbaYWX06sywzbFasOQDrRLtI0n+rh87L7ATWHIPsAYaAeWF8Wje
EM96ZMCaYdzJ1fm+Sq8vCTKW5E/R6+6+H7wyctXGybXyfftnStp0wSF39Of0CavhszzibD4tmUHF
DLt54kIj6TQMUe1zc/QYpSwTYPiaA+9hxacEfM0MLdODFcSvin9Edvga/FTdsimGNec638tvifdn
w5XdnWkpdHZyp4NXnIO//pVHSkGEfTX+OJZRSo+9ntG0JHhmLGEUJVybQbq1/SfZoy7v4Z4PqKG8
opj14p875GpvV+UV/SHmfqeXxBfSLWZQ2stRsJzK9LzaaqtnsFnwdB4W+pXK/hbAXElagoFE32kG
xho0FufphYST3EsOwG0O9MsLfbj6TN46h7NTPWRlUDL1IQav/vqKfB5aqKcC/yXVChdqU9/cyGoL
1HxPaJD7sGJJ4zWYcE2w4uISPQWt/c9rngNaAWFix7R/m4Uc9maPX1gVeREZMdwOsc/OyacE4K9e
t+Kl9SMsBhs/gRTI5tlHCoWfW2MWf3+grrKWYH2gZVoBBjbtVjxRXQ2l377Qf1a9sQ4xOZtTP7FJ
AF7eGdzCp0HxVOLnQ1VWJ6LlWRhj3NSTKpR2UTUc4Ic4WqGPf6bpcmLQ0SZY4UZw9mReamxiI5FQ
CP1L1bCI8MdYLjQVw4OKmF8cUglKRbTkr/um6RHqZiwwGWZL9lRxUMFxr95EwiDJeWjO6bbFHISy
JNYxQdcYUy3vGwDfwtSBHBdQ+PHoj//LgBB158ajGbcKAFl4vHydsxxUDfXUHJIw/6XoDx1M1+kc
qk8m2ReAJfeyxhM950fYqMrUS9FMprFsUfk7LrJdQ0s0cn6fYLAnD7SCdqzLxWnWN57d2UDf5Q/q
ZQbjTFVlAsAQ63vMVTgjnbgh4GPl+ThHZS6wsEivleMr6mlLi7ZX54E+XZqY02X3hOK/24Y6ny+R
afsGdPX8F8zgMvnYxpQqgk6o1Xt6IiUoLgC9Ik19LufSnYYC3iAZJnRyM15wMGhacyG2mViyNxER
vE7tcCgn2boUng4cT57ewt7ArzfBOuns2AXF9SqDqladVINB+aBd0ClPRq0LZrEmU1o8VxXp10D6
wuJZ8jwZtNl6Mg76hVXg4HL6MCp7U2zP8kq2598ujniN8N1r7g9IsVFFdju80kg+ikDW08uuS3Oi
1zs5TZAetlHkJcV5P8/l/kInTcICncPFzx/71rAin6Awxqt8CPlldXmvijrlweT/qhZcIiELC65N
E0xSo89y1aexXeG79J6kl+tUKSoE//ZQvajHUiO/BCcIVL4jVzpcYlzDimx/fdsOPI8ML9XA5wv4
JFbZC7m4OAOWRDSpIGhLDL/jaRXpiubWgy1yllbtpftAcfSZJzE1mHNzd4GUHbgpp9CjssnMl4uk
TagWl4CHdZcqnsJ4dSTiRCiI/9BitElvOnYTn2oN8o1MjzrfM7ECS8/cadethhmfJ0eveH5EHPYH
eZjHET+dhBr8FUSw75UfhEEtbmyBLf6f0i2+mt5W9FLgIIVxQO+apMKY9uj5dIXyLwsT8vAPHJ9L
kpM1b4dUp/ZsnkKiH9MZIMXa/Wr0IvdA+/cBQo1zoVYGq9JbToO28CZQfEN0yd768DUTxzI9K5Gh
qkRxGoUp2bcNtzJkKDIWnksdRyAiqVauONiKCug/P2ICF9gI1e6srD+vZTQ03JjJyUZ7mEqf7/g5
YYfdUCPDjGoQSNTc/awA6nPUndyR6o9HRfzixhCpl9sRYGyijU/rr9DOeS3VrcZeyvglLvR1+tsT
mHMc2T0wWCVQvlx4ac26IRhiAPLhe5yTlSce9WfxiRhG4j7maOvvMgoU8bIHHBLTJpupxb3VQ5tU
t8xYZUZnftVAxC5viMU2nx4Ddlzfp+CXkkgy2lP0kSyY8IxHCbqZqg5x7Uvll/A4uWz3ImrIgX5H
tHlkg/psPJ1WWgVgdWeAnMKEmyQurCADqpzG6PX/ToDSD4+Xjb6mvtWUzLhOlg+eD4rZzgMeyhsD
RIh5Ru492OZMIrgpUq8agqeFl+/NSSAhxLDZ57c/ySsUsgaYs4y9iqYOAM4wVheAhTFswQHxK98T
eqZakLL1ce3zzjuFfhyPJwOq2z2tqHH0LpayHFcNdAEykrmvCK+5IicDosBkhPF5JdFt812tAPiC
+PG15PY+uZZ7D4kZzy5HEKq1MNYlE1qYn3VaK15nLMnhSojoM5MdLY98UkAABsvPyl/p78nxqO46
6uksSgiRrRYYCqzcziNQFQpGnvKuII29WtuP0kToVThHm89sphbYvD5RxVBvIyIkWxRFHtDJ7/cJ
sdXLWIRYYnmoEHfnot4SI6BCuk02qkO88MI5L/ecSDPQQO8GU3wqTRVBUve/qOtlzW561P3w2joy
mQGMD5V1hrbCPoLCX1w77zi4P+DCuaJ4r4PqMDvcC6Gqcb5YszbtrrIpeevx4/R41e2Ym3o1lAo9
O6gD++OukqliAp1QBlgs5SJJXKX90pinqpJarsDJ5EtOY2h0MMGJjMj6cWCoiH0yF4Mm56vSMkG3
92hvOYR6X8dkBgbfbOnOzOxjW6/EbtdbCogRafhP8EBYKE+hrz+udd3MKNv7fk9FJTXFlPnvILsO
Utyt9s/ErI8Mlw/IIM8S/AxOaWxV1s6CqEhDbOwSS4TxsmL3BZrxw4DpwDYeapacDcjqSS30kyrS
BSOMIFPg22gNCrkvZ4Ibq6U1jTxTPwKwhMVkzDoYuTDefSqT/+L4PE9g2qrsGIn8EtrK75yzNDbl
rA3HFbygS9O2GRy/aUkB5rdeyA2TPLlZvLrN3Xx0STrLSFd1zbCBCF932wsrs7pPnb8yVTMkDMOt
8TLIiloTvj/LAQ0Nh/ezq7JBn+H0cX9QoxwEQ6K7tdNDFhMyAhS23KzJwf8nnly9Sy75MIFeQkG/
l9Kfgqwwre1cQq1Z1xqEJX8Ro6qqJo8B3Bqu/7JMtfb/Tfa25oZQ3wjpNFu8BS+eZ3g/pDKcM7QM
wMAlwmvbI5+vwvFmWNLQRIzxNfj8+uAbyYRwNhRMuFU6DS9mFEoGHYluADwm02559Se+5wZ5bHQR
oI/qznYWEYa+i7zE8j4vrhN2UhKDrL7TzpH4dtUZ51NeZPQFXo3aVLk3dcSK/yeUSxTVcfeEGZhX
5g85f2SNallK+6B0mgmWc28zgeOqbIu0iV1bFN5xVuYd3UbQsi1SQ6UzYj3PYJetq/l1jGVJkKXl
qAF4VEGAKnUH/3JeURXsZCc/en9n91VqbnrJ7qykKcq2Fvr0FCHfQZBVUycYW9BLEoh4nBREk+mF
pwDdyMrE8k2WSbt+CqFmMsREu/Gaf5N4gYOdRHrte8FInsdpcrYF7jA/UwTnZgUn4bxpFtlu3+iW
iSvTrypTrGBFxz2yRLlNrmZuzOIw+LiwoYrY40aoSNmw/XfMGH8J8YL6z5ubUZ+0yNJXn2S6rYLL
dX2c8+f06pztu2ZMWDZd9ZBQhSi7A3ooBwjHkUjgF1KLK7S7M12vpaypsXIpPcwLnc3WrCH/rwof
HlJIU92kpGuanTYYSZG1My3yqRlzzkYo9w1a1XeIsftIUXchGS6CYQxM9tSHHoY+J3esBYqIDMap
m5wBZpI4V/pNAoCVj2sOjqb4QGSLwCVaINAQIxrg+PTYeNGrEbiYXQpcBsPUsaRs4rEKE17u+d6x
6X1pLCUvR2JfjxJvigs8GsrB3pljH1XGsjnV5/OraZ5D5GwCAo/uZL5JvJzkYVEHdID6mWaw2jeW
cTu67rj9xCwq+zt1M/WFcH74Zb1QiKw7p4bPSkLTEb0rmsyTxcrZRhaNgBPamie9QpTmSSJAa4Yy
1tucUetyHYaN5xAvnKWBAaeY6mKsJhuOtxZySZvObKpsMCDILvPt0lHmuhnl6b0B1+O6mKFNQoEg
IWq7tszGzog/BQc5TR6OgDH4dSrCUCKsE2GrPbW1bvBaZT2l+xjYd2WsXkVsEI2CEa3dKWkuLGRv
oy45bLtXHVBSnWByiPK3fw01wWlpWNa0a1sU88oPgwBqwCUQ5v35/lIS+lLr8dD9uYkKWhr9E7Qh
fW7kAydhmS7OywYArizgzQ0ns1TUM2MYbh17usdIxvXwZuIEn3qb3GwHtB0AFqdonSSEBxtkSLpF
HYYWcnZoTLQTs40xtOU2Q6POKChxEwjVHDKUCgK2iYo1kaLywyxCDuiNOjUCDdZq1IAo8qHPz6Dc
czwtcXa9osaYKNB/cWX0Lo7HjQ6PgTX/07UsTlXQTx+W4WKEW7SFUQYv5U/7tD5p+52yDRb2CVA2
I//3UvJ3ZNBkbmMAZpnBXyMcCQM1c+Qg1r8fP1WVzUYslKlNxghSrQZOEFCXonM+YOp3e3aeBNGM
klbZvPRidB8LNUZRfFW7CDzmY08nQNJ3FzexE2qptvGqKJ6cNDyK17n84KdGXp7ZhKvfiN/LL0Jb
wY71QeWV3h3dn7fpmtSiZM9ukIJMT7chStXe3ZMP5OJfVZV8gz90bw5oA4UmwFfPERRtKxoNATON
W2y3X5G5lXP8c//k58xMv/gXveG17TKFrR+LfkTxveM//KJ4K0Zo4kV2rKk61lIx/Sxt1M5d1eak
paG5i71XRnfZCNrBQwU6XyxUFck3surZRJ0ZfNVjr286eGWUgMSM30hUXjTGwjO12hhc3IMw2FUy
pjgiUSnD2Qm1N++QKLhkQzFGM6CpEo/1V+dlF9sbrVdKqM6H8SNMuWGAjhcdFk6Xgw5w80Ekzcop
jgAzSkViBat016I/2knffrJou9QvRLNs4MjG/QXzIPrD1NtyRJzrCBgc7Nn7ELWac3JsKui8E/rE
FVHjBCyRKUavg4J7Thxq9TXi2DkvQBnFtNlBv5tqtECj3BVumjL3kVJwvxRfICK368TPCTs2lzKC
pPpUda89E10vAn8K2mkrc0JNFDJ8z+NPOnS5Myr0l86F6r8ERSDQ2nt5h/0Y4LmW9BVAYxIdBs6a
lj3GabqvS4txVkZVkKLJs5cCZ/iXrHu0JrwZuy7ofEIi5R7i/artoIHXP7IvopwYXZQqIC9OjLDx
he7tfIf089QCwF+9s+xYyFzsZXJcQlLLBBB6Z5ADV314xcvDb8B4x4i63f9mQlHzWN2gavtKSoW/
F5sPRjm6VvC+KqyUts1CVZfVwnKmK4WFPLtq/7CQQ/AKxhxprgYoFIzkBGnFDSnEjtdqNSgLe+Lx
8ZJ1ysGVfYHbyg31qnt/Fdn1CwWLv3eydTiY+ZiJE7N0L7G8kubdAvFqA2vqEB85UEyxM7P9paTz
htQyPyoolMEjhmx473m+U6mR7RwcVVdvp3q2VAuz5pA5RZoB00T7WtYKR/AhwsrBWQx1m8KDkh4t
r6dBwpiV4XIFabzIFP36o2QHL9wfZEfSEqcMCgFcRTJEtnMDMBijtoDzr4/y76n5Z49DfVBKjF5Y
X3C+BtaoAc7XtcPSapZPYtZWtr0TOaDVIzky29uAFxozgcHHiAluKyanRGQgmPnuyiU2AGpKGLry
fzFBIREIxfB+4d6kmDsf+cd/QTd41FNw+bMJcjsgdovPcdBxouFaH57ceIIwv7Bz8khjctRREJPZ
hHPQfotkEfDlrFyvd0quS8UCkSSFgCWasQtlxQiV3cQUDtCr0boB/MUf5nIsv8oBOxGTZjNa9kF9
5Rk3rPT2pjM/BGoVX9+TiV5d556AA/11QRW6FTCY6IraN53PdgbJgWUbsHPqpomzDxJEWKNhjAf1
uJzMCKfuIvHlkR6dcMp1uXeoHE8EPYrg7G7+FN40VcMnwzeRNmEft+iKWPCqvOncNQ/pX6vkPCpO
I1teH5L/4nmgS1an4y9yAbqL8FJIKtT8luV/ToN4CATSFYnoHYsekl3HpFdN77Pb8jnRMkZ5p+PH
XlKrnZ8CAkErxE7m1yimJhnKYZFbDYlyJAWxVsUZZzYQ42taTOF9CRbHONF5GH3WXHOT0ntsL29M
5sWMWzcLtNcKEx8+vcx4fKu5uvnWgXkvrqe4MMUL1HpXmKxbg7pG2jrXrS6aoebJCcaTBO4W7l1X
zXzQ0vbvDkFK0Vvj2kVPjP3VFgAhIZLb6Lwo+yMBh31upmJ9kkgd8W6Dbi/K5N0d85HLSCP2ma6H
F3qJCXdCaXufyxBA+hRIZwdyENOTq26/wvomXhG2PrxXtFItcv4GhwR/xVLBO88WudqlGhVNTLu5
+kcERe5sIniXDX4DkRbOOLfnpyxsBFNz6JW0A2ciMq1UywPzvqCZ137RxBFjM+td8hh2nVG2wQwW
7RLWIcXoMjdHi/vJxEID0zBck8q5CzRf3aCAT5gYPRS2ZZ4ds/X8dTR6dDPJPvG2jc6gVd0HQOav
DAU7bFjWTm3arZVRcEkWdTnl6/IsKz3Z8JHpOloRrfcgM0KkMWF0vOmuD4cfrwaOniU2An4aRFlj
2TJ1sSvuoRCy/Edi6zL6h6vsqYHY00Oop+gLVWKm9bdFaIDSuM/qEpbHOBXnE3+gXmmsBqYwlN7C
3fTmBfHOdO29Epp/8VB6EcZxfgzKEs/zGEws3VrGEOnkSP/Ez7Mbjzpokk90W8M66qmuISnco4EZ
UOanPnAubGvYsso+Tc27DjXRODtrVxmOOL4cvu50iTedO64ax+76p39pNm1js7GV1WKppuElDk2q
6CuV9Gwydrg/PKiTmEgaic0tcijiDTivhylT4ERShQkM9I/A7t0tB68uFLZpMlqQGenF6BvFnWfs
6sZ3xOpyH1bc+NdStufAiVE/p3og9NISxs63sZ+Wdqi2XVBMDw2cnMb6RrVoxwCqZQ/aOk1SdT3r
phz8/UBBW76+XNoTdjgCbiyuCWLkvinlHzjlb3ZKs4c9o569H3dwq0JGdsQ51pQrhBCHFlCN+spb
oxcEpPc+TKXmEX6LYN6VTxO+O1oedjK9O2d26ehcjNVfEKGOPYyFrgrrjUmdXx2kyAPcFcI/Gwpk
KX3fimTScI4MH4H7Pis+NaQUwtXwmPf6F8zIjpMgTKr44uharyEomJedcKgW1EDNNq8wgboC7/vv
ZB+cf+0oG1EcTYTMle+ghsMsvGf6caMZoV6BPNMtSmQXTY5QNBOM4Vplu93JV+fbrCjCT9AlQi4+
v7p3aleH995bvoTsS9SnKyMmK4wT6sQLI6Vfmp+CHkyyFSKGLnoaL7i+adJ3XS7at5CfcaVnzGAy
X3fxRkabc3rA9albOMP4T0G7ZfQy8YLvXdTqAuWyrlpR3NGSi3RD7fXRRTcPuzUKGZrkVx3Txd06
W52p7uG+H2O2EfOiKClvJ6avD822LxgWmfZ/mkrRh5DzGh9tu0oS/A776i7sUugIo22597DxtV/I
TKHRuPmcTGOgt6Co/ofvugAkuS9MDb120/pz1HKzVPqVX+D6AggdhElNsco9DQbBxIF0zGfi1fud
dXyNlyQDrBhFBO9t/oFUkr+ME6yte28Dq8r6yUMI8ut50YzSh2aymfHrtZiURXychmpjQenBljGB
CeZo6WrZvGVUpbE4dDKZQbFLH6sxBGFMvUHnQMM+dv8X7wafqmOe9OMmWJJacX4c9+7AT5FGRvwk
nsxZitkZo+2sI6gQCRx5cJu1EW3dOl+UdUtsG+QmovsTQt075ziFKeXwiRufhQiNL71CUhhJAYvn
Dv9Y+k5Sdr+7oWFcleJKahf7weQ4LBxpIzWaga8OGoCDd9uKrvGA6zDJfMUT2rmnaIrHwJ5qXrpd
7PYuKRP6WW/SLGf54RBJJ5fvhDb/Xh+C9BEQNqsFct+l4elbntEPA7Kr6in2wdVEgsnf8tMlAYe2
BTmWIE5mBM+cdw8BxDEKKr6JvIDWO2VYBnTw/QDnKyoDd1i731nL3mF+FEj7yM79oIwcH9lGxcEF
j17tRsr9L2bu+GBgzNVIZOYcin5BFchtadaCCXnvz4lNi4RBmMBhDE6wLk9Qv3LjehN8hYkL2YQV
DxUpl10MuDR1WlivCo39rFx3mB/qy5jvaj7aVmGVDmFRbTc0q1/IDevI6PLfhC4xt6oojsy75ikX
1NSIMJFKTrciQa32zKHYkgEcbFq1DUvntUhPGKX7TCoChbdxODFVbcJClUJlV1Nnd28ZIu9C0ufF
xov3dXK72i9xZVaHr26SnoJP1S4v0QnERxYvVpit2dZYjbkrI1s2b9yMAkGBrhi4DyKr+DCWLAoV
GQWNAEPloLTagG/1vEeuG10jTS+Wi5eZ5PZ0AMuFvoKRFhY+g5vTlmVXGZTiY37pjbXZTzfT8DPv
aCQ0wbAkosZ3P8jwfPD349cZEdVO5x8jZklZfvhoHr/ys+gSX98dyOKYbITolmSlg1cAcOBgOQse
3vlTjSNpxFrqh7esLb5rwBnwk5xmOd0MUVsnIP1/PS5uHkwcfBLUeg3/W741ckyGQXfv516ewEdG
AUb5twMF2mPBelS1uvY0h40blp1hCFI7zYch8xgwB929qtPJLDBJHl679PmPgG93S+6IdQYl0qiT
90t9GGgY+QDzcG1koTYceOKpl5s67UtrA7Du+D2CL3ptQvJkJ6biYniHVQ0bUlqfI58zu5WEfZoM
nrIAUd7i2ftj4SjqMC2At6bPqIbrlGTrz8wilsHZnIphKfOJ7v3ZdbOgOEAdhXujgT60DkQ25IfS
oBUISvzpuammSlzGsGp0d069SK2ovQBdNgXQ945vyt6DoPhKcLBv4HmHJL1fb7MttuWOqdlwJl/B
dqQMSCKOx6plhmgQNIfF2BfBs5EEoLJ0sA1xvi+kSvByNGhm7o+qDBJNeimuxnnKvUE5UWWVPpxT
qfb5d+VywxqH5b8x6+BCBOCREt7yL1z+IlWNF+lc6m00escWUjjmZv4UL6wJ46ll4PBMqrkyvVW2
QMKaQHmB8qSGEug+v4ZitFSCYyC2vdQR2reOkQm4bj2ftvQzO3Rbs56bGgPuV12WftGkEXv+PNft
KnvX9wuSfJRVIiUoTwNacXLOqYQ329iMGKPrK0zZDH6B8QYf+l0ozdl+ZNT4uxuIRe4qdLrAcGR8
UsYNZLWYhghpBjej9uo6zuNRwupg6pNqeGHae9OSp8SwRdD4BQPUeHK4R2PTO7sUJg6e3Ctd4wvo
F2h//V10ACNvLjCiq0O+JsFHlpjaagzOZrO6F6wnutOXCZgPjjS84N0+o3iIVrASzSjmO+h6DVhk
z+8s6KpvOtxIpxxFG/5OXF2MkKSL1jsdvKhr/glfK1gS37rnZFKHXRDfZg4uBodtddveOYiadWNw
t5E2h/ISguZWhYVZFQXtLKzbG1ToM5Ql6eQ74F6IeEoO3IibLNQ9x+owYUGrA4NbecQvVqMUo01L
4+ugO6SyfxDVhczj4fILSlIuenChsRZai4N5RJCSUTxCux/DcfHHpvzaBjufO62ixfZ1QKHp400x
V4rhAXw1SkK7naAMDrXVoYgSJyQQTodZs9m/bmiOAdp9vSVZLR4yMTpicW1vqs63/wH/GT3QXC2F
40Srl+6l4BU+TOIh/2N3JAsCu/mZW5LcBtu1yphi1ahmK+R/XsM0lb6zgj2yv8QVBmXmzteKk3Ug
04NUuKUyg7iuDrTXzCyb3Nfh9olcMQVZP+5g6K7gHtNmNk3JnWctp2CGPdALnaWB6Xik77i57Ayp
2b6t08/99TUh0RdKI40UR4S+C1MjK7HEPZhaWH4jAZ/hhTRLX45678zEZr5bRZycGTJHdsQCYM3c
rmcSodK82LhN6qWPqLKgV5pNSNx4/klNNeiVSMkeDXsZWDF+Jvbfh+W0kY/PCFOnMS0SHmUv1RBJ
/fR5jGPEQyD7Qx1ga05ZWqXJgYi8PgtbyhZIoRPMn93pU+xAzMxnUN+kj5Z+xu93YbiAmVhXDIaz
yhBZpnua+LG2z8CBdw01v8VMqpggT/nbdY3Fv1IYkbelj5Snv4uCfD/dnyWcP/LCgGxxHkLkrUTq
ynQzwPHBnqLyaaNAn1+zX6Lm42nWePmIwEXBH/3A31/jPsQu7tDj3vC+fh8hk2oi3QfTbVSLkQvj
qqP6b7LdnVCWPDN4qpcuYO85JKjsBkU3z9rK7CXZZLoU3X6iDjR+p1RjRXNZSAiOwB027/LLkGP8
STzItSpQMMlIZ2nTNkeYOal3t2ik0kolL/zf/gU3+M+XiKxBwk8/af13meLFigcMEvB+/uGeVpQ2
9YMnO6w1RQDXjls0rNJa2h01ScbAMW5rHUzanUvrA0Emz/27Z9vzy/RiDqCmJEqkhy/SdukdNPYH
vrUVa/LpurNaLYAJpQA5OPkKyB8RAn4X8ydAdcv6bdX8kWFhJgxfPsNyB4FR+fE4PMTj9hlmrkhR
Y2dIu+71z0A1VN6DUQ9UONc4FN3d+GD7Z2iSLxm0DfXOJf+dMec8DPvvAEEPvN0S5eppbhIA8nC4
g+vvT6x0QpRNPTb+ZSks3w5TQwZYA6ELFLAE/mSofG/SXnRJ140NUORxP2YRTW/Hnux7v6T1jyco
o19NiWy+uttoEPSgTNCKajJwA3M9Dxc9C27NxdDfwmDuknZ85qwGxSotY+mlH+YOMHXrds6QBI5C
Xz+s3PcLlMhMOAjQlsc7cN3js+mPrG4XuHV4pr6Q87tzH6zIr3t27DHvcw8UqZepG0yrnjRJR+2N
a1I25dhe0KGpthGd81XfLeSdgz3abXMzSCnBSQIB8XVGatwoiY32zb9ymYyok8ljheadvpCVZe7z
mJbUhR/cda07qFIJkAIBKlU0iJ5NXrlMPHhPCNkEsroN01MF+B5n14/CiiaES5R+jT9s0C1RfGzE
XAYmrEQ8YOJsKF8dIaQnYM1RgOhHqHpPITzTckAfeLCgaZ224g3SUh16IrfZpYZXUt4f4s/TLWbO
HxjvkoryhxSWELdqmLAuygIp4SEpj6Cq8epMWqEymhEfOxwaqgeVHLK4CskiAW1C8IHWwKlO5vJo
nTL9U4ilV4gvfHx+CpUouoMxfNciOKmkjRQX+3Rds6ENP8igMnPSeSPWME2KVC9k+LWkwC1FXI8q
6P0PLJLHH7gv+8z2ofvQcdOlC70LrhufEopMMdHk24dFML/MTbHenLXaYR+6N+gToEzlhcoieXWV
ZbeJq4NmzvI8O6+dvwJzuKXrp4n8aH8Lh8wbioRIBaEAyje4X9GOkjjW3LAnj/6NFW50OPeIymOF
xuzbFx/at7TdxvTm2Si8/+R/sESbKzhPUNxyQPuxkNkwVIB2IOS485ZYP+46ux82LVEH5ZnU5HXr
5HzkpBv96zCGASynBscQNromXNdHghdr/W7LnWHIywjK49CaV6OioyKhtISXohjbO6nYgyxoVZhq
2Cyre0uJ2QZRHrb8FuyCGkaTe5T3+EakEfqtquhbr6DOkBSwcM4RmkYF6W/XC80vU9vkbnIDdlgg
FIT0+U/eCVirPnMJUfLPmuffwzYA3IKKkV4jmh7OSDryHo7gLVWNKb3UDghbi+uut6w2Vs3+w0Rv
QDKPE6pcehEOhiN4hJcSwXZ1sDpoQk7T4ik7H/YDpF2oe58Gv1t/hTOv2Ey7Ssw90THl1F8L1fNC
AhajxOJ4SbTgQYGXI6G4LeBsYUKvoni4wuYyol1wBT2/wyZcfPGXwAjN5T9RMigCpw/0jwtjAFEl
5YGTfIcNdjoha21fWDNjM3OnILC4mPvXBzip7b8u3gd/ZGDywPQXW/EWqcP90X8QUmfqrmutpuJO
3qMH/H/n8khit6XwxuSO5oWgFf+qqqeHEJhoQFcNMrwMJqcdPhDCJrx/gwkSmbAFDgxDxZ+H8H+3
SbGYhQ+a/Ai4n8/XjwkX5iYlvRxZ0PMD/FAipV4UB6yqiFq9oWu+Mqi2HVQ/b0XFy4zvjFOVwdZE
UZKgftcc0OM3O1E9KFcv2ISPNAJwAvvT4cCxG7dCiS7AAyOyZZBl8aeNF7cf5rfTxrHSTtEk08ZQ
39d5U33bO8iCnVMKiZte0xeJTmkXu28TWlo4aMpyfzuyXDlVcYOHQ/grtXcETH3yjPSv3DZkRi9N
GNzB8vKzxS816vi8YgHEI9nQuaC6ump8kZ+E6PlFda7Op1nGsiBPtFhqn3bOg1Kr3DthmhwlRCLM
Gpw5XPLeqxGpmJ7jcxrLE+qiqUVbeju5j/INcDHycmNnXrzG0HB+srnn0a9lZWr1WPr1GQqAvvWx
4IFISIPeaqseCXvuNQAw1tvEhYCUFkYRbToaYw+qaBY+BIH2Kzw6U+bd9WZRjuUKKaScTKJN0gNs
LbgPUQqCc55wdgzkz2i18WgIMTh3qd57z0rgR6ra6seCXOfyHbYLlYQdHuKJap5q5H4PmWxfZnsS
hOILf2VKMBY+UjhO3KtXmiWe0ilMPE3SRAuokmNOXWvtxNoWBc6ZM8NjBkc9K+lcTfbKY/pTJYDJ
wcyi2UsKHyLXO9RhGyjb2eDU964HkoNqGEADMZKkaE2dhVX383Jhv++TsaUQnDaqilOIBhD0iLtB
v3WqiRiSnNE91Su8jX0nCo+NkdfP2VNxpHMAHA5S60azuSiOpKIIfs8G2Or5bZY5vgcwKASA5992
xQdTxHbVeo6BrIPO8QFXVMrupcEnOl6WaTGrcOA/dz7vtLAZvCCjInF55N9PeN8OYoXxziBdpyi0
utfMoK/bsKrnQa4QNr7rr4bOguTKLDx/o4744ynCa9l2zEXeKK8AThTZLuLb7kGSlybQhDodJf1y
eRJpSZmoKLUQKoGC5wgQalLImMJGtNPar5VbRwYHttska6YESsE+WkzpiiqVocwjGv1di30qUBLi
Q68LcGWZ34Dr428N8l7x2Tat3NGJoz7zcDim6e9An9uZ08M2zTZvYv4EZcE6yn7om4tYGbq9XONm
nYGOUrVUMz81N4pDrPRhpOrTLkO9y4DpNhHO1O5U/Tx58gO5Dr0x4v91/GcWHWfTOk7WjWLc0QWX
QY7LWt1Zl1cEXKl+YeCY4ukjUIpQNQVW7TeHhHi1XS7t6SFBfeb4raO86kYJDDLf2RACTu5xkEpy
3ShHrODGB1oiSdBQVyY3cwLIKEHxqe8aOfpMlsfkY+LonqPUxBMb8AZ/PEdvInvfme4NETKs4hhw
PIv3IkKHZe/WcGwsMAQ8AAoqshRypc8N1OL28tqKSJMVq/3BjnkIAaAHLu3ZFOkXKAnu2VaHOAQn
mloDiVYjP7Pj3NU5YPQHy0Zb8jtEImuTlSbp7P0OMoyDx2qwPBvoqMOm4lGaDWomk6ZyreMlO9MR
KM1vjBalEdxl8wyI1IBtKTZLCislOkHmSh1xZsZ9YzMlmXgm0PSjhoU1J9a2jhlOnCbUWNDMNwxZ
Hxn9efMyvOt4FPh3HVE9LwP961j7+HrIYsFUG+X8JBiNyRdTNxXKS9c63HXPHM9Pm719VEKmv2ap
j8WNdgVHNB5JWPH8RaHLa6t3F21YcH5PtSiWvTEqMHpQU39UyPkGU8y7M47kKXa42aAT6nRjMJ+B
zi3VR5GTbqbE4ZEA66KnLCPfyp/mPogHrIu4uubvP4YkoCDIjsdzTogSsrtBcLB66eraWbniMk+Y
R8CDoorGIn+8CgJn38KAj8WIpeHLqZWoXhvLyTuvFSYOLxDG+BNzruNsgoZw+GcUZSbRskBetKg/
PdrtGQFrWqOMb2ReW8YMC1opC5POAyckgw9HK2mqnV33ekDlcWwTrNTj0HqqCcg5o6uGc/W6mc0w
UDBSxnxPqc9SwftksOa+xWFqmIaK3vl2UdkjfjvO76VxBZThfy0g/kL0r9wvVoWu3KOYJy7u+GeB
vj1sT5TzHRpcVP7uzE05vGU4OZlnXkfhIW66idV+iY0IuSOJq2Dn1FMGo4FcHiksfXsC4COKRsYi
ViWhl4epFM+iTSl58ZpJNTLwZZaQD4UVwKHMrwCKr+4K+3iHiXKWWs6X5QCmFRCSYktyDQnNFBrE
b6EtNLmKDj8T/tlurKIjB9lw8RiLIOwC7Wsotb0eoDqAsQf+3c2IxMBcfWE2oSl8SELcwVeznfJt
7LfIX80xXVu0UFbWTMhT6hOqnJVKCR6I5Ou2ClyGIRbFzKp0aXIIQLi0DFbP8IpxesrDorP/UYZs
lmitlB0/1Ud8yNelZVDXW/fgMQlCqJYj5kTkyjY3KGvff/UbdMKXuCwLoDXOl0HofdoX5YcPOtMI
K/V+e5dV4ES2wlqIgRgLTASUQApdRYXpbwejPPV5ByEp4pS5dOeBRW7EYJ5QoIi556TpN/dhpKRX
ywQtX8gYjyKb10XbzgTENpdRY4hBxvZW143aP608N8PMetbj/FzbYjtxAsAzr1UvDwsJWwFh3q4E
/DTiRZtZxucfx62PjfO/iDz88u/LFDXdNfbboSQMLCHnjWqJ4/758vh9Qc7sdgtD6osv8NBhzNOk
M80wQO17pnYRzoilgyswRiUJs/Syc1TyPCt0EaQ3t0Pfr6mJLzG8VXB3KxZj0gupIr5oKgF00lv2
AKx1GgEdFnJQvT+wEEIUuPwEo7mf8yYXh5C6qrzCZaNxaVewMsu1VRcdskS2MMOmGGVqOewzQu64
zAnpyfZm+dR9Pxyb/pMPyKL/P1bNh+C2K31XIuuPD41YYwwxYHOYtPjnc8edHIe8NosnxJo5QjT7
U+CwSlmK8bLHk93TMhAT8+DedsF5VHOuuLThl9DCOtap9iJaf9s4nd/ZDBBwW0HF5lTNalqpSkp3
sx+82Chz83UrzwdpGYQUj8vprJsm8aNPOLJCjDxMxUlDt/Jo9VPJww6a+2QBGx+9i0I29/2rpEE6
FTiqgUoekGohVOMmPhyy7Ko1iz0cKsskE8frfwtIlK6++kFjLCB5Tduu3A0gV5AxYbnM7jWSClMV
OMoH9DDrMBxyL0hbuOhLrGTzN+H8lDfKccaaJOKHfgKeinkdCBVDjDfbF2rrkRbU8HOYxYVWxIIT
Zo2eCrxS8oGQ6juA78SVxqXMfKXsPmjvEEZ81LYx0uJapeKfmT+MnbxHqPGPY95yO4/kNWIOWHXf
PNk8Nj2VFrYJWbfqvTAj4dvt2jkCQ1j1R4rcxkiqYpq7ZsZeIVJkpqZzu5TaSD4Vd397hilP0uy3
HflcF2LJpbmF+v0KSDuVzphMRg27DyOUpNdvoZipwypgNOdQtB+8GwiSzWtuDvTh1hIpLGzfdxB2
GGUf2XuMMFNiNKuSXWbxoPvZ/EbtBBhK6WW8kZir+nDD3a6N0MHoYlETFxZqKVkAUTciO6tRbpXe
qaw/SkDY1BgAReVn1NjewvN/Z+vgftIspziqx+KUtts2n268TaJ7RK5FHFuva/SCNbgUptuIFjHS
y5gUlRAuCwfhbYFokLn6RF039w7ifeTeH9VADKc+EQmC4u8Xb7JG2baKVCPu2M7rEMnJsID+YxRM
SckgZEfgvv6PbVP7arrz9Y9wLrr0AqgUWkZo1XcXFFdciUeYRRaJR6P3VVOhV4uBnG0PDnFK+I8f
u9bG7YXO75VnmNgFvaidQG5B3ZPfI1FT/9fp1rwuAB6HV6hW6mCn4hpWtGX+QZPXS7RO3XfjCVGH
Va/LW6IaVLrocnLS7SJWMB/YRivhH0eJRDiFmQdi4fDfkyjgZ2pzre962k4aCPykJf0dzTaCRK6C
22Tg9FZBr4clEqWdjV5wM8wcSkUbveIjXo/Uu5uLqhSGbuxAzTtHD4HPaEEJrTCLoIbLFmNiWTrO
zhAfVq8hRFro2bj7FqY+LrFXRRopKSUq4Qx45iRVJmBHiJk9iItEPJE6mJXavhLphTYiyPniEuWa
+S0d0Ml5PQuzOnbKhwkPf2exJdwmZmlSIxwMSCa/DLZ0igbNLMXzSeZxE+Qdr2OR/YriRHtaQOIR
XMoFwth+5rDdJLccsY8ESbGtLL5ppdAJGTwb3Xy/49CT+8xX5oWjN2T6Nc3YVvFmsRIZX8JKXj96
qaCRBOcRhY3YQG0YdEaXgDYfqsCxAeYmDXfd5EJWmgc0b6uYwim9iBbZHXHLbmEpReaG1WIZqbTG
Oky2j5NG0KB+/QRdDlS+RX1NOb+8y9vNvO32pVlp8kPqVCTbTCCisBLciqqrMuJZtPU2ugYJJ09j
91elS+fzC6peGSuZwxHSetTsVVy7Lz5Hnv0cy2pW3QUbSy/Tm8nVF6lGOsgbYNmCoq0HijN7z9tq
5cI4Yi5pd3Z60A15Cbbsinu1ppNcOC4fye/FOyFfKoMXC41Oo8yiICfrBzi/L+c0z0xMUtMvTT+W
zc3yHhKTfNOENEw7XHPcp/LkfDzZiwKA9gyXurlW0rqlSjPtoDiO8Krw02b3VymknPpNWikVKDnw
24R7mYZ9Lf3Gc1fZkdvIXWMKKeJTRM+/3AzYZ0iqxcmvj4z3Muza9C/G0PdRlwNhsOb7tiGJqIaQ
aGHSitvOfoharYyCJ9fDR8doihUvf3DLd3S7EVbEzIMYop1AHo8oP6foNPgBw2m99NH6EdxGGmmr
nPKIvEKkEDya7LOwrsmO315n6LUIDMNU5yo0/vQmsPxgpuxyl5Pas8bbjLHEo1yuXdA3N6m9VlM/
Aash258wJHQ7MAFcs2r8j94NmsIAFOFJLpibrwO5eQRdHxb25RrdGbMXvSca2fYAWrb5qxTUB76o
EgTAtJMhJjnfp3zYmlBzbQQeIUJZIO586GxZuGGOP2OEvrh//pevEtbf4eajWt5BSSJbKMsJcI/z
BK37RPL7lz974Cu9eaLfrNshRQb7EN3GNKg2x+JnwpS+G/UxzFmm+4BfXKe8F1mdYbkHT2aRFkm9
XJ8VnWdgxCVfn3vFpQENKhjf5TItOU20tmeBI39A//JL8I0spxSMGo0YYoZ0DJf9tS45RlfUsibf
G5oIQvn7+fm2zENMAQCmbyLBi6mtH7wxC7OuWKm4hUl77omx0bKVaaEuRejSt50Vfs9yyRLqutmz
3JfXQaTvKab3BLSbu+W0D8H6NraXVZa9AYyXVO54woWKwaIeVDJBRhonCjxcg4XurBgcQ9A20vab
LOgv4EhovHzJjXmQQmTPBY2a9D8QNhefJS2E/bsu8UVQRqiEK3A84F/LZv+9iefeM6TqglEaFXmT
+udXAtVKukdjmpKmvkXQroCGIN1n3hJUO/cJrnkcplF9owV+kXcw/Y83OvDYArUqBv1W4CJ5CnNn
iqZLPatw0C4SELY+S7xMIHpmZZ2sMWrVJlrkaEDL+RDGaZhnxELKv6NkflFnwlptUzG3dpOmqwtJ
s2vxQiNvopzMFZwpTeJAOhcLPMmMQVzpmui7xhdoBTUrJtmoPU6BCnw0JiEnE4hz9fHEuKHZVQkg
dAUvm7rY1xOcN3XiexNhSpYl/oI4hoPEWvUsyItBCNG2Y1L46U0k335p8IE4H9CEw6/8nZiNN2Jl
i86K14g7S/Xw9qMWFKYuF4e3Y1w839pR/Pwa/H4l3Zf/YZXmX2w7+xsJgvY+CnvR69erXfK9RXU5
w4korrqFRnpLs6WwXGBfH7J41deTwOrAiFWGcjFvkaoIBaVA9Ku7Y1taKcJ7HpgFfCiphJbmjZe8
V5mQfiM8+1pe4K04CrQUvtl5MOnjGaN0Acnn2crP5K4isP0vS/qGguAEv4FVpVZpX2cmuCwKoLSr
syF/DjjeUlqdb/Zj5YRARqioztHCK0MI6/FI0ugHDuWtJMsMWrDFDvo40MHhW27I/eOnkt7gSA4z
9NHRwi5xWI7SHNJ5//Hyju7D3unCKz/xW1lORH8WBHOTenRxOYEt41TUoOU6U4Kis52lCIcOsw6x
t9ky8FB9rGinJUEetLBoHQ0IcdCu12YZ/3FDldaZfRzSJUyAPSyVlfIgeVDfnfKu9VkE19y0kCC4
/XIQOLqdeBimEUkVGV9lXeuGgJswdzJAWnz4dj4K5tIGClNPChLnmLOHC4J5wzstuJXzMONIE7XG
G6cOgKgeMFsUNbEtmlkOM0KNDUwjyP3QOf8xkhP1vw+9mTosHV4KV3+8HpxpbsQWOGrAeVZ7prEI
Zqvtk8ZwLZB/wRXTGVnf075G46y1eKeZmNQ0DBXf3Z05kd4yFQhe22In5Xr3Dr/ebOj6TR8IwJ2z
vAJDaBPX7zyoUqEOvqd2hp946Ptp1hktC80/x/EPUEFaT4IsOVGHnzVLAAWjFWJ4G8ZMO4zMUq4k
SHgbxvlnm8HAV11Kf+5QjfyHCs2IBmMpaWRC/n6q7IhFy1vvjOvThbro6bBdOCl/0lFvfEodZVXM
Wed0Zrk0CX9aUTiO1BmjxRSJnSkjOgl/16l73YTET3D9tkpHIaZHWyfgf7r1G8Z/AtF5mTK3eJGo
T1k6RuvUORBjtBS+witFMbmnZxa6qJIA4gCHXXnN+vCnFcTzS0R25lYymW6UipWxGfFA9+XE1/OX
ggMLfDkppKo50CvaYYKDizyC+JidVjs/ymb6w74G5/d0sxn6+efw04xWnRCMZriasxvz+2xU08bJ
8y1mh17QElukoGGeVkAF9HiizqrINpsvZZ8xkr4/qMEupsJTppPeuoo5Rl978sBWmpCF9rmEoS9F
c4mSs/sJ0BQSdJnfIjeklIKcnLv6/U02AHOO5wAhR03hSLMnWPnUd+S/z6b8XcTn7fUJ2ymuE0p9
aCwPN64YqlPIXD+TETXNE40vMwRjcT+0/AbHUyY59HqiDl9Ou2+vpHo5QdIWivLiHcJ2zqnXUP0k
/TU8EoSUjkJEAeVebav1uVhetje7EzU4mWFEo68oaNy6XC6OeNDLox05HUvcHr+pE2QPdA07YeVy
JT1UN0/7izkFqHMciR3j9D6fv/6/eVBnMYJNKDwgZHqGyYhS/fn+phMYZYjpqrK4yNdZ9kkTDrW0
OaPU1O7TLGUAKT3jVbimxQDCunWh0+oNghPysOvDYjrSJRMpV2fieAOVKqG5MWDwH6ryYpzC+wUR
tr3/TNstZpnboPBmt48gGPS2cdGD0g8l1jQJfRpQ82erVMEvjMZvWOTrXH2DryYH3dwMO8zHElN0
lMtei4JjxVEyVSasuq2BzJboBgquOe+2WBit5QTywObb3o2FEd+jKdrt2EAKTh9i+yL7oaw8AsS7
7edF72PTwDF9d7uo1VNPA5SVkWAyOabVTTQKtR2QkjnqJ4LT3PELt+m/nRHaVaE39TBujY9vjR6v
n6simuIcIxg1RvnUoO7xIhqPeiC3vJ/OZmEs2VI5usPBrq3+Z89ZrONF7ZL+4rIXof4PynvtYIew
GWPiviMY2C6XrOcA0A+qfH5rG0x3j63TDGF2ikLo3wAS0yMgpEeoI79PTrV0VhC8KSINMwe0JvX5
IEMNfqRRgs9WMvMcgHLlLXJPe/75E0VgY83QjCabeUeI4dTKFei8XBlFQN1Q86d4DxwKAX/tVUVb
1NeIAvx/DoDIo3qrsNH0M7FUlpOEaFtL+JKMjbSbEFo1vqXawc9V+3OkrFFa/HSzj/w6ZGLFqfKw
NTQHNfJYhoaugsMrKyBywPtkXPb+z7mXMjBIhI9KcN3li79p1o1vxoskjgvx9oo/00a3kmHxRtK0
AwIdcm+iEp090rjMbnZdP/CszVIS8svbOx/NNIv2wb8pVvVpWVpt4+2r2tx2hjRErs7OLB7WbrYV
jIcJvorTTpcsP55Wownlcols5NuvpnZ2ajXq4PTbNEFmUg/uq2GSV3yDKJxf/bo2xsK3LS0LW+W2
kMAMsQ4q9/j0WFJPshwrshADvhx7JRyg9zx1NO5CFvGgNaKnA8ukKHpeMz626Rux73ly/74/n27x
Wx/Ehab09cer5ksr5nDk5VnJNrWoQI1KwzMDYCjXPMotj4wjiepEZitwpWHXdn6r6YwaG2/qcHMQ
m/2O8Xq8yiWPO3zGxwKK/422kVI8hs2cX4J8Wra2cUS0Rq2bHfrQPSWXP78f0Eh1LrohK+weBCY5
5dpRIDG8k8oOxO72HkqDlu90wTcXOUcYl9evjeqNNh4HqQluZyOlF0sC5i5J050VfeCylt4hTjGr
butib7iP0193JZr+cGyF5ut7Ov63Jx27Ust3PmzW0iTTvn9sWTzcE6IdevFW3IPRMUj5Gp6eZJBg
v7PoLuPf/jmq+BRkcFahAK+HvAHQ7sBHF9IpEe1LtwvriPaOg//NqrYOGX5zsTfDPaSRhHF86kcc
ZuMSFxpDRPM6omzyDA+D9cJMzwJhMInLmjQoTmyjdV9LwohOUM1Bx6BriZn77PFORzlth2WQgBNy
rA+MwHmUWw4G+Sdn1SuVk60g2AXXeF0jWM248OouQ0z2pRJ9itBEsVgHAYB0dPj2pj/S3S+Qja1P
g9SIJ6DT85HmedXkllIkaEKys6bsVGfZ4fGkbqcdTdyaXAwQnHx1GXAxsIrpOjJe688XBFGUYS84
+iJsrysRBNXaXvvWnE+cGXO+U4qTGGL9YSH4keBQH3236TKl1HZ+WrO8RPWxe9A6N1xgg+aRm2q7
1JnJjqrE9jh8i0cVzcctWYWiEdSy1bM90SYOp0XZA/I6yEkL36oH7dVl0d0iwYzASdMvJig+2pwn
yLPDePNzblmbafh6sU893E+iinLeRucXBYYUsmn1nWadDJHsIdSBzYH45n9SMFHbBgHkbPkVLaHY
d58gscT6QpFaOZR885bnZwiYTv0qKJbbIpopYQ7hvwYt3DstuM/oOlla75kqwAjtp+WOYYS6Zv9e
okdI5ewLLGL3t4zcXIE6vgxuTE0U9GW0wF4KMMkrAwB+0l9e4CnWM/uAopNrGyC6dyrSf/vIYRhQ
C5Rr7fr6cMtgyb49yRcVA87aziZvQAGBwQ75YaE07eN0qNF5WmieShWvnvNiRnAfwTi29vkVjZ2p
udtJyY5UGOBfGuNYr8BlaIA7N7wXHCLo0iAXClPC8Vekpz4m9SK7sJQZ2DBUcuU9fs0JQCHXHBr0
9mwW4nMaIidPgxy+C7UbzNyX0YNx1KXcrDY/STuJxGIii13bMsvEtJWPTIJDyrwdZ8+An/3af/QD
mMFGIfvAQgRVjuqqb4EC81lmpwSlJvJxGGngr8H0iTpA4poK7AZ5dcXZsiSZCDxsQsFlXsqBvOyC
QDQl8kfb9q0+hcC/VEs/Getd4TH0hNM7ElbEh+lKtkDWorecyhGNWOloXoykAmOUv/9CFPgfD1mY
4itlsKP/M+FLMyD8zkDUk97UhpHLpDwXb+16IBAFlfaO/ScoHUVMlW2rulFCgPOVqrn3fpZ7eOD9
zoRcVOL1YIYJgVnGM0KkaTNiGQ3pUrDH5BaMq0Vn2EYXrpQcXPXDxsau0RP6+YQtkFl3hyreNT6r
TTFWiJ2l4dK/mDHKlcvxul6kwHKEpVmcdbXYPGAj9c//pWT4BAMvuYhg20T0M1Xar62ZFXSTANzb
z1z7AAN9iy1OIh1DPxV1gkAvDKO+byakjIQ6lFKGi6gyhDf/JEn0R97K1HVib/JFeykfMQFxDUmT
HhDqlDThq9UzzfdK5iXmKJWpDeRAhdircp+AWllxwu0+Q1vrnCHtdar+UUG6784hGJAP7K1mhbaN
w8CO3JyLQfNscAIK1hIYKPraPLZZ5m1gsWvea8GQDxjWR8xlOlA8nSFyLQwVGzHGX9EghaRex5c0
eY7Ss+SpFK6GhkABG4RlehxHaoHngxQ6Ie12dTHKKgYdnm4My7W79cwk+0zG93N1Cac1nb5OT/EB
49O4+qaf4x+X9bKYSHkU+NSqqmgTDmN8+MqQZqekpn3h/XAqAednOc2ByF62Fvw2IHeYsKcJtwnw
Yn/GZI5TFgAtfvFOaYHTXJS/Lx1PjxA8FwsO3rkrMHQaTIAqiM8OoC/Rmo3rNnKtfYi5kTn3UEX9
281d+M7uu6sYO+vnikiipV/Y2pv+giJ16v4F/9yHD7GgfBgsKccnKfax5W7spNdrwduMlt8ZKpSY
qrjuu7QuFD3+YCVhXG1yzNf2xF2ZEf3oVlQWNyvcpOLS+/8l4NA5rRzyFfVSyVoULKNt7t5n967E
XNVOxDsknozSH8GVyQMzBRvDnjT5Nkf6XIdthJ9r/0nBInym1gsOP1scEFeHxFn3N+PY9rLcc9+K
3HO47AHj3HtjhJyGRH00GwNDtiuP3N9GYyIf71Fl0chtiT4wKExdMR/pSTX4XhfuE8PqUOAycI4J
CdB+ClTFz+2BKVIkaSLsBtfniW8itQ/H6633LE5BS116xjElKgfhK+dtHfwuescXN4mso1YtWtGo
iEqFZJI0YBYulquIfo5NrG/e62/To9mpN/9WgdH+oMkZ4Ov+MZmKwo/TExJs2HTj84kx3WrMmhCT
jiQu1tNUc8aJ2tgDNufptjN44lexDPWFw+7m29Ee9mXICv7wSwnb6rlaN5F8fR7h8F18lEOrO4sZ
NUfaPoLI7MeFHHPJpRfM+cp/jvFn3lQ95KoV49t7JHr1IsThWZZRGWjBmyhGKEOAeuKiVKNcK27a
lFmGdo6gxTyAoR3zKM97sJe3xbIvpCdhK2mGJFRNLmbehO9J9R4k0sg+w64PokPUB4qE+Dd2SmYP
qtuSGCZq2wuVg0fKcCQ4duQYzDQUmoNGHr7iG14tpSZA9w37Cf/WGEEzVXqwYO7fD2ciytc1oVtJ
9tNzvrmrGPzWTcnTbgAjHSYjqaVO/h/OChw4bEr3wp56URmzKq+7PTT5+uJ2aX0c4DauXL7mK8cS
dQBgnrxKS6kvD8eyjpvKioy4JXk2KhDPbxl5d/gPNaaYO/3DienvyXYmbfQzZTW7O+kRe4Yv6ikG
gKv9D4EXUw+NHRCLRRDJQvsCqdipS6CGzGGYwEQawjeDEqGnQT6bg/NTmf7o1rKJ3fly0EsV+StE
ZgYOUXtb3M0DEGG5OczDtEeJw5H6Q3CG/PkBLQYuOkS/Qrt0NEUqUTYneHBuMMN7od+JfEKgSd+O
+NcA1ssowsrhWkkNrABm0JcZ4xpCkxaBoeHWwI8NE55NzgsqsM3a5qJbb7p+hq/hBkiWFdyZyRNY
j1jxSdLGGqvvJubhEbLbwTFn4N4+8eubBt05dSc83aRRQvdEb9c/Nc6eVVMU1i3e4buWjxlMdea6
TBLtfZLcCx7zj0xY+2o+GZs17efPPkfH8KiZIJX4issZ3dm8dmAXkreTdZkryAJ+Qkqta1m0ji9X
7flGc9Soy0nknoE3QkzISVxfdbSAXH9jrUN3u1rc2c9joR1YJnQ7TqJtiMiMpyyN3rUGph69zosu
4Ivw5EliiUl+jZn2gxzZC+FUFMuMJS1wxyvihEarzUrhjSjLf8aExF+ArcAndAEW5wuqSJBlHfvZ
2yiPEr6Jtk0Vrg7ccwOKPmdm2oDX2WR3WcI7TMnQS/0NqxPNvLjzNrtpROKy6zwyQzTXDB4G+562
th/b1hO388dEkHhR4Squ2b6qoL3koHPXNg+anDlFrOCrjodgE7wUiTF+74W+ZVHhsy4dGzdOUTuG
GPEuvMH3s+MMDw1a6JJvm1AjBM8Zfqnb8atEMn6zjtLI7/PZtgjGBSaHfqbQQCeSDvUjFwW8dFN6
fOpXeZRhWobvYi7RdOe6Z3Agq2OwzktZ5SxIAqDzGho4R8zZ/KVrZ8asA5fGrnWzmcDwc2Igdvpx
xQk54EcoRqZ2a6Sm/eDxF3PwomN1VldhyU1ZLziukNniDXdLH6VVQ7Uy5yj5P2PHZvzhkTMcoPRM
7nTIViN0QOgfKyNqJy6V8MFv9HGYJx5FvP9wS+0cdg294r+1DzKvSqnylZTuOUGugrL1Wt+SEp8T
o4hzLPctCO02/S576doW/AffTzdZcNCwPbkz1QhGEHnOdpAQI2N3oDTMMt17SGdbcofnLQ3LLaNC
d25yVWMS86tDQpjpZJZoMlEC2FW1y3wAWhTV8V/fpzv8bSfSdb/JKWm1fuKYgSaMcCA8wIvwJOdz
7kiZEv1Xb9mhr2idBq+3xamRHDLVbuoCK9Sj5Z0mOPd/pUDj2VEzLBRMwSCy3+kLhiwcO1eCEv1d
N8xGRc11OsiBSFWCBeoJbxgsIaqZfC7bjwI/BTr+vSopiR3bFrgVD0fJxAk5cnqjY7lx4pDU9BNq
RdB0zysT5sWMvPBHumHHqP/2lTPhh4p5DjwO1I5UXnXVuqGljSSkaWZinwvo4x/UIV6rcsG9XV2u
FbQ8XQeDmEhwbAoiUri7PBOvzebCFBxAMrXXk91xP57KhvRjuL0nqZ5OjNuvLg/03INjDEusTEM3
6hu9zVfqUZ4q5gXCfyWzpyCi66iahj1PLw6NvvEFIAJMpvpOoHkwyAgXY/W7Mx5k1c6w6gN8exmT
BfOkQA2qNqJcbcbY5QitfrDomlROxKQzffxYdOPW7SzQkE8L5WRGAIhMssIlqmgd4CmYKHCR5Jnb
C5aE0NipHZ2adt+jehlTDj5OTg7t3KdNKpkeO6NpYvQmYhaYiXY+LXOf1vyu4poAGYHSWCIupAqc
yf5gx4sWXiyfBBo0riCG/cOWwvlKSelt9sWCAlggACGGj/oWutUIdm0HVPn5gXviqmp+I097goEd
UbIaDCzWH5NB7QO4bq68MUEti5URlbmEVUsPILE6lq9RXITUOFwm0ldlmWUD0iiG6+TFHui+7Ow1
UEbRBu6eHh0dH69gG9o7+0flN6aVi7jHyj5mPZcxbChyu6alHz0zgG0r2CraCZkglvnX3Fw5azJC
fKz70Kxqw3Taj5jSdsUAb6U9A9lApHySoehOFmkmRTcu1glHl48/isgKhCAA1LYiBYhVIH4/5V2h
Bmhz91qunWv0Kqnu+yPozGQXrG60/I7auTDJVa9p5HmFyWt85JtxuR7GHE6amgTk12FbeAX0J+Zt
kVLr8gBxXTxnVFWRV3MTW9t/1++S+e6onU6+36rrCMsmMXQtTusWalGIZYxnU3U2l6jQmQk9NtLj
i9Qa58JeNuxPf5FfxmO2OAHdKKNCHTieOW7B7UmEeYd6SwqTf76JjuUSF33SBGTzygqHoXeXfyu5
Ij05bWosPKPy1G/Vw7VF8W1+/ztQ+H1cJ/QSk2CTjrijmiUewcYUSwDx97a3tcN6UUhyDU8Ob1WU
Op2NmpeztAOogeVjHkhoaSZgua8XkPAVl26aK3HJP1iAJux1BC8krTOgDg4WErbhLOHIxhnGm2Jd
+nJdqBJNS/+WbSpcyuFYosLtx3Bd+R+SNTz99SUBWGFGFMylgCEO5ERn/nBdboiV0grQcE1flj0T
KCDjiUSSpKuWwj3TOnWBM+iGkukcHHEM863oF3pRh58l0R0Gqfdv+KP49Mks+2eCyKMUEoUoQXiP
oUO4rpz9GwPh/w54qyaJ7Y3wCEyDpGaAhSF+uQQRVoWtPbz/QMm7kfA8ReKJVV2ntGSVRBmw8wgQ
Ju2XhsEdWqg8KP8S+/mUPVxRZDg+LeRNZYK+AyjZ8PIBTZpleAhmdZH+l6+qvSHQa6k/N/ZE1VuW
EVyZb2DGi0nLIl9/31EeDMAf8pmBubeW+kNqIES9ULwLxaDruXd+q2IgldS6+ade6vmNQs5Bldt6
ZxYhx8greKMXfVCKHFst8JRZtazJpLdT+Zbv3OjQUVLlhsa1eGxJf6mHylN3ori5jeJAezRyCanc
VV5wv3Xh1eyfwJj7o5M3T6NvpzYE2EyVuDNUv0DBsq3Axfpji/z9tFKSRS1bz7Mt2tAotHKyq6Pl
VIYIfL7+zZ1k/ZYIt3gWWBvFtkmMQEMKY7gzQ5pH9qf1/54+BYXmhwEq21hgNxmtliUgoSfM5FJa
enlALTX0+K7ekJEHLZogVoJODNJ2PwoOnn20fyeQPTGB9hqYKq+JgxpRhpg+Vap2pZFa0am7HsRR
+rbbmx1j0PLPGUzbkia2/kfbtz2bAxddun6dI73igYcAlBt5HwmcSftV6ZTiokECLszFxwRdofFA
C2a1Nr2sKrHKIBs7CfFhwE6WNmLl4WRF4BoS0wZVDkg/eBei+mYeokRADvTAPkjKJWzu/VsgOef7
JXFC14zZwq5DlyYxpIsJIyh7JznkEgE3PVP9vhzFucHH0z8K4V/zbYb2XOTn//jnyPvF70GXQYwZ
crG5VIQjKf0lKRuHYgMZeQDWSnr9oHBeV2cbjlE3c9NrVjkpPSxCOVUYGg3OC/l/T7oJqjolHaaL
tBIxrabwH/A2N0CbALj9DIM51QnMlmrezAx/cwDYzBcgsH+YG8eJUZk740/7ZFm2h3biAZEbCPj0
Spb+U6U+vFPCnDdml7g5dkS/SSrn0Q0HwuNcQI9m91Vn2tG18MfPMXz3axcRZkpzzfvyXJEjaOt/
ARdc76pKuIvj6rc0AWL4FQ4C7YUzuoOgMDPJ8sjZHqkKB051pCDysuDgRXFnsFYRB6tcHPHRAcfq
wqZ097+/GwOJRfkdRSgR1R2xwaMU+Eu5D/TzLLIu5pnooDTA55+nYwo8wrfcws38km0ppYn6CbR9
muqnMTLN2HIt00RJYx8Wv/YF5EyfFazToNNDIUQ+G7dQ9kehk7aGFKCytyejZg4o1a2UasYmUFHr
eNcaO5hzJh+CESoB6MNDt+6TxrviAwaSN50ae71ecChUv0gYTXYd/WI0znu8OQs+ZmzB5fC5rzQs
an0sHtmQ19SFbISXoS3JgxKF+yniDFelqC8801StgIMiXqiU7OgnpxhsNB0RG65gPH4cwCqXe2Db
JpQ/7TmFqIwrlUQYvGKi77cOjyJiFVpRTtxDOcRjL5YqcwpjPArZNSn0OfOdJTea+0BA7g29kC3t
OKLpX12TkWS39yBchbPmosWBLJkH4ErwjtcsilvxwSiMhp1V0aobEut3vDy9wAN/xxJDEmCO+YJw
yI/d2iUzVNFh1eZB6WrdA/IfEPdyptYj6FPd+CnKFdZ9hOHbXIC25mMcjB0vaqmpBDMLdZwJUB6Y
DUIjeXIFw877fUYuJMcuJFOc5xaiM4s0fwgaTAuIs0Ao3Axe5EY4x+Y1VXPL4Si2l8CUK+oYuqo4
1J0JI8jW4rAfbyj1fIbY8B4rpuCgRqlXhggCfayrS5wpoSjHXW8SVZShecsxu0jKcSu8qPtzBtTg
IuEiohOGV/Gqq+n7QuIyQyB7S6sf5s7MxqwDuzIqnhEA87dgaiXwMgS4g7yUpAyYF1+sTAxmabq8
dJss+peBy9/hBVQ9xOapEiOPsi0u7YcUkHOrhRc21Z6RHodKAyo0nJ8i+EJRx4DrabZ6L13b5OVj
J3mehtHpPhOxEZnVg1IU8rHntEI1wYw6ThCa/01p7t3hpFYXsJ78KWHWw+YQ7ZqZ21dx4bnc/oZk
ghNy045zqcobn0VfpWsLXJsbR8pwsECIhja4IAUFLZFEjp09+vLtunDGeTwT43lyd2IDYbBPoYNN
tLq9pB9V1DcQwDmlKfDoYju1ddhW1qS9GOnMILU174BFYK1/iqjCtUFvNksdLtxxy4eloWU/cHS2
Xph1PuX+cD4AZSQNGj5fcESb19ZEqBJa6DR3dofbAEP+ns3KrOCvZ/3pPCwEYgarUZ/Wmqyn6UyH
3uBYufJgP7KnMhlqehVIeys4Iuv1zM+UA8jDLCsYnAx2zoOksKODgYGZKSiWMBrt4Tb9njjMO8GR
WZ40pVMi85onmacTm0gGg9hS01DhJu1hqcnziHkc1Pbz9BU1sKyO/+eG0wxae0ztpGLcEKWe6fz2
3QuhQ9xewR6xEr7tJpqdvsYXZPN+zH0ks4UKOqVGmxvrTgPILuJ7iqAl/Gm/PW/Z/afXLu4BHwRI
+NZqvTzVQYv8nwUgDjmMon5kZfTNH48e39luFNmKYQMsmCogDxsIWqLYRirafR+9bZoAw5pcjFit
uCGY5gGwjVjVPjHAQN7aHqcJwmRn9aPWURUN48l/meb+xDuvjdOJ4guhx8XCcG9QS5e28ZqxsJHS
YSN5eA8qcaSW0vN8OzWgu+WRJZsUp10nWX8vefcvgFKGNR0zjqmZPhl7KO0Ugqc3j/Tu6Ih6FWsx
zh+uQqADZUUBPj40DmNC2IO/bAiVj8BAEa2Cuiu30bQmgDDv1iof3VTcdKp6dW6RWmoKr2ZIWkGI
fYFbcU1qf900XOY3/A3/FpYraJLpICUihmXLAe3mkEwENIHRRKrxjgX55e+++H98eTWG9W515k5e
xiXCRNDc9GBhCMFzl9kRzepJGHSUpfh107K3/V0/FMuDSW5PZQ98gvUu7UuRilDqZ4hrydvK/Y3y
MRNpGivjbZDZ/wY2QXzJTyuxSW2pNwkxxQ9zIEjJ+Wo0RFUTpFX1bynESwAQlq1AOEq3uY6ZFq18
sUYBXdeWNpisjUsACel2TK8htBmOnLylh0YTdo+v2kgEt+wTduXuYf7IKqZfCYBGbHkOruma5UR5
8pkVtPp2nzZFNGOjtjPN9I6J9afWxsb10+3f1IuSa0Ajkwpr7QVGjwuy23hJGtTvJPjMUifCCVJy
xe41wPjaRZeHJoPccbde3/T8hDXkIyf3Z6uosm6Jd7Sw55lGo16FdtTD5Ek1GxAZ42Bjb5zBcvKs
mUYKrA8daWWxZ9OzOGA8EbuH8yaAHqx5yMal44+cCdb2vPTn/D6TlvuEWZ426cLPRs20q6zBng0U
AW5Ioj/aTfsv8DkKa+7C/buwe8jL59PZEnTTWQ08x3HzwTzCDMnD+LNHXO0QopbSeKTEBi4aRAQp
pGrak0regMDJ/eGfpCIk4z1jZqNlRzMEhv7UmXSwrxuiLMUz1fqDdf3Ut00hVojdu5GR5f5I3N90
VR9oHzb3ThRdmdx4Df7C0kMtRwcUhkUAwt5hahaaM9yfaLKIQkLbdKRl0WVQ31sHqZDkBhoWK1vm
wiR58NYr6CAkuTSoFHlDBql9kyv/RqfqV7yQFMf3OMuQHwYlZdAs2Vm5rpp2IKRGx9H9n3F0Txgn
A+X38ZoQWBlHakKz+DOzpV3EYojPHyK6sJVVoo19iGEfdunLr56q60EFWUf2puXOyk3kaDW6zfjx
kqBZNwaUhPlND2fAelIIsjUmW5BHCgGDiSk+GonnpnjmIHxCI3Er5zX+J0DyvniwgdAu3AGduNYJ
cfKdgqeY2+croOUA8GKoj1dE+pbFkBWvTg7fmnkR0mXPF1D+Eimk0gMHantKy8a7ml7eCLtxjsCS
sn4FePPtFo2bqQGQ+YYGj491KW88WyKqCcuqrbMXY5ZabLZrWhBkybMKgYI3K40kfH+yt35Kp92P
s8KzPE2R5vK3BVEE2w2biYTWqY+qCqMXwg33CQgbaPtLaiaKjXKuKu2FwIvcshMkEw8VjAImkm2F
JvLQdAqfl5ZkxzhLXm7zQ4YJERpt11KxOS36o3KUXMxhGN1a0DrK6S92k7+6EoVgzhWtIK/5AzBz
98vVg7DaWA7mnHV3AKjVlwiv232Tj/71Clcb8nCA931Bly4e6usk5mWqYp7j+gPNgFUddvMG5RaX
xZrIackwEN5sRbcAAC8u1Cw7RLBj2GK7u3cLx6CU0bv1uagW+SQRA2oXXiYTOgf0WJ62LZvUSNBp
LbaNJsnHfPhvbZ4qV70G3uDO6yMbwwSCqyarKQBUQpJsX00tmRKWZms/I9o35iw+RLvnJXv+2/wY
cTt+DfVm8foIgQ3KcShb3wPz4IPhDXeE4lDbobs73C+nBaiGvW1SaEDrR1RS6q8iE1KDlnDVAWfy
1WW1syEQepfFflEX5nNu5ZAvNGa2JkfIeXUjBB8JusD7hzT/nD3rw+HIrPEUAITVP2CFgiA1N3S+
qIgFr52bvMbEmGU4dQjCeytDK4fSGs/xoii02bKZMhzyTdvupQpDyvPV53WTK+T8eZRgOh9cneFe
EV02XlD3lD3R2jjvdN5QFfb9maa6VsTu2yjkBNdnRZXJ34pUF0HFJ57KnueiHwBXAUgeTDWj7q9c
muBtua6if+4x/7M2P2eThMcuah/nSIWW+sqIVlVOVd9vF6Od3dTMgprIjW+oA3Evykzuu/80huid
Bv0lHKBOLctDBMIMf4/H30KlxWzsasFElLewzNBA7B64iy1CkijDNbiZXDByqO7uqRyESH1L52R+
m8gHeQgN7LLpBMda5sPoTu28wLF7iYSrNKixqiletq3wXUNnG8rc6xWnyDoJdsmLsjRldSAu7Jnv
8KaPYk1F4jPmk+GwPTZ9PZIvzwOqL7KmR9pnjCxSVTxceaVTQHgCSRN8hlhJs+MAnQptegxFK44m
KWyVav543REhPfukB5GdMFWxMo2CssEYdL1Ga/HUbHWvOpkkJa5q/DosUpjZC+C1FAiD988/5e5+
aIznHQPvvUxb1U92PLaDaOtNsl4e2AIaibXR+PNtruc8ROYyZRnFI2LN3DXiOlCB4hFuE+N3ceCi
77OOY6FJIiwiEoyh83b9sOOxKZPTLQaZ08+X9m6PKe6Yy1snNSWHGI6nGIbVE6308mkQtN4uVc5V
Kq6+Bjt9ltkdvyKtVVPrzLHVoJWbLWq4Mg9ZyibCVz226DEXNLNDyIEoOdmjeq9BASImC1STz/WH
gaCinHJUoUWJR413B82JAuo1S9smuELl5QLm1V4w461GzyRumatFeN4FnOozr3IC+L/wLnoWrOpH
283jogzNTsBXDfdXjyVUFaNtp4g+BwriBCkuOa/7SiaFA4M2YyoDanwST2AExgRr8bCobGKRWHx4
FlFcsQ63c/NraRQeOCX4wxbfZom7/bc7JCBWET2wXO6pWKXdoPAuxttSCQ5B84vZohSW1r4tkWGa
YECny0w+HutAki+zt8/7SdybdnQ1UO/PNGq2OqIQsWv2uprbHw8OB24BlVq60c5Y255t+9GXb4qy
E9pJjWuZdRfru1mtF9esBYiCId4BlrTgO8AdWt/MQuzi4ns/6IzQaWiUcoNKPEtj2VJ0er8V/qs1
8j6jlE6HgVVtWQgkZ6OMY0txRBmOmRJ/4jXtW1Fa3r3DZ5TFFT+fS5k0ccC0z9JzkRvL18+ynAGW
7CRtxNETqG12YLrAi55FctXDrF/1TTHYP00uq6wLYqVeiM/ZNnc0/dhCZvwf4pzmnvXsjoQllfwr
pMQEgs5DmeVrS8q/BkHXe9HkJuUyBc6vrCIavMH+wcgwJzE+0RanIPgZTy7haPfK1jSwNod1uSqt
+m18+vfbV2TT0wyptK1bwt9YWcqNSILLVpIxDej8l2UDiJQOZFG2eCoG2PfNyucaxJUVoWOO9san
HqkXDxdNelE7TEHyEP0ExuStH//B/eKx+o+HsgL1gmC3TAXGyeB67ZL7qs9BkaSQwDyV65wZ3nzu
ymcbN74EIVr47NmjCGy1C4cht2yv0v/VT2P4Jgm9r4rW6o1vuVoXDB+0JW6HbbjHRLywGN0f67ll
MbQCxSVzts2du2G5Qs1rDdtmsafVR70u760Sf14UAscqnwzEUPpxlw5XmXmJdLER74hubj0LK3sB
z6wjEemnfaOEXXLPgyTIU01tJB58My5Q5CgMKxWILuI+Uyb0+c9623ndQ09+RkTJuDVvK3jccvzd
1t3yNuLUM9S52DeaivyKnhy9tuKa6UPVg2YOeQaHkKLvSt9ef6KNHWgHUFaWh74OvB7A7k7D6KHO
qpmEGvkmQMAgpEVHDUiioVgXx5C4imIwE1LUuxj73gYJqWLlNeyJC9+1l9dZ6/9rd7DyxvV5Hh8I
Qix0djTvKb7zytercYDr6bBmpOlJMX0R5RN+vwmmTMy0vLMsIUwO47Xg8jiUzsveRVsUMWDpyZc/
UXVKtJbQhPAmDBDdZau808ROtLh7SsaWNOU0YpIdaM8x8+NQUBX1naAidPAS6ZDb+T7MdEenvJ7e
H0paobj54Is/O9tWjuUWShtOURrAcYJTaAxvewGLMZ4352k2qIlWTmPTGNAOcsAfgbnFiOcW0hgn
y0QToZ0Qp7WB/3/UgvA3hEAFAzfiCA410hZvEogLDLlh5emGvfuoCaTzuDktawVRFDL3g2GbEv6B
nucuDJFZeUKVfYyp+dGqeIt1VlOi8Uf26ljcGkCTBdvfMW+OGHAnDVvhfvRWYNydu5eVO0tEgIvw
jRGvLl1ridbJTfTGBvCiCF8vuZVfvsYYDR7wUU9A6MP2SNgjMso+ZZNr1LWZoGnMKk82oB/d/V+F
PgwD8c1dCn80YSy2A87msVt5wEmABmNll9V0JWYIjWKpEFKNsaQJvclHH2/EdmgtzCBiDvxuftji
K5NuHpzBxEe56pMFqwlWOdXxbVjgC7gDMzH54ilJTXGevYaNlgX6f54m22/cG50ggwcIKgT/El5t
yG10t1Ld4FE32rjwtJDE7wKOorFjdkpGK7akNs4MtlqaxujnJ0E7+GaLHM8lhq99MNiu5BhUsU+5
h30pkpagl/CUL57MKi9Mps1F/7KL/MQKZA9AMJiM7hXDZgCUTE4msjiC0D2Jxm4sHZEk+MpttyNj
mBSVVY+amR9JUpvaa52NP6sOozs8XNfecOvRXJKeDiHy7tuLzwNDhjif/AC9s9AWpliH35Kka4u0
eb048CtDntK0jS5oPg3VU2WFmP3z8ImOJlchkTqKKv70RZtmVkiEC+K7syc9pobrTSj8DdN3mQ75
p+6R7c3ZMu1r6vPwDGrBYD1aU5qD+57jwYlOdaWjSbrMbGp/nQT5srwmzaSa8evAuJAtvvaUiGxH
04bX2wX0SLFAaStb1xCtqbRH601QqeVpgOLEs0pmxKK9kz7htcudxQt0njnhhVWhwOay6ShIHYQw
DZGPhm1TqjARtByLSzztwXlvwrMm64PTVQ0HgZRYpPinkKiHjo2rkgzMqS5+u6DsPro2KzDiPcF0
XFk09G03QdaSh8DJIQlrOFXp2BbFfj8VNY0DcZUEnzkFQwn05ZK20AjYW1meepz94xSD5zBgksih
yINj7ksXuGpgP91tsqzUwzJK3rkjA9gxk5FR3r5qPQg6nGNSPcIQPXtasv7Spp2dmmGTLHazsoyT
CGyFI6u7oLruoVH8AcsV/Nm8ZZac+Pwq6Js4Jq/ywMQi7VkeXYquS51F5XnV+xjCkz8jTky+GzaH
p3ziEyBtFbEZ19dRgu+4lmdZ8d2iz18bndnD21YQBDSOTj15MS+eaKbP0gu7gA9YIlyqN2f+rMiR
MtME1ZzykVER+fBFf2uxLpNOXUOGTnEKzeQC30yfSN9rHWJtiCa3H3h/XxPNeuUKKl8OR4K4Mae7
JsqWD4WxAyyVUNLXLU1TUJGwODU7GBYhTaXfA6Qynxmev7umfpRrxaoobNNaGNes/ve1509tk0GN
Zsc+tZT8ZNJzsNwt8G4okwMKDsovxnmPe//KvcYevlFhb8upSbmiuf70hWBputuOsslcEJRX4Edy
30r4fBS3hxP1mzAKWzBYXZTMSxj+izHC7d+AenVKL1gRf0hMMO9ib3yEnetoBGZh5afaOLgeoGDl
d1Oq1FycmYTEFCE5419Dul2Ug6TU+DxdkzsyB4UdHODpgWWfWJDZooapu75n7kXxkbHypu1W24wn
PVNYUTfAhdgAFFK2wWL/LNqh8Bi2B1VgKO97LncatRp5FiZoHX1aeXfWSDd/0lnQKpvXIo9skgYd
zYa9XIIFrz0uBhWrHEOaV2NWEjXwVY6xpVkk7O4bel5SYRb40Gfy0npYJ9ia96iNH8n5cHnKxbLf
JenJ9QQJgKtnse6UIc7cplTZITxVy6szOMMw9DCgi3M/bMUB6j+ORMgX5GmNOJVfm5I0G+Qjn2af
zb4hIJsjYvTTh2EzLXjQnA2ZJlnp51D6XhpVFRxSRNPDziyCOZmmUrkQYNt49MpgkU8ANi5M+CKW
IgFvfOGzqrqZSLbmrGqOjMy6sv6fEKeYcThfjpJbUhAW/ixsq+6pOfeEt0WP4jRxavVnxqCCnsXK
6G5vSvLFcFQia2kaHa0Dvf2/fy0xkgxjTHtjt7jiQY3eOJmLJbiyzqeXBKFG0wzM5DbWcwExuVVs
Z/9GxBj+s2c8u8fSlilbGdYyRHXaaAKMbVayuk+WVbk4DXBhwbN5KlaBb6SCbVcBwdvrlfkYbpPM
824Q3aTP8Nj4IBo+f0k6d+ZmtYpqbQPpteK/35PrhaeqoBFySL4M5NBNgbTILcWldAOlRikFQFO8
T8l9H3bZJ2ofseVudmCzNh/F4WiZtI3uUtR2tYTm7LhIngTVhlUxma9BJ5khL57v/010uGA4y/+H
CE22ZRV4CLt6Mx8/HqC0UnC1lrrG8KchzkZESdMdA7kIZntFr24sqY7tVRplRbmmuK3XuFTx7Fte
aH02taaSn1eS5ZRyOesRHUBOU1Mlg+9byeUFmOOn/6cUIEsz6A3AS59XqQpXLinP99dooLGxL2P/
718F6Fk7Yx4JJ/cMBnlVNrlTp+oRD019GlmlsIreEBQ4gP3Oqh/LQe1cd50JE7nHde952BVZONI+
MXZ+BzH6Rs/jNWjXp1wTD9gGpiJe0Kc0EGfuv+ewTVkaexG7/Nne51oGVsbKhIsuSlzSS3b91Q6s
Tf+pqv4oQI8fg+7kSC2ilG9vip+wSG9Mp0+MvEyp0o6+d42WlggL9Spd892iteoNNYSx3ScN+Jj9
bcxUcczHpPVf6xVHYeErNQ9NZJfu7CfGWMlK0fVpCzyCAH8Q2Iq5Eb2Yz7UF2kOrZNHUDxUW8kga
ANnIM8Ju+/Y7GcPmpxXcMX4Vu37FoE5bBt5mPq4PcQktQUPzutUCBBqiKX1T53Kb3Pe7pybIAs1m
tgVP6KuEmYgRNLSq15EM3FjXMr1E+KJgBJuu13M/h3I6zDl8CfUaU7msVvvMDx+LUMyF0Y7gaGuT
OqoWD/dae7V+Rn8QUg5aHzr2vwaRGQB4KhkUP2dJA5UHgDkJAh1rgB+iODjWLAY4ERw3Ukc2hJFj
nW1WbFNH+O+eHwEPQ4vSsmLBDJoRCcxrnCHy7gsSaiIe/5QgCLkOKfE8nz8ySaE6v7xxrnFXFAsF
WcVPwlvwDj2HYQP3xGiv0PWEkULiw25uJVart0YxysmMwETqSZsf8s6LZBaJOEbdZQlyBxfal8Ho
ygobznUqCe7HoW7zGhFh9U0LPk49SyHssrPeVUIu+/V7B4jDdnfbwQx5xWceNS8kcfsqvMr3RaIi
C/qkVibjs5KeMr0SuRisChOFXQ+d26ksO7cxpWWsVolbFHEfATqo+lhLzB+4t2sjqp3j0UI5Djyz
PnVZoEYuNxgnW5xovoDT5wno8TwKQB1zb8Wt5dRixBYX7nna26hmM1D87bi+x1a2/kXL0LR0+X1u
hgg4DVfptp01gyhn58hnfiaDZXDSGp+4yq5gdpalgmJemq/kE3+meye1binighU9c9og1FoK5oMR
kY2LFIzoFFUmDSnUPKF0ZosZ9LiMSpEm3S/mqVJss4dngqLKYdILCJzfuFXn+NGYBCrIfvo5XuGh
GDmG1WNYLWJL5GRg3L52Vm2AFPKGjVnYoOJkijIo1NdQANVGE7czruQwhrc5lL1YeNYdsJDkvqwO
MznRjgWS7KuPGNCBwcsmk342O/LCw1kvTH90weSck2ya1M+u1aQNmKSexT1GShRYS465pALF+iAz
BjUVlZT+WkHei5NazK0LbqBpx1+gY6HD/rlS7pppyRgK6X9pkygpGMtRaBWIozKPbxzHN0qcTSM5
RIdk9cVGSmJfrj2sS1592nrm1JJQskEuEGe/Faf3RU2+Qq61TWr5ahTZGHujF+mIxjAmDDcU0jMk
yHuADbN35QCzmMNzyvyW12vBZalBh4FLZhN0gXo/DjaAnyeJcJ3ZpmvmISgSM6FONt7AsSRUe2ha
rSaSQWK15EQ8//IaNFGqjAyx16LhAXeJv2Lx+uOb0Q2U4Ap5+ef77GL7wQRC/kb2KBnon2hA2veO
d3mZXmyQ5BzKKcD+6K24+yzGlg6U/2NPT2++xP4b5u+JbZX/23nA5pGvYS0sXQjfTfhqVqFc2PCL
3Vc5iy6kFTfsnugMx2udYHw6X2NXyTHC3VyzEwfpN8NiLDjSX77NRXpPmP4IB5Lz1QS3pjz3RdTq
+Lgwu8KTQiMvldm1/i8ekDPOv3zZFWWXA66Y9Qvh0VAMdmpoz4IUe17c59j7frRfNrfMmxzPzitq
aDQ80xuoI0szIMJG3SKJB9WmukuKGPjArqmgizYpIFAEEvSRQjb2B82PjBjv/ehXrRCFoupapufm
zY6iw+a33dnJiW+oell3iWHlWrO44OgucUFzqPH5Kfr0GujS+hv3caNSgKCr71bmXDwFGzNROPbv
l1eODkNmGCwAB3dZkbuG0AAXLu6LDd2W66YC7QbtiSJ7zBhxUxQ6IwTO59lItwBYPZaJmKzqYrPh
qCd3QOneljiBTZn8wK+SLu81msT9A8KicxeVN8Ac0ypq2MXyRHZrzM5Ot+vIdKycp39obJffLpvc
oGghzI/e7JZ2pa8LQZmyUsPT1TbcMmjPUrP2LrByQM+izDjKv0YiIeohB5QbHyWaJ7XElL2I6Gbn
iEXj2ao0OU0MfUtYwOsdBgWAHMW11ZNXbpalhhF0Z1DTHgKOL3qDabOR9MgOi0qzcviEFDM7fK05
P2laP5ja4dnWCCjGdUixqZ4TBCKyfcU4voos7QlWZxLsEQz8NsBr7lr1pGPM7rbluoZxugbJFQWP
lqosS6RnWJRIEJHCElGZtxzar9Exb8xFNR2jo4O1fMh9UYtD2zyVGy56fQDPv8lBguJv/TZqO0Um
zNxLJvlEdYSENDRdq7n0u5yx9vOiCTQGZ9hCzy/A1GFqT3d/K6ahd+YvKhKCygU9xdKpHHHdryEG
24sqOZuTSKeZYWyPqQ58nZRl38COP9fZndkMgchx1ia74hs59qyGziy4bh723lUs+czec1GPMzzs
gKzu49DWYrBWCqLY1n8v7bRbY0Vic5US0RrDQJMtCDckYD+xuuiEJkn5s2Y+Ai6KITLZz+5BpYKK
AGqTrUfklb1e7h2CtT6IO5O/Jf2hIhxrXKnfMZsRH+mbrtkfgEv4N3K5etubmvnZsgpB0hedyuPx
E2PYKdJrX5VcAbq6T5jHxhqH+JFJPKvi2PzmxhJJPCq64U3jjGNzSSsj/lJlGK/TBg9BPeFijfBw
Qtl8wFoKA8nOeU1n+lVb7egqk7ngtoyPjqIwTLPlZBmesbXUc45gwbUaKZxVrcyk8Rk9mc/VYp21
YMX3xht13qtUpfCBA3OVZ/UouBfFWmT7WT2h6THrwDEYcheroerqt1A3LjREXyWE1Tmt1XrOGAK9
Y/26TnZhCCBe9OLESMmmutOgR4Ss3pfVGjZRGgfV2k1e+mQilpkcQB7plZyIoosrkp5taun5e06w
LCIrM7x3+heTu0XlcmkCFlsF117rJgHd8PcmVv4puuPGTfCPF1IOnwdZZbqGx7M9kvyLErYcMdXR
oM4sq0K73F2uy/jYAGd5dLJF5OOntk3mUbBqLII6eYXRtJ331Fy/3BsXCxUoFemBspkPlBtJi+ZW
/Pa/adKC4JvqOwcBwprLRvr2s9KduNGVJ8G6x/2iUv6AtKBrf7vJS5WpmLw2ZP6wA+n/OH7GJTdp
Xkzd7A42V8vqZVyw2ecFKZHPmEmWU/E2gtXizwaaFQS+0IKW1SdxXiFjuaroQVu9dak3vZLWIhkN
oZ90iqOJfxN354ZkGvWVZGp2x8+V062iBPJvsQH2D+puCe1ZDd64XoUA/R4ujg809JLfuANBAZYV
KZqtYnK12IeQW0Y98SgCDlHed1b1lHvqdoSTL6RDxO/YuRdcBujdV+hmyO5HTZNov4Ri3lasU7j/
jtiPGW3iWtCegBtGE6OfPObjGZVlnuhjeTOXs/0WZTO0KGg4JOKLp7uOO7fgMlGZR9DglAYStnCh
q/w8/ZWeiKnCYwgceyzFHoeJW4hWObe+y5P1FfsUJUHB8dWocnN1vXF3beszOICr+fCnjK50i/h8
zRllCVFpYV/j9qbMBk82uR47DclHlw6KTymR3Rh0P1U4orEbxKMTnwdd8OwEcOYmAHOCiLbdOCje
eTxx2ACA0PiDLO25MbbLH84ZT5PfqdiFRM3rprhqM0MRljqf0jCWaMm6oKUx6gY3BHBQUK4mq1NR
VcvAA2m19LPODg3lxm0sG18C7Q1oZpx8INlAFaZkAR82IbovShabHm2AdiqTar8I6pUAhwt7Jkn/
7vBbjRi0oP8rNQsWmvZv3jjTTTHAr/PEoGB3lCddvFmIOhnXF85JxE19nq235Rkim46pL1JfjhaS
lkpEHyt+STim77yCbkcX8W+cKC6XI6WnlLCd4L7H+J2YwOmhyGTeWelsvfy3LNhjmyi7QqqIskBV
DzUnMipT9/g5H2fJkDbRvNUPzYhLjq+55OqgqeFnkG27YiS5c18VDRPFH5S3cefCX5Xgkuj17mrH
PmRa+Kii61lArD0feM3s3MPjoB6w2nR7oPjc7Xo+Tu70/rrJIzfPrObcrm+CBMHNz4lTdW7zSqtq
56AuMA3yy798NW+R8qM4a5aI9c4bdXNbUYS0BAm/JKnf/v0EfsWuM2/aQsiWn0Lqy5gr8ZvvJ+Ue
L826W7kB/Prq1WV7qBa1oTDdAnrnsOLVOh5d+EmZCrZ6kag/bIl445xu/u0zfwwGgcugPbYYKQo+
ksbLnoMl0Geg+qj8f44XDYZr/8epdYXgIVvam2i3pMC0Jc7JOPpYq5G4mfYqj2EjUb4YuQXcB3gH
tJGCYBn5/FplWwjt5IZM+PCGSgfBn++WJfBF4SiDwyOpij/fTbbCz7vj3QjXMwDKrhRf7upZR2WT
aHYcT1N9YbWngrlQ4i8138r02RGLIDAcQ9UO+8h3cR4xkm/Zei3RLcNHaLtsWC0vvUw62ZK+I/Wz
WStoPmpPKzkos/p2qTscY5niGlSfNm/0E4dMGP3ggF1/wWGZjjbdycqRKE+5FpIyY/BbV0ij5yqO
HMhBsanxrTLksgzspzsYDwHNcAan8qOcCfP15xLI4p8RiW5JiOpGn9gFOlaLA0G/1aDxF/wDYtPl
oPsyMb+mjM5qjMJy2V1EiON8FmAcfWJ7fP/lR/szfPoE9YAs5h0oJ6QgzCbOGnMxHLmJw8B38kTi
R67SPGyqmsK5b9elBwCH88q+Zt14DmBKBalyQ+reJf0diSMbRI/Z3GYD9Fdr7LJoAfNHIa9wt3xt
8v27QNDFFhYUK9m9Heeg0pycUQcXNg923/sy3aGFwUYVL3/w89n03pCxFNe9uQbVI1EV7/P9q3PJ
5Un3Pkz6VRu0A1HLRODS6OgRgAPkjXz5ygdaQVMs7uSL7moekqiKWtHrVnKi0C4ueHZI5aKQPcAv
HumF9qTyMV/S5bhk7RqRLYIkyxJhShdemNY2szlGJk4NKGxDYEVpo0LkP3+JDSTGL7PhGv3nimqN
5nbL+WA44Z1EZbcYqL9CEZX3WF5EXXc71JG0duKOAVGNzb28x3zTLFIC/U+dM/V7uoY7bVMnKJTC
cRZ4sZY6nHuKfiG2dtGRuoWy2mjbA1bQrIX/gh/15FJb1Cjw95EURPDvc/PyignBJixbPWaqUTsY
B7qf93asqlbOp8D24JptKT6/xjGkI1MUVXaMBiVLZBYDrrP0uHlU7dg/U7T1dgqqnfWaL/1lfDsH
dZM6ODfR98vNZ8NoegwjewxQjgwDuYXEetbkx/vvs7aYwieQw8nYfJ3BjevPvQst5InTlyZhAFjq
3aWN4T4ytkslPC0TPnXdsjNNvDXdvb2vMDskMGnbTgfdco/nYYXbJ4k+q+nEjA2PpzHZi0NTgOck
cI3zE1z6rIsz96O3l67dZ8fZFZVXbs++TFohj+JMqekyZxj00ylMBpjM0buPJNrGaMl8Ts3za00X
bUG7AHE5loBeCjXhk77/sDGuFRddMCE7eYtO+Tna5txQVr4odd/tOv6CDAGEyj7pWGacboOUBmA/
RWCYa/eGk4LX1pui/C5kYIiukXXNpUrunb4umRej7s368Mii1JskP467yWdfRdbpZ7+wXHRzIdyC
OMEap3Z92qHCW342birtGU6nmR9R6KQsC1OUkaocvMwA0ipm91usimlymsI2DWnG3P6Bpy1YIIkX
DlMxcWhwMz0qEenVvheYOOVOylMahIo/7ycoj0LvJYyjBFjVakAUWZoW7nlXT9WhV8/Z374YH0Z4
NfflBLQtN89eiaPgns27i2JIVIUBuvx+YKE6gYpfIs9QIu1o0G9JJJ4wfHqggYeHRpUQaGdB8C9Y
TuObTIOmTFivbB821Er0p4XKY+4bLhKaN8eGwN9Flp/GvFz6VdVCVTtF10auYlOD9xxcT8YyUaV4
NwD0s+PAgpoXInsv3tzlqKEHplO+6lHVR40zyvzu6BE10ogcEvKM1rod7Z+s3J5l6B+LpCdWN7+H
upzYMo5uxKyl1We41R7OPDLUESolveHfSDFBtk/9bfwd/BFzKUVOKZHeJBBQFxBfDJgHbxbnk03O
3drTu7PgaS3kMl4VCWuNMIkJUu5PZAH1oGA+5vUu8eyR6zM+jFK/zYUQpF/yTh/rTyydqrunyfeY
wl+MI4ot/E+vDlqymduBPSwsAg/1M15QMm1WR6l8W9tqJxnsgcXjV/+Dw6VfVadcUBUytKyj5h4G
yD2vbIwgcD1WPvODCanNgBQzkuqMHJP/Iq4kCN3ajhNz4a8D/Yzj+/2Lt27yDBy0cFwl8qsWK9b/
HQweGSr0bIfMz/J9It3zRDeHKTwMzYhz9iglLz5wJmNDxN8fhW0en6iO5Ecxw75t6GOf4wwI9Bn6
6ZqHOEblJ86BM1GnTXjxnpOoOe8SHPx0xSFz3WPrCABVYKqU9drGIlv2jFf0w0tU19t+Ee8rEPFs
SZiBf6ACIg6k+PgZ5ChSHhEdpvLaQQXEyiQLq5iipzrpCxNbRpRfMVTjEXN6m/YoMRlEsxZ/p27O
xus6YgHbPot5zS6rybhZTklCu0Pmq/YncC6otEvrebYffb0PozIThTT44hErrFnbHMyGoVHMktG9
rVzvoZslwKd2oznCyjhZceOC9BnY3t9PxEkedptfIlkPsnmev/OsXitfgKHYZuRi1RMu6CYyKdDX
CfetDDdhpEJi7QrDvwjPe0BVd8gc/rrED9wUmc9yTev3d8Vy4sW7eKtXJZIt0gnQLErPBd/UcZDd
obDLb7IFVEkd9vushik4yd26ob7TvrIHLbKXWZaM6xRJ+rXM2pcUuibvliZJ5wP/5sBEnWBcMj/+
VBFrE9j9z/9nuEggUFyrgndND9XxRVSikNFzuYju+hoDwxQO7nVsZt2gXjkJ+Eeu3fPF7Qsxs2Zx
QACTA5j+gyeDuds4LZDc7HtZnAuUIe2H8bIlLwBRN7DUIzvpF4ABjYqe9cFduxuMmH/FJMfdr8Yu
e95oMMfEvjx5poR2A1mxucx3A0co6NT8KhTFFqTvYM/bo7EAcqLJRJUxuJ3SR5I6tUYYUHIkf+Jl
EPCKaifn7YAKKk6ErHr3KoZO09hBePa7bfuOhv3KItaTl0W0Ci/m3MjNwXX6GziD9NOkPU/yKoKv
KyL/yKIukR83jJj+P++Oemk6NVv1vC65W2ZQjSc6CMtkjh6vX92xRzJpVM0L+a6o+hYO82VTwYmf
U+JHZHtaqIK+xIDMS/EWwyf/boxDCyx2/MvxOuaQelxJCnNRGRjboKGK9dISI9jkicy5BnxYtIZB
ll6j65zY/p6YtHoPTGRQr9gkTE6xbLRst7iFGvB/qq3/xsRKQdchFdLROw2heOICqt7L56SUi0GO
6EeMlRTxlZxuFYDYhbvmixkSRL1TRHuBpn5IGi8IOVtG//L80qa4aheOqMP+KKeDA9cYr77/gIrK
2E47jBOry7f+fnX4ORJLE5Xr6geG8+WQKtgSdp7Bv/CVkaIXQ2WarXxF4kT7V2+050jkWv0+ZYd5
2FO4P8lxgcJfUMyrvofvONauz5hImT8fMT3dOsCeToycedgXLOk123tQ//C2d8OdfX695tw0lW/T
TpSWq/3j1weQfDlkmvSZt6fAUe7Wl6OTjzzhwESUmUanoY5DS5FnKeWU+ftCoMbpihmxhk/Wmudl
kzXe+vel7Qvm//irh4IYtyJWN6VQW4NNy8fHRcghxTNE7joEFQRUKpwUZxTVqx/qU3t0MifIwMgL
LUhrCJPWWNbiok+TtjS54QgcRXBJz6U9lGrlML+Lb1IrANo8kSV8A2dXughvnwauU/LPsXfMm4iV
DN/VLHOYeTE3GF8I48YhxOTxv6ab3ZPGFDY/gK+gxOIybg+JMVf/4DApJOk3PfJ9Z1eznU0BsADf
CE31xl9xsyFNQfiSBNG8M8HNCZ1cHsA0afglKyZHd7hG9QDFR5eW7i0BUa/hsVH6F4wjdeMZ8JfX
SdiqUVSjf9wzJtnxeEd1Z0LuBQc1Pt6xZb10Mg6CLJQ5YZoMLx4IzMfcgw+FMkEufgarqYcob5tq
Rx9AX/6HbtuV7PmwU1XsrkZA4sijgrkyJCByt2mpjO/PJf9gykby9ZIFEn5qouEc+150+9DEBg17
JuvB/lM9COpBKRkBLPYtOxAFE142Gt9VOq8BBNeVEH1ez5zk0sR1C5Ir5h+G5fWD/kLTK0+cXoqH
9H6kNBxPUkNpyKQbOcnKsoPvZolu3QCjsAgdzwUfkEcA40e+qTrbY0QdXfURcY5pYzghJszMJl7S
okC/GlMyvSZxhn2WDGogkzZnXMfSAR/uqnJ9wqvabUZscq4nSU0rUQKS/FavaLxmxYZrZ8KbF63f
IU48mqUO0OKZXgp3Ve9Ro3WCTaz1HWmcxxdcr1XZ4RymRZG8+Atm2DeQ64OGoKJGMAiYqtaa8rw3
gSymN5XaVtzfCk9wxptC9IJJbVWnHhACyQlkVEf91p3OFtLcLVjKG2PFnot9oiAngjjLsXPTj8il
A9wXgU6oRBHHWoUUbFFwC5GB8FFyrmXOp1ZDYXSZPgPKBYvOAv5p/E4R4sXZ+nhC1Fwpo0cTQ2CI
/yN2y257OTf7HF6/PsNG8Sf7pqjiw0OnYoHQcnKLJWypjUMKrfthkcVMGswm0sWNQFFZxPkiZ/B9
MeKYt6yd4XuLxECV5BukKX1o/1KrhLYerZbfa9ifktEnMrgmkGtnUl8hkYiV9iZNqjD+n0zUjZyQ
jvwQidJ9qToBj/6nGEH5N03SO5P1gWaRhLXmJYQk5CnCQzeP6MsM/80eAQrobzhdGyv8zAFM5kj4
f3JG146+1KISnJQMgOz90OHxiLNmwT/Os9RwTUv/K4Jb3zWk7OtmcON5KoIQ4VDDPiS7j5zvXxTK
1AIP04kwO6LqBME7C7bid4oeQ5T2wY4/QhaBcJoQUBvdPubFZA3ufA+sLt4+ln3xtqgjd6PA5Pfy
g0gWYQKnGA6p8WJlCQYqg3oCEGabob13smvlPGp7cNGa9T8kVb2tmw1wBhujuv3YQYhCBH1Qr0eI
wA+GcySmpSrQe4Yf5nz33PGoLSTzT1E9zCkl9UocJz6RMi+ZDauWyS117Ah8MISyRAAuSuVmnhZ4
c3hGzHUpLcCmA5NE1Q3EtPZCLCjOLuB8xjNz1CdQkMO/f2x7OAGvQROiWPqPPhPcycg4TXAbBPcp
2gzfTAkqgsxVpgxHFC0Rk01K9e3EtUSSUGBgC3uTetcTcq2YCaH9nzEEUdQ5jYDUf9rSvUX8VZie
Vjc+KZbl4Fz/AXaCNDJSyUwpbSiNAMT1JSvn6JqA+lxzr8bryYEQtWwrI4UAvL9etf0WRNsSskeI
IFdMIt0FsLZRXeleD/3c9C2mgc8cLb0xMGah4kFAubiF4kvRlmUEJkKabnfct9kfKDbS4MX9QBwo
EJ15dFgW3s3ziky2jkKGDLaUqBVCjQng4rgeCFFZbx4iMkXIyPfbUbjtO6eKP8/xJcCfvkG2Za5e
Q21DUVI0Tw5rka/rBrJwRsIKSUcAqCcJ380UFHDD43TYWLLbn6IfeR5Jhw6CvMwpsUNmFpvQd547
uIOamUn6qv5W54CGWy/JSE5LbDnxH+nR6tl+dxT2pxBiHna1/RpCJFnJJxbOPddKHLZhn2+qoikA
5Aii1rmxoICu1+EKVDOtR0UUyqbPOCPC6qZR7sU8FgXBQMPaw6dRuVQqsNOin2jGuM/INwr0EVkl
LihsYlRoXUIGBkpLrowTnp5i1MGwfG2GfhLFEq6NCTwGTAAJF1ZkMcb19eBppfaiZi98Y7wJI0VC
adDuLnGquamposZDZtipNG+HPJLdnJ3ODKTU8bTYuwmjPvfNJ4WEX5ef4rR3ioJs1i+uLBEN3qFf
jZtxMesZOdb0XJhtKKihmUjmXVW6y1s90uXvYkXN0AurhSsM3g5UB5wtGQS+ET8V8RDWOgZCdQPZ
+1ItvcyW56ms+FRz2CGMClncesu8WJ2rJOXtY+YLSZv9A9F9Opkj9edwQVVvYS21b6s/Vkhm/xuX
Y1sR6r7rmgQ+Ti9wzT+xGOVcDWp/SxzpxvnzX8i3cV0EgtCWGz4ZSXdLMhifI3gNqrOJ5x9spdcT
SFbHk5Q3DwBl7QcFEdE3PizDdXoDs7berk0ejLBrnQJfrVxjD4eqdAR5EY2AeDP0mrfguFqK9Evw
anvXFSRzpqTF9wtYDKrCvFMPRdzi+6ZWv4vrb2TT0HNhoIwWRdOGiTOJuHz7iNo7nv0d+42eyF35
yh0aN2fVVmwD2k5wGST9aZDpIsnhGxtFvqkbwf68SpkbtXk2vc4oCFs+DsQOrj7+IY0u1Oo42Vis
cYLt9pTpFuWACeXK2FWZHHSJdX4P+pMHEdC3jqTZRm/kTOHCOZjZObswf4T5t/XUZZ1bryFB3wlH
iIL1WQv5GgvMGI2ZVffTdk0SE0bpdsXG1NdmLpz3cvLZuSeMFiCvKkzNx8PUn3wWXPo9UlBcj9Qz
PnOENNmQU/hrDL+oKWOadHvhk1ZH2ZzGVO3sN9sB36Pl+6mlNJldTN9EPxu+1st6nQA/vB1PwbT9
Ed38RsZTC6qC2fDRgutl5CfUtVWGd/MZumyNNh5jhYn/751oiphAZYeCwzs0mYlZGlBjiYC8m/+i
j2Yjj5IDxLxRTcXmf45NGH7ufmqwuSMe+cvXQPS1Q+SmE2owB1opJLRQVv0fCHOYf/a5PwoojLFE
POKjoRSbzboZKrehX9t1Gc8OyX2cybROQIF6ZeARCI31QLSXGv2W/AwUc0Jl5QO2livP/kBcoyLl
sqQFyv80JMRb4PiJodIYxfRIDi6suFz9t727erAPOIRrFeJ9x/c39LIKxBx6Apq13IBrqg9n/hHS
LxBzEURlrlGFVz1m8B9nzYidUzMXHSJch6woICJ8TNSgx2zor7bZkYJZsf71lcXjfrgNbTiro0O2
cmFPaURGpcWbHsITkGb+gsmrkNY2WDlpHePx2L16G+xj6JboNKAM+VnYpn/UhPh370rrqv1DEEbh
v7rZLgDKlypWl8UrXtxL04uVTqCMP4ELyamwPQaypHv/agF8s8OdkOChLrZjvPOpC7IcqZ8Qd3MJ
pIIdFuzVdYbOJlUXR3YAucl8hoFFQdkU+NMli4TgMlE/t+oIvE22t96/bBtgFxgdUy1VlGGEAL2n
2g2tUV0jQUfIOFsT8eGxidQ8N/LaBkqcqWinQ9yVoHBCzVmCc+bIopPpGqt1RMHJv9OfnDNjhyFE
QiHMQ+0LRNi+vduC922vKoBz8BvQNmuXOILgvnFVHBhd+4Bk5gSGbI8qxxUEF+fS2TiuL+ffx+eX
GUuBtWhd0qfwJNiJoo2f4B5I1h03KQyC7IW4WXvXBZkCOxWFoqQdQafIjL9owAIVhqCd7EXuHfMH
qM/mcQ8rJ+EBwIsZgPycGeZwmkDoolfqBg3PrE8EDrqHKnTHyJ2wg48sLi7o2DK3QgnmtbSb1uQn
Rm8t/9DnsRcnCaPXFTnZEUB4vZby6lkGN/ORMEihHQnmYSajHk1Ng+pf3YHC11JVOjM9AuE/TCNG
ho5HfpVKzmWAN0zDxJvKiGGf8MenOIyeySJyCchBhqXy5Ir73BBGgD29rPV+/HTkG2YOl4S5fckq
JxHz/Yk0ks+VfJpydRsPIpqIog2NnMQQrFF+hLiFcqvX10aOXhkM2FQB1FvIgTPw5gB92KjGrq56
6j5Dwm5VpCltQ19CX1o+P6RQSly7rZIPl9P3VLY0pBUUhHBttCBGZgnpZMF1ZKEUFLLiOLbimxdA
F4mqggL3UwVUPyV83mNRb8L8yPjq+Ed1WGBzctE2C0YX8gzup6ZYuChyal5Klr8tWIiv58EqZ/N7
W+nCmzeMgOxWPheHKnmqz2MLAfOkpYiCvvou34MmV/PRBxNijp4HRklMvhl3JDVnzeXKeOYqaSc6
Bh5iuIwB6JMJ0Xy2vjZH9/J4Q1FFvKdvUmx/xh5Xdlex3A8MUSHeISjUsjKDi7NDz064LRRgWg5W
6wir4aw7JQAuqMYOtt7l/ZVn73uD48U4KZOkq5oNfagB8eERhpTaZ9Nu/ah2NZXAvPtXdCoJtZwG
CO2gqP/qFS4ooHaQ32S+KunBNu2n7+8lHhV0P3dS4uezlLq1KZZubtFXyElg7Tk8JjQf3x3KYWdC
eW5fpImkaaD4w4N6CdSe2ChAIuK/gEHpZhZVNs9eRrqd0HiwmUMK7aQhPD2UDUpvs7OSeL0vKfzp
zaPIqRzheIlOff14OxXmILoFxBw4IWkcl9vRE3Zqno+PupdlMYtDaTpqvFsrLXGnawD0ZVw9cqR2
c+D+kv+ZfAoRsM/CNG8sG49DuPUXJxJUrbJYpDY/Xrt1utOk0yobMzEVzRBYGD3aVI/ztENqtCJE
QYUerWEH9krvpe0xyASvrVM7tulV+6+qQGZlkXGj3L2cSCi5KsHke4Ewp8l2kirb1hk6eC+HYdI9
dqZ604qV88GYJ7zw9Tjv+pGaGhZb9nqSzLx10w/jhnEBAoJr98h8VKgIgRGdJprNTPglSjlO/T39
lBezE7uly1IYmTat9Yos7T2FgNnXNMelmox2s347vSe02zc/0sFZydYBLjPtOcA2kZK/Rg65pp72
p2iEI7UhP6PyOplQHTb6WGtzPyMaAvL7I/bKSXcdmyikzqpmSqGoPi3PGWS3CeEbfutts2BtIAqr
dXC/CrJiJTpYJMv+UQXqaw1pB+jQmpEi7tKALMQJtm2ZJ7rdWHR53xAqXe1GAntPRCYynQo6CNjB
PYQjEVYJNhAqEqy/HCHHFcQahJro/vT6ZCjgeInRff8Xomg+t9mWP77wRO+ti9yi5ahbVhk6VTxs
tl1DeEKHj0AxR+loukcPvx9EHfffCvuFmgfvcBTwPD33xinCYCW3DROaHOmW21uR5NbQ083tLX60
rUBe44nqTVMJd/cXBRZuonMZgknnsOk4kS7543zCzr1iFm6kE2VQA7emTRuKvJai/lLouhKdebyl
z92x8QM9odA43tq8W/zw0j+qupv8HB42BU/GBY/IjlU+vzFOe3Eu9iA1BstyZvKUy6j9qm9uUYXd
q5gFbM09nKMZLWMaVQOerOqkQdhYIpgrjP1bGkhAtd8MmnB518K7zoHluqxxpVzsUIoNVlFNdKqk
PP3g/bEiV/Dsf6XIKJimy6/Vn9gVrrJHpBLSsQZusd7QHiKsBtU1htNGlXzMq6h2E0BNt0FWFyxq
DBIhc96TfweFlqMHkOxBwlsfEqEhYxmFo1xHH7ZH0BQi4mW2ZpWi+ROpvFQQDY+QI17eSdKwiuol
48wAijv2QpwWV/LnLUPWT1gQZ8hC6BN31RUjjMc8Ol9ExhNP2KKu5gIM/KMHH+E1u9sG5ERzacaE
4nVRmhLXdP4llbB1vG6nP2dbCv5bKxm8MUrx3P4sRM8dbWLCrc7Pn/f6RdLA60r3llgygfc9K6h4
Se59lbCS+Rkhtp1BiRSm7U6eqhgCBXoPk5HNPZjZcNTFbcBscWkM/wpV81Xj2sPD39H/2B2gLX6s
isQ6pfyRhV5eMh7NGzGGqLHdXXBAUrufqFrWStKIpnVqp3CeTEV5F0H0efzIIgwnagDOT32kdsVW
2xEfehHHkznfvB/kZQJ8/ptpXEZ1Yj9YiUW1BUz1FInu6LtmUHN3GLlyFQwDrm8rDcoH8xRQ0YpY
+dE0R8xETp4pNQlricgmO6cRuPnjhuP4GTfcnpxhtsxPIm7Cj0n3eMpwxfSnfor7IKQo84hfg829
rqDUK5RUho9yQw4s7hGotk1H2UnuSLRwL/spWPaesfVgneHzIHLm+65ootX8/BnOq+XzwHGRJjHg
YnbRzqr8SwefiNAiVzx9SWq23jCvpTykQRUJ0E1Y21GtL0tx3kFkvkOWmUBUjjjrCHm/qF3YRL57
3ExdSqP17TuqiYhgqLcYXZxpW0TS6mcVkXqnqKiqy20AIGpFuWP7lAlx7R6UiqkY53dtwMJbT7iH
bSTtygJZMm6QSG3bJjQqIkikEXQ34zx4ZzwPgK60fZHI64UNOnL4RT/N+tRF3x1v6tJIQAxF1bM9
LSSBpjLzJKSXmYQMHbdF32PLoOH6tGj9FI8w4ge+0aRrzyy2brusXC3kuYt8yNc0Z5uVyhNQXxuC
PUzZs11SIXFJg4Y2MhAOLUZ2V++bUX88OFfGmgZmNlDFMCHqU5Kudt/TC7D1HWwFKd/sZ35Ave8G
z0WA8ZRJLYWCa1YFMeAdGeIV2EY6lbRfSuo0fYs9hVug9bXNN60jh5H8sKrfIqAsApA9uLIg3khf
zBsJCwwrpiidZPGeB9Pj6ODicUhoHrTPsdBPtva1m8RQlRpt1k++ASrt3qgCSiVfkQUmmGMhrZK7
3kLp6nGcH5jrKfOc1YueBAKOxVRu1JXRUvkNoK0/sH+9BhrPzQbW91sxjuvdDg68FMUeREsFlAP+
+cB1bvmWonYLAZ1h8WrDntPaFDNm8HJOEXuwVDpY6KJW9+K56MAVEpPlcjamNpn/8vrzBqxp3rx9
6cFHF5QdOW9CRcHL/loR/g9FA2l5HSzCCISoRkWBr12glUM6+nP95Jre4vQEoxjVzoKwj4eOTH0N
85qfc3s4nAg3I0z48bABkVidE3KwFa6ot9ZwPiEJ0o+jIi0NZaOLLy239yvIeIcb/KRn0cJOiWCf
YzMN4xD9AfWVn7KBu1eLWR3+dW7eIRUdcOzmMv/kYTHkK8e7zcC+yJBKiiFhKzc7KxknNxxsWEvR
b0v5KGbI49rAHemJa2tezOtZ10f8w+TfgcxDPDf8jeaG3yeX9Vrwagai+tJdLmwOQo/s7z1ZDc61
GDg3xaCl4ZyT4V1Y7GLvI1u4c6MV8JtnB+SIzGLx2UoRSSN/4KLyqE0nVekKezT5wFTs3sjkiMuv
F9PjjeAYOBoIXXj4pZ2GEnzaVLERIIIwHkKk/AkoVNrnvxmF7XvE6oNv8HDOdk36K/oP/7ghAG4b
3suXSSvX5Z970ryQV9UOgmxkvTc+Bcm7bXt4urKQh7XF4aLmWiB2Ln/XHSPTf2oK5LOngVnuV9hg
7SnNk+J/Y7vHjzweL2Q7ZMN8FDyj3BKAudsdQIsBGH1MipTkGoSCUMfbA8+18EORDTxZvDcBhMGo
2BOo7tm4GbdlUxjmDTKNj2YN9a8hmpnUcDFKhXuSu/Hxh2zdFI+Eo70QetU2nc0BJz5KCnh9EX1j
Nj36+CjQIOZvqXKmprQBJ4MT8SsKQJ4xLMkKnISen4syEtdRMJQJrPgh3Qnl43demcwpxbl1Q5RR
Wkc8pGJcPwo8NhjUzskEcekYOJbmH8P527KOThJc9y4rSgw3LHvkQXXQbr/nAILMZ53tUjdl4yJj
Kqz3nS2Mftsh4CDAdIeD/+P1EGwZcUqRwvaObjUuxRVtSdFMoikEU8Q/CZOfea3x4zhs2E/HjIYY
P3OYBhIeFrTDlIqZVtiEv0B+1APD3kDi7zAOEw/ijHu/IpycWwW78U9B59XOOhQTYS1ka0z+plC6
U/vIDnim4azsrC6RPTSsuflVg4wi4bOHKmurlCcH0xq96PJUjhrQ1RNUrdqTl9WhEqwdZK6KRJ6t
vjCqG1O96evCeQfbyS4mVYed5N9d51nsJDFb4JK84YWXMS0JWmq755R3A4mpUMbt4i/YO9i//9SB
Rtg2Sf0zkTWkDELZKEkcgp0mRLUWtRHTNjX9ZFGPrJ0MM+wdMxDh7X4b0Zi3QOH2r+ukrq+SlUtl
X/LBMz5rZGHrKU67iaDapO3N8r+LiPtb1IQN6f3pdrttRS/Omoy8HMPdt38QWBPWIBEjX+JgE1yw
+fV5nkKeeoADRgsrvL2U9Iadllw0D8quTAxfcOaOGT6djeV6RfkVj4wOHpgggMSTfnDAl60+IXdv
gte2uPYLARIvakptb/zcjVEaXEPgnIzrNG+l887EKoO8p27ULZUpTTxVqO4HvdUKuczuaPPVXGbc
3nMR89Nln3aX1wj258EJSmJEpc7AqH8l8grhUXIZ7jFG//lmaI3c07NA5JH0wi/klIyev0VSeOPP
hLwXP4uK3DInMpMzqZ/GTB8CE+BTCiIO8il8nkZWUyg4sTRLOpPaVFia4fyP9CPD+5kzGzbYT3Ex
w6meKDfx446xjWLsAd9zrnKjveePERq+DRqWObed01cd2PpT9Wmesi0g5pEmORVTpHHcv7nI506J
YSFalQctCLFCbCduq5EuaeuPCfz4LylyfVceKbhXIZzAaJRh57F+WU/iNTfPgimNC5n94mB60n19
DMqCqglhnsR17w5J0vIzapi3E3nBSeEnOnSss2oobMi+LRfuGe2SdNnHNnFkqtMwHUYzOBbJWD3J
mb1mU2O1i6WCA+xl9mDcFyApgoeO/STIe/cemoWh9hUFZ+CSjnSzLkkwVxS+Q63x/0XRcBBzzs/N
PNvHVS3ZAY5wOOOxyRg7QUsxYotCCp50aEH+vMQTFFgfZ50wFaKWcjgnJBznqJ5Uz3Yg9LE/S81H
oUX7wPSdXm0AiEhSlz/tHI7ngCn3yhYLxuh3ERYx80FWZFmtAUH5nxhAx2uBdwNDHc/3mxuT4IwM
BtI1OUq3kpNbWbKpAn940jSON81ZvKrpAGJ+geLV2NrzHXvjheL1cQf1i8Et8FNlMJOVNLDlKopz
v3+NropcFi8tQzRal9O3i/2rCFL5EAOgSqe+5h2TuZ8Kh58+SOlIkJHUGRhlH3fKQUke+YjUFIJd
XfhZGZJaK/+ogz6kJtTVGMjANT5G9o5BXmNdo+d0SenUj33sinzb3ic6PxJBEBvg45Ak5O1xVey8
ngHXgfgv+lqE03Uaw3CSfYHezXa+7RuTcgOh/A7AtQ54no4DQzySrXXcAMxIeRugUkpODZr+uxiS
K6u8xxPIuzKo05GgbogyTPbCxjg5aM4bLeS3D5FGK67k+c8Q6LDI9W/1TA2375gmG0sv9cf0O9O2
/pXcP4g+wY7h73rB29fWwNcRNUYU6vfLpiL6cbSbR7+p97cq1ZU/cYPaOpVWwMIJ40nqGmntAH31
WfSQ9GHL6FWd3bhALTFpf5r9KI0Hw16V5rQ7rB+Y/Er3ZKn4yyYGD+zerZ4T5EFOGliNVMJxJNtM
Fv+mI90myHP0UBoDrsPYcR+UTOhMRrspO+uan/S0d4oE99BSGuDo56S/KT5G4/5dv79+ZnqnYDiW
lyxbuqg+gz5FZy3AigIHma9LrDhvEteudv87F9eFRH+bfrogI8h6qLMNVpMkUa2o333jyxx8VMzr
/3UqLTiRyzjkTGNhJudaXp/EcrNEoN8qMrgbOvh1OhlPQtYFITiuPeEREplgJuj2Orh/Ckl9yyS5
nGguCFVxO96pBz4cx1Z6PIC1rUb69wtCnO8Vx3zs+NfqI4Utbn2LKeSc0wehRm9Bnj7K5ln6ieJQ
e8fZ1ZHccY0HBE1oQncuk5AdRcH8TvWMbZZ/7lMDN7ihg6xAFv5o52KMMJ0acsxXuFerhxZWjMGP
sh5VWx2S0xSNvybIWj8Iy7TGDALq1XND8arnGhRZ60SDXVLLNvn3Kdya8p25o6MTLb8oP8Ylu5Es
B7fK33RwhWuRdWqeAO8CrtQb3u8365p5SzMsakvvA+LaSFvUuYiWh14+c3pKSPIwfIiy82MSOX8Z
1IS1EhRw42ZGY5mjhRmwF4bsBWT/OfzSMxwzOmOB8PWWB7pmCo+J5VDhYnipu67dxFcK/UqRIJzk
Smr/1jsg3QcaPO6M0MyAzsl0leQiDXzHRekSgGHQnyBEGUX8RJM30yUUMtt4ogkrk31ovU+yqRH5
87p3JfaM2/+aLQsOn7UmhLrHFaf0POUkc7KeP2ooTd+AxFxbEJ07HnB7sF2aua/0q2Z5EfCpIC0Z
tUvYvdnmfCVkf1DFAly1kNVBW82gmVMRUAp9rFSARdQumUyIhTHyjLnooMwCHELq7jNrLI2fX+hx
UDbKESa01tH4Fx64qeeq/eKwnGKyqNYwu7hNyOIkg7iYYUdpbmfmSmxG0+z98c7sIgCMMA+lL3bw
6U6UagAsQM0KRy/1fhxAuyQuj0wfpGvPCN7EjPV72W5+xul4w94MvR45vfjr7sQ/6ktaoNd0Mgzx
EdkQyalVDCGEaXSV19YhcIHyEX+bNSBl508mWWAot4/XRX4fubblpDYxGc9yvORY5NiZajkxexYF
ExlxraP/Z2oP7qZt7mjkOdVphX/0OGzq6kz8BZmU5T6STz4pCrAQUdBHtwWu7id2jflDPLS4Aey6
miJ6nhJTtXtf5QsJjknb+KabkXYd29r9miTvy4fB2WkE2RrUyo0ISdRozIVm9YLObusP5D1HT0DO
2Lbcxm2wWMM3dA0nPsBSLwQdYZ69rL63u8O3+NGj1eDnhztmYZcXLJYJgJqWaYAF2YOg+tL+slyG
tpzvDVEBp4jjn6K5VQEc8zefjJ0eKmzSD+S2ErX6N1sn4xILhetC/OGFgd8fGcsqnLr9dVfXFwyS
mHkSaQ/eL0PI8DgPFCJ567hZRDNTqsa3WQRvvx8TJRMrF8pjzUsMlmOZKR2FcoZmErqnFIjQ8U9i
2NnCc0kzfQCtgNsVjoo+YyidDIt4oqmx9foCnwN6Jk50PBaryRh3kFWRp49X8kYmVN4n0YR5dn+Q
vkMNT3Ul77kpGa2OLQaZXPoblYtK6dp5T+2eP7oEVoUgoUox63niv1MelLwm8vvJogXOSJtQMn4X
5IKbxgPJpG6dJvmy3iRvJlj1P+2j/vtWWRcuzKbrwKpZ4SitT3yxmarEg6zOxW/o1r+w5OEVk7Bk
OHoUSRCYoCYBdQFLy99qhmfXKpukq1X8lLMx47mG8VgqC3R/dH/vglZqQUCcS8iWPwW+LFZ300U6
tYAiOcKU8P6spqrt91oZZLBRjmFuqwKNmNipsCR4FTCmH2W9NjneG3nAy5DfZ8H0K40C9q98UuES
557ab4HdOpTrLAlgIWbnwFuFdaSiIJGzHt72kN3OpmFDDjT6LGx5/Q/ifF6EXLOOA849p8kbKuPa
w+1da+HkpOOGhV16np9TaX1VwwSW958Qs+cnHc0yzRnjrAdaJBXv3SSNtYpmqvZ3Mf/+mn/7NPCi
Numa7FcQrGrRb2GUVj6AXpUro2SrZ8f0uHhTD4glsVvvssx1hm7LYonxqzrBJc8HpqyPm2MH6SSH
loBBMmKStfJUpiIBUajtW8MAdI5oIalwZt4mRqG5OitxVMggLfcJmQJNFsDZMTt9Jt+DmP/eTESA
lKvPpxrsgWGcvNAT4S0CqMBYtwhbcI+XW+2DdLIh6rsN7P+BxOtMvbKKhfOPN7W27Lx5B8aTehbc
GqqRfuMkFGFRlnEaqYAo4GeWIdey6GuAZ0ck0FiqykuUgg1DjHKrjwo8qIlsApNVt1pWd0DqprK1
1U6T6bT6eS6YKVCuFxO/n54OlQvtfqv4OkmXKm0Sxpa9kFISXFPQBA6z072FUEnSDyejeTsYUIVU
/UynksjMqrl0enlpWrzghj/lAfdezy/csyCWAoXzsUdzpX2CxLv6JuhyzW3O88Kvzr1XGl2z+1Ki
VzUdSJklihCiK/GNzMw0qiTd5eWmVLf5cOhgDsjSF6qF9zE/LikETvWzdvm3ITWQi0WN/ZaOAP7J
4akx0X/Ja52SNz2Ul20x3IkGf2bF2ZteVABeq2wH7DQ07APP4I3aoq+StfseSUhQETMr14/qB2Gn
juxMZ4rtFCPa8IXkKZ84UvflKs4/Pj2Gs2qM/LEebxoLocMuaL77xeBZ3DDAUlz9xSL7kKpb19aS
T2t8FwDeUZO5omwoL0OU7VuiElUVs0McZlpJYlUshKfMvHxkO6MXiluFae2EUUahj0PjWq8ax1xR
kwUW2ifEJdrrvxMxr40XAvtin6994asAKpg6o7HGjY5d9ULUdMhJVC4sMCK/1GVUUL5lhBi48y2c
LwBVC2M+f0lzpBo9U+3NG085MaI3vXjBGWTrhPZ6EDO0SNAbdxz3BhYZCxRkEaSUFsRWX4YhvJuO
aHJZpLnahee4Tl8z8tohELd/LM5Y6V40bALqHnuqFi1wpro1PHorqsQpJpAa+jo8wNkHm2xiTKzI
yrFRNhfS0nLsrKtm6+X2LAW2wfw+BUI3KalW2+Wjlm72PoncMJPlNgfL6c5L+3XHQmlG7kmH2q51
aG/PWCAVngRXQVKAYeZeqqTPhn+Z5rXQLguxgTEOz4FZjVujNw1wm9nn0mJTZ+EPbnLw2IHQpwFe
Q10faJTBrLc2jFXSQyvk63bOYcKMHrDaCAkGfu01LKQNljmAPMZH9H6MjJ+hsRuvg47iRzmgnXQE
oI4xp6n+zIoQ4MXnhTOA1sej9tVtcB2iwz5yhsZgsFiB1XVMhXk1j2gSC8+i5CleXupzaTeY0OLz
1e8UfGFn5QBzyg0OeAyUo8WqUHpnTH6KQk4D/XanjflCaRPUZnvwwh3Rqi0K66TW3Ca62V5oahP1
Itd2iPUVAc0VGMqd6PVf0jdMl2/lZNN5qWfD3FSwoz1cxrRnO/L11X6OqAWqEeL4KOaEAzpYOn+J
tnuMDXWSEMdvbj9Lq9cIH1WHOSqn4v4ne1zKyDv9/7IKCCfaISskmugX9+iBkJryzzH63lG6R+83
ImZykSSiy/UyIoaiUHb7sHOINlMrmIzfXgW32PRWehWfxNpJEXfnqyK7XBD1EL/T7uQi+tEXMR7a
+HQbZ6G0iOPmNx8crQJylV4j75WyI0XV2DF4OKiRSb5oCruwongOa4Otf9XSFKI9R60bGja+l/rD
LbtJTMjKvuzafGDhI6FvuSFFsadxHeHkcokAaWiCJbmGfSYhF4wbl+30oYDnzuqEjhVYnl4eosDT
DeeiBLk8txpopZc2GVnme2XEV0e4mVZfNhcvdsvOvFU1Ycs0SlAgZy5kAONQHUQXe3VafLqagiDZ
9r3nYOH/58g1ahKuzQzofDeslISz3UqnOZV4Oumm5Jnbfdgl6yu7HkvtfFI2cwd6xVnOIlXAlcU9
K8QMeR9Rg9JH+L8t6Hwn5Rz0X5Cf95QTrmrYmJRR/62H7qJ/4Kofo1qK7JBprcLJsmKjPI8HLWHk
rrjqv96wm6nppyku3/IGnHJYGCbx/gzHVFo/s3cWY1oEGUSasfHcfXUz50r3ymGJB59kcG2uBLT9
2I/jFytUKXpRlqj5Ck6GDLcr4br+JUWbwUjFlHTTjQ7MOG6O766nX+I5iVp+/CsFF9o4xeuH3oZ8
bLEPWaU5RIXMg4AJtBA+EWXTzAZuxmSnPGa+aMBvlPugx6LZRdEeGGgojtSguHF5NOsCfEQE8uNJ
LA/lT7hnHH2urdBq1KSrucaEgmw6lltGL9MtlzI7MjWqcDGIUQ6PoDDHoeGTJfTC/sYig8B2x8Kb
0lHXdPqhk42KdWNef/zPH/bz8UMy8s9D9i89IU8RhSndLzxIRfBpJ1CICxonNslYlywq5Sch2QlJ
kTQJDIkyHFRGr4B/RwrlVEoUqHHuMr14JxkVVR0DRmG+9se6WVuO1NcKRwRWWe4wsThVG82rOsC4
5r6scMTrnv9sRmrW85bHOnbbwMFTxsv4S0U0DcaHjxL74d+A0joonAYYSAZwpA0Ax7kK8Hffne1c
5z1SWE+EM21Lc8c6+EEdbTxkzzp8H8qCyASaiOc9c8PtXYHMlU/0VwkH5pESiCU3hRWifJdGiPj8
YP+mK9eQZ/wKh1o9OkI9u6stiXd7X434jFIekKq4qDPbqP+KXlytU2fbM0fMM7UoYFwWobpKcbVp
v9dawvBkv+Yw2JTbKaMB5YoOvlWwWUC2+D2/pdRkUwVUOwZXxgiUzwT+kSVwe2TQslLolvo1kh0Y
2RtKjs0290yHCkZFCXIncX2KOaVM5xxHp/khjCQLl0tqL3QkX63RnW4MEns71j8e6AD07L1tDasr
zRXNN/5w4xZNukjA7Cs4cphipEM0JYUFLa2gyIJCtUvdQkoWGcx+IIS71YsUsEf/aKu9RhY6lvY8
/CI6+LQjj/LREYe7q11egY1PSTLoL4H/SHKcBnOATKwMZEIz+BRxwnA6p36r0hIMoT0qf+Z1wDot
tZJb/VnPf3cvm1FAXIgmeoa9qJvULGcP5zq2QCJExVPQkayiG0DexBEOzdDOtf4+K2BST4lXF+j3
93uRD0MQR/dZ4mTAiV9pN8JtnEjB1CJvrHC6xAvuMZ+RUy2YovrEkMqcHNz72hI7emgs6c69Qrv0
GwykUdI92LhlY6/32lrVaQF0qi8oicIhUTBtk9caugUelaisjWM13j77cJhN4o2/C0kUXfxNOc2w
i4H0v7WFgULAt8bNxkFLMD9wJH1Vr77TVrWybLZDMVWDpr203vxEEjqIquQ1TdAQoBlwnJooIJ5C
Yn7BB9TLz4zIQXGWAImcy0DCdPff0HeyXAbI+1UqkDCvk9MBwAxb9L7FqTSPbucGkG9afb6FQ062
m1iQh2nwq0NcZMsZ3tfY2ipVQuUUHE9zZbVbwHK7iWDWuvBncCetBzf+97Gb0NrpVBgjgrD3j9YU
lCsgYdrcJkJqBLc7s0m87O99WlQqfTWUmkaQEMJ1HDqH6CdHkfgdwRJq7VVpx9xnbb0SUel/N5+D
pJJliBv+zW6ZszcAWrYAc6eYvnqzVpEf966Qc0lq0tsh8G8mVwI/U4IIOqUxizdu4NMSK6LXCA0a
4G5iCepG8t07tU9a9ilp8jXfujvhd3v1SdmLZ30ixRkunNSHndhPkwfox93e+2yVxpKN4XpxhRMJ
xw3rOjX4ka0YIJk/pWzqPMSONfIocilRO4Gh1x3VwC/928fWOCxUstCPxP1bFC5ioGaj8ryKZUPM
pYPd3zHb/XhadaFZcloo3o248qE72EvZCefUiWOFevcg3zERTqZ8yO3odPYXeqUi3FLXivgGWf8/
Px1r5zmH3xbgVmmLTutsR79+cznjCKoAYfNPDhZlmXyPAjDArvvtQRGpWSMX+HiFmFjy755PlnIS
omEkWwpLJyP7FSgmGi8VQDKTo1wlF2eP0L4k7fLpRwsG48/I+K7RviYYKk1OGpYxq98CVUPE1S2O
+VOoo4QIexlsTQtFRI/r+yzBFOdDbLlLONp0FT8BhY+5XQYZyUrOSP6ESgHtC6X1Ws+47iWQVBWF
5kJy0ukKRMVK6kG0H/kJz+FKziGoLeGMQFLZJaIkqfHxlizvHixsZwQC8SxBCCrqaeFCD/YAn71n
Ao9nZB6rnAT5wCHPHJHmzeosB4zFp4YpNN/12UfBsd6ucPr7CcY7J+m1xDthuh8V+jBW7cR6daDx
UbWPcKiF2osU7WRoTLvxFq/pI5iKO6fkZ6uTB7Uwqy28gdl4rIPLYhQt9nApppfwGclHVvgZfZca
q5DqwJfKQKz7IZ9tkzN3ATwbKB788PWWRtLH4nj7MqIXCjbyTkfKpS8KU4laWOnIjo2GFlJ02zmX
9FueY1Rz9Vbf4sRATInOzSXXVOzIVH6AwG4SRlVfiOoOv7exVw2PM1X+isKG7/EUVxMamIgAT+GG
mi0Mc/PpP62xKrG7QB5xjTxxwKPwgbWuCJqt/a5L6lQA12X5egpetOVEgyrV0RHPUhPGngQDfXa/
Fmmax8n4xjXiJmAaBbhQ2MyO5y5OxtSnAsmCbvH0sGPt9o/LaWCyKaKhKlv51qFYmjKvx+xozYLN
44RVW2Lx3AEVu8AIitLdelotxQ+mfdxxNVBpdN43gLIQWBXa6/cs/ve1ezN5jlE/XGK9Hqwy4b74
fec+HYc3qC97it8PCAvNE13zApjkG7No7ZF7Kxv2MjrTI12APkk2KCB188g+PQdy4ZrH7+lHIFhj
2WoTJDKI3vyTepCsR2Zqp+UcPxsQbcyYiZibgFNDGXOT8InAKTf3H5aNugIE1hA+uYyX9Be/kZPy
+QqHEWNDLFZQOIOiyU/MNc4XOSN7YxUE9xBvRVjKHSDe/23gUVara/FtAhwX15/LJMdgkWzgZAHR
JdQVK1Fs/7cteGdjQozYGgvrDuZHjvtK3kxpA9odvNT3PgNTxN+trIOBAb09Jnu0fFBpSKTIajZK
26VTIQwxiuwX1IM4StnM0s1UigtHbAMESlmU95UEvcgpd+OvP6c3Tr6XxNfSQvF+CdW25Io0iT21
zHFLcN0ef64U0we+KR9h8uqLFMKtOuFYWsD6ON/4l2/arOvC5rpbhd/5ST9wAmFOCqUmBW6J8CHk
krHI8Wyrb359HrOdhVjgg4ykk08HymL744zm+NGSu0NXDcF6gtXldvVL+l5NcceO33Qcg6uoDNqc
5pQs3+P7WEpWsdt09fDf4JR7gSzvb6mb/vscrkiZiIq3j8hFWO6hhRuKpQNmlAAafXIPGJ5E0lx/
JXvKsM8HWW1JYOHL2BceAoxNNk1adEY49KWxh0P3z8SynD4wbeuDj6XuAYnjB4Xtgi0cUF6JMujI
GE7mxRaijcdOT48JkmKddvvDz8slMQ8Xex8McWniEY+kHL8+szl/8U3c4GNKTEM/f9PkmOelxbBH
OeUYwu4r+e3sYcEPkHVBTjsobMJK1s2x2C6zN7YjXt1XgMNXuArx1H34b3YAA474a3XDDn4aOLej
2BCwAlFuXzi5JyL+XREqX4f9qGuOjaOrfmAzEW1+qzN7NeO5X83hP/BjV7s4lKKY1iktnNjwtRFH
gCV2KDE/qKUjjejQOASy4ivfmWgSfZYBpvnb4keWvFI3kl2Jgfef99Y29jUD18gs86cqpIbyJIhN
jf+kp3btCch4zhtMxw8uZ5maLW/ETYiq09xJAwGNAwD+3IVBsvfb5AsdvAoMZG7oKNA/lhj4N02l
3y7St15a8S6kq1UBtGrZK+D2X4eZ6Ego74F00L5y4P+2vpoYbQzMxbJqPgtBtXrfh09zoKAI7Y59
tXjNt5++Iwgy7DDukCVKYgIsDTwe4dK89LCt6qkDpFurMhMABzmkH6MWo8mNZcU44QSYtmvRX5PE
RNoxPOlGfNUStDuTgVGeicM88XkpB/xQl1dlJBxJyu5moJzcgghxd8JFQUbzYJfHuqHxp68BQGHi
qDLbjkGyg2S4dNagtYdg5tZ9TNdXEWY18Sz+/+n1xqNFI1K8owaoKXze+ZKR+KpKEqkK/4o/ItJV
3fzjRDwDkoU27waJf+pDOtXHpgMmgj4+fCXgPldC4rP9Dqur9Wwbc+bfBkQ+dqc0o5L/YE6K0VbE
0OPZ4mh4AUOHNSiHmGOKDZlAycAfrzCo9GkyhtSkogUKO21oiupkEkFaxGmFW2Dm9NdBDKaEUs1A
uH/cgejzds621aYfo4wjecxeFi3RvAwfKuBnUlGcdN0JIY6rYt5j2hUfxOU/eZ6NJIMhKpH/IjtJ
MQTaZPLLO8KwgdIpLmHlpv0qlNTCmvg+cpAqx3HfzsRQDGJmoStif1yGWPc2pd7FycaDiois0OW1
w7/u+raGveC+ZAvgnkaBrUe0ACg2LxNuQhHBbk7xrF9MUVAOgyFuN4Ae9DIlPX7wAnXl2eYjFgST
82rZK0kkbt3Ua0MHlf3fSsfbP86l4LJhPdaqcvNldnvzAMZSQv0xeLzoFiYDJlkDJMuqMSyNl8ie
Aap1IrmRF6IROYOxwPCVM4v0/H2CcT6qEKx3lvA3Alww/q+Cn9dhQgB4l/y/0Y+2L3wNHdr9+rtO
NL60h3OygfXkFvc9zLKJl4qLAsIh+i9B9fpzPFKGENRBw4Q2ivQyUk0gsze9lcwnUIupWRa6k3IZ
5KvS7dx5ao7diDBSAr/9PMAy2ENOo2xaYx/X7/2QkY13/54MrVUHV0HX4nrtU9hfqI3TZn9Lzb7t
YOq9xO2QMXbU8tR8yxoQAnITYSQ495+cqetqgTOWhjvuHEsJBKjceNKA31mwf5KwAmpmG33cbrnq
uJSMelSqr0Fv/CcEESJrX994cdD27JAOcV+etlzbnxtxCylJ1sgq08avUg99fbmggJu6BWLGqnbR
dnNxd5dU9ZTVtnJ+wVhwEhxiKfn6cUEBK0yUjmd+yq6kG6sNWOKV0wIPuLBLLHnsSS/Gt89gqkAa
3aGXoymBT4tB7x4r0TUM+7btSPL65yaP+lqeLDimGBXBr/GNrrBjzsJs7wrNl1cIxvFcRNJyipof
bIvY/IqRFNol3EK57Y98lV6M17Z7EdeRu/egl0JejabZ3XlZMmSGWakfCD505CMkyU4yQZA5EhA5
UDISRhtYvh/NFKrNe6+KeiUoKp4R3MEFUcOoJp9ck5dkhCIidD5+y5g0EuwDtmSt8DSL6Fgq1rN5
bozghnp2ACBb2s/SeS/4SzkAMnRbzItCESOPnbZtjVZ3qzYgCeOxrzTKAS/dH1vSEtWrQNBe6meX
2KU3Wq5beKyAB72HmagC52K7t6sMZ6WX0oDwtX8vl8SqB/Y3QKvKPeA5BI7KNLSAu7vqc4P18f70
PFvUQR3C9SHOZtsdRamzW67gbKUFtnO+A8dcGO4jvULj2UPXhBkEXg4xs8CC2qH7GSQ9FRJlzg8C
x2T+BXnYBca8h+kBkaKRLgnorhMo+OrWDMNcylB8Nh+42fRPl+ZGaQIPV4RtESejlcITH7hNxkw8
4pA/US1/K1tP0EtCt6mF5TbQuULal0lcLAlEGPq2kFGlwHkkDFhjM4v6qFpgZYIn56KTCKaerzrR
GhLGjFiE16wOGOz/dgkY5vJeNhaT41tQleC2ijl478w+NTPP40BaOgXKLwUxRZ9CvuDHtocKfmlj
YPj5HakymRSAeYEBmwAM6DaiKWnHZvCNWV1uJtciXIgrVgf1EPkniLGEgvasBtofT2w7+1ET3/Xp
WIQC2HoVWeFvLvZNiubsOt9h0yU1ukDV3+NDIkHRP1otlU9F4hJskFeA2IPriQYEUFPtdnH9N37u
PISLKUQvouw208wFTy+R6m2G5ZRA38X4VPcGc67yjDXhSAQSNmFBCe0uuvBp/lDj313uGHeXrRXD
6YbYeobz8nDAouSB9CM/c2RjGkUgjyiNaEamYBG0MB2jAe2weEweb3c4aSgyG8kajKV7CDCLouUn
8Nvl0bYvzxo98s+rS0t7PJg+xJl3YWORDOx+iyVi/TZPugg/AOD20gtx4DlFiDPBa8pUuYJ2AWwk
nTmlQq3y5lc7cvKhuVNcdAGVWPRBZY3EfFzgK19hfqGaNLefeAZPDre0RVyL8A+c3TnbSURW8ILk
uSbqhHEbXlsmwwFA9m67ljVMLJ2HP8/4H/23vzW2D3at3uR+m1eeuev0XPojtLvMnqLATn9Cyzog
wBSia2wtoa0NlKoYBNHAwL9o77XvJZzWaFL1DWriThChuionkO6SWtdMm16s0axbIOspTYT7ZDkH
K+vD+GdNf3pYnvz4XjtFlkKJrPgc52z1LJUSZAd86JzOGjKxp0Td+L8kzl7OwkqePeFCUvNQi71+
wWpY6GOpHN/VkoPqX59j3ZrfYuZcpTLgQeY3bKSRnZJaaQlEcHH7I/HeFV6TheheeOlC4Ss4loB8
biLMU6C9wk58ET7dDto08MUZnIlpqxRMWwy8/dqJD3x+VKMBjuUL4FYVt2nnYR3SVAUUSju//ryl
u6GxpTnrkhTuGcGSWnsZ2cs02TLdd1epbmu2dPgnc4z4C3VuEpP4oISTX6efZs7rMj/3bI0ijmF7
Dni4d3ijfXlbeIWWGF+OdS1Zwa2JJTmQDVlrX4pFlFOC8ruyt18gU5V1XR1lLF0l/tpP1XvQFYWK
tQmCNXsajY9iXUufh2S5WIXkeMsjk+H+A4k+Xqigr1hh+epnMgOUDwEEvGU+Q59tGlss950HqHL6
CP3uWYnMr+JHiYaLXkUoCqI/9lof8psGqALrF0tBaKh0b+Sa9qkc4vSAQ2m74ZatsTcLJzCCzewM
muDwzmhGA2fx4YkIm077oZcou40MKgNkOLEESZvrWScGTalRdb0bxkWhzLecpK8vl5S4SpKNLIhg
5pqiTrVPsKYZ/EzHUyrY1pIwzqe1o4tFxLhOIICJPiveuNQNMkOSLb57Xljuxxthkk2n4fwMFkG8
BoqkxugSWr9AcbdhQho01h5RTSHETPVDNMf/pcVPFlFOIfdFr9yyO35QJx8boM4Qsb3ySM3v4U00
2gs3aYkTfKl/zNeLWPJpauHGMHsiPClaEpsaBAu4ApXDz5MikzWoaPP+lAOLI4zElH00qhPgUGI+
HiZLrN7je3QAIRfhMNEoDQx2PeS4eouCPmCVAptAAxMUjp/INWaI3QiTuXqX9/FnijbfFC8TnKzk
r1ssxKnCyoHNVd2V89IiDIrLp5Dr00Gi0kTHti4haeQT1Guv/NDFUznaSVoq69p60ecoc19fzzZe
3hQQWdHV8TMDttaplPPKOoX9no9lQbutasbAlvzwPk5zJBvNxrf9iGx8kvbyzuptZubjk7RObyUy
CtgiSmjDWmcX4ld5NBOfNrpKwJN1VYC84Ypxfa5MaS6myuoPLMp0ftJo3OvxOFnbST7HaqzhmARx
p2oeUosDfCrXIND7t4L67qZDsUHDbRC2B1BauSFp/rh+oYtIYuXfmk4Y8QjCXF0wp3cSA8+PKsic
9vvpWoHfXiVJ4FdIztkoMbmpT33JCDxze1zub+2eHQ3ey6FUYPfM8oInal6HH4A6UqPUrvSkhMVh
B6ztX5UC7EWbvaDlVgZHDuZFW8TEpVz8DCcaQvCfX5DETB+iNqtEASBntdi1GI87n/WGe7LZzk5u
+qmoh5uFSU3EhjfN3KeK1hgA04pIP0r5tybaarY8wEhWsQmIMgcgsSDvp3BfkauBhqcaAkdkx9FM
feHztzlzI5Tur7CwqtbXmHUNz+klRATeY/KWesLvn6ydME94MkLnbZ2L+x/jM74mTOSgeyAy5WW6
fSiMcC98QBim01gXcY7Qpap7Dgu2EzeDlw/dAnivyInmDdx2lZG/USiRi3ipb1gVMpVxUMpc4yZB
MmV7GVPceuME7lOyvwymP+VvGT7OZlHwLiPFtfLdRoYTmxIZ1mB7u2T9tPlFxb//eHEsudgnVwQv
VWJChForsJN/+xw1R+rrkUT1+pgz0yYhyNveJxOB76iNnUz8B6HQ50dnwIjiX8p9kmecpN4EJql5
Mp68UWqMg+AwVlM7DIyRnA1fgbGaDskLCXNoWJrAY8giiOSMRyRKEw/ExF8IgntrmjhQmTTigw5b
q07RsxAnrQFYM+QsfV/hUHjtyc5eXkPhmT19J26K7naulMwMS9WC0h1cB36H/XX5stCTbnMuEJky
mIhM67/yR6F/phXqlO7r7bGt4vKjOX7tIOxHP7HUd1/lIMgoNJ4E6rckgkwe1fJJsX3gaY44MXS3
dR/aKLo2wspibJB7QP12FaiXvxxpEiQfnOinqb0zQOfEK2VgLqlTln0/G02a3egnKW4BffmFm7ei
i1e2IVWuLoRdVfipkJVqRjEuJgGHbVGfvGoXc5Jy5WXYoeimucqYrVfgoSI6Eg+fGKIgvtjzVKFq
26Oc2q8kAsN+47w+bv8V9KpedG/GINtfNMUOjzzBocYf8mnVNcChOeLpepPI7RkCL2cgQv0xTOqI
5HaUCUmpxC+NOChog2sYLDWTF6fvv3f2e4aV4DxUfCKAgyWmGgNrnR/Owe2YzrzCsoHInMklqWyC
aklsJyeZtrXjiXixh+mbeLAu501RS0B0s7SxRZNYv7VOS3h0dqpHnK6hEDyHSZYdcXORoUocWKTJ
S0ci/zdBQXaDWN3umbdHnvnWyx1SvWGz/y+5dN2wLu7AY9R3KI082b5ZV+/VkpyOWn7u9BC1W4ip
RShTs0aTY8TbNGJEmpmGyC/ErT0oIcusYSSywJS2KKiUkN6iUcvg6q8ZKxrKd6ZSp3lg22m8nQ5U
pOuui1hPZ4QNd6PqooORxRE1xAu9Of+ToKpFBQGOUs051oXr/BZ2EXe9WNH8LOgKPocY32HmO/QJ
9qEBh3LalyiLm23pqJFRlfD2bKoBDfeg4hLzmVli3UTFV3Za1m9EkwwmeBG1cmWxvBrm+BUl6O+s
H3rf9Ar1SOFS7LTsIyCWqK7KUVas4Mg51o8hT0g97UZ/aL3DxA8950/TkXMgNwZSBbTZ3ukxTEsx
CbFk8tvwJtDQF7srXCv8zBKH3yh+vX4BENXnmpgNlWJFS78VnOfzUWIpIUHQFFT4NPyyynPqYg2A
Yz7Eb+VLwjv/ZWE3XdgyfQmfVdDPPK7R+aWeGJp2dGStKD6rxZWmniHAdsBNpdt2jprylSfYOruu
+UpBAEsbPF+r7j5JfqAM2kD7uDVh/d5ar942JvlQnCHD+ZhLy31MrpCpIYQg2lThe0dN380QRSdT
PqxmSWse+E8hL/vOczHcu23ZfjSdnQXtnHZwRAOx097ic+0mg9ddNwTVJ44tWsfTxwyi5x3n8jKz
hgJ0Y96vpxvRfFLcOJrbvmTOtZH6hCrM/fCKftw0oUvgNqOt/SzEyljSASE+tWc7iFye0LG9z90z
QhB5FsvwPBs3qRTi3VwK+Ig5GuWF33qK9rOAEoiX6PIO5qicZxDqdUYa86JkaBX1rU/KidvYRrd+
jn6Ho2eM+kE5yV4OeqUstXjp48inyY/3CrBz9x0dbfkixQxIrgYI2G3f+uDnjFgL6R9EyeJ5r1yY
j+i5fuPr68cixPEmF4W1EPdJnaQcUa3NTVdl29gc4ff6EV8JknxVEiHcCPPLXTlxnd8ShfagoAZh
kzsejv3FC/vq7Znob3KEsBP5zXbzaOuktr92lNAVvQDStlrl7f/SMAVx7ueOcZFtza9p6CfE0+XI
8L3fAqNNOd3alDYIsBUF9RlRhao26q6WDjQG0B4+y5jcuYHD47SVxWNvun3YfDcbbmqQu8JDg4Td
V7VOEKuHLwYgKt1ObiaPbxuCyS8/Q+K0nvWhSBtnaOIw4unTb9l1HU+RxSIWEY7CjHJDvsICmktE
Q5Sx3TtgFOo5IkASBXz7y4iG8gI5NSw6xHhEVzTIgtLpmTq7EHVckGEIT8BHfA8Tc4ViX607CXn6
03cQ0zo80+2tiKdtJ6T3gU69nEqZUoM+E86e0f+OEWkEVVqmtqMppmB71pr3ZzTZ9QynfLuAILVY
JWYdsclL/HWApRgCkpieAyE3RNU2j4L34aRA4ZxLeCqdtBV9D/sXCQ3B62rg60eYynHt9i/ib9AP
Y/MZ053iORwfPaejlUKGOwE351GEUVQlDOsXgzuUEtThdo6P9uMs4dySbVxpNRncWsADQtL1/ESy
E9JFRXdIiXZK27qTEgPSefDabDwkQdHvlrn3lM4Bag5ooJ3UeHD5chq06l+QQzyf6z2OKfDIa8NH
d8iAvMzxFe9m3MxCT+ZJs8F91un6hbLT1aREScvQeseKT1gOwm1JzmOHjnb6HfN0OeZ5XfWx5Up3
INinR9p/sNoHhVKZMXhN4SNB8LC3PCqie/hm961qLiI7iPo1tcQ7NBL2ilI+1m4TCLDQi/xE8rc0
vS4XVnoBdoaITcTldNi3QNwuyAhEpiXOIi5v9RBwSHxjZ3mut0RQ9DksK6PtoabGzAG7LnLVoGNi
nR9JPeNNDVre2uW5BsBfCFRroOakyyZ2iHTyNQwTCns/72ApxUtBF3satg7/phSXZEBqV03PwwGX
yZVruucW0w/6rA2ni9W3Mpa61GHPDCMLvvI/NC0tvP4r3zxAekSqod3obXrnzFhxzm1NFvXd+R0O
YMpTAi6Z33XcRAh507jiG8MA2O2DPBtyPMfnRG0mNxIE5jwR6d9ExiPU7yoodRuU6OS0F0067Rwg
j2BnvJnwV5xrNFaEQ0Tb02XrnGqNY8/12K9roWr4wQF1qqmnAshKTvPxGrhkQN9+Js5WL8ADDZWh
2JWH3DF41NZjpSrT/cMWxj2nD0FPot/Bda6jwmSXc+izj8Gp4YQUxSvtBX65TVc81nEk/u5N3mnw
uAgRkKVbcgHLis62HSOGZvMBQLSpvWJ1LoHAPON/n9+XANEVyFeRstWd0p+fmCjwvmBI8fPMKCEx
W2jf0t7O2pQUcmYDqyYgT9L5BKt8jRlx/khy7RiVc1WZfMehHgBtsgSc+G7LomjjCFBfyzk2SQ7w
RmZSvXtUKGhOVppNw0A3sWaQoEDkqQevjyRCKaPg/qCfJwPMeguZBjelPYzr3ZhpJcsGgvahAPqr
aC+6/fxepr6ya6lxV4Fl/TfZMxV70V8YSJcBbue5dFmW6wCavC0MKeIkkoR4bVz1kESUoJPqTwZR
h47fTs8k5TAxN/X0OnKDKhm/kkEnYIld3gsmDHzPTI1AfyS1REWbQfm7qt3FvY4iWjyxq9RK8Vt/
jMxicwK+n+v7GldbJywMBdTZIqc1X+JNEbHu1enEE6embyqfO5Jl7QFLDejqJ91AwfpjRtcJE5I2
omoJH3xvQ43HRREnQj9OsQnb6Ir7YmcO4ej4z+qIDxInAcO+/oqoYHuTZWjUT9kCjE0hvoLjio8O
Ix/ijVFC9FX12Xn23Wnii4oi6SUQ/SmYC+VcdL2WKQkI0X4vZLwTFiWpJDXHnJK537JdXv4Hu178
6Z97QLaFxLJ1jnkXQQ9uKTuauqZnmDHwQVCsT0R0EKuQpKyAPLzpfkmsEPpj5drq20eF/iXrp1sF
VymQ5p5NVnGaPWYIaNmzYlA9bdXzNDroggXkisbj6zB+CvfiO07YBESCfOm6sxvoffsNCuq2Oudc
5OhDtUxeAKCWmuKBLvAdIaJ+P77FJ3QuTbZqL+yKpW1moTDnLOfWJ5BAw6KX/78MNcTVFbW/FwsY
M+8Mkbw79bGOx/FF7HgYX2tgRoa0bpv/Zjvs6esixJnFacJ6pf+scRNmsrvQK+4+f6V4cnvjj1Q8
30cYKdjP74+T8TJnHP5SelbXlEHdto7brQvVRq6FvipFJw0+CKUUYc6vPB0jLKmZ0lBk8Ki1zOBH
ocy+FcvINo71UxQGEmKUzmJRRdhFmegzF5JkszOwjTXAlrpzmjjIfkg7U9snJErX4cx3nlO9euLW
wkEO/o3RV9UTHCL5aOAgY1K7apWUmIkPLBcIEqno8fLBhXhFXf+W7heCWVWlZm/i0lE3rfsVgCq+
kIH825dgpQHQLlL4vUq251IiwPL5iUihtmG7yM0f/dEvWWXUx0yeC9v8eY2uSLfXMM12/NcIEi87
S6mPVwrTOrfE13DpjmZwbEZ0rosAIdxU6zdxohIotm4Rz6wLe+I/oUvXgR2H5x17PuxKD5+q6ldp
uXJWKSvgzh7OHwVh6T9jv/q+CjmnzGVAAyBu9D6Fch69YHKj3eS6M+N1Ftj6zWYqzndS1VGPImPq
0QwC8K2xTKU7KZLgRW5OKdn2/1QRcdZAzjidiT1U6N5m3TlJeU5m8Indh0sTzp0Raiw/pyPPpngi
NINgdvcyv72lDlqUoju6fygZ2i7DpPr8eOpGqBWX9yB4siUOfXVhgxkf2EiWcXjx1NBPBa5y+bDT
yk7edZ7OV13lPl+qm02Ll2H719MjiMV+72qJcGjD2UjtiWNUxkY4DOBe+KRRPqC/80RdZ/lUujK5
g9/Qqz3OT4o5nNJHyR72YD+O3/qMp/mlC1CwK9avVRJipAq9w8jOS4HuygJ0yCA8GARdplHp3CC+
Nsux6Dvu0+yuIp4CjBWQM7xiCDjblUhm83q1FvKvhhXih4AisHOWHfr5kv4n7EfR6NVWtdXJb8b5
ALJMmVXjyJHzQX6+yL1/m6r53XRo5MSrZeBaxi8ifISzf9xNdXH7IOUxIDV7fNdfW1wfM9DE64t9
mrVslJu8H1b1rGq+amtLSZE7RwElesi61YCZv1mTndnC+bqq3yKYaTUnctPpBD0bkbolMALGJbyT
XqDFc3X9JATiy80bFF+9+YQmP1JhOyDUXK7+wLnV2iym98L1+qE/Qx9+aaX13ac2NqFImzqoThFf
qYxuScpSon+s2a9UMwz2JYuddi+rRshLFfLkaj1NrYUWGHFRJG3WQPCXV2vDpm/9d4kVxQC7Yo4a
/YjGk6llV4NYdz2R6EfNIZwaqER8EU3e1zpbLpSxEq+aKVK83TGiHswvcy5BelVYV5b+4ooKdQtw
7Ph33lT9or8ucAz72iHQsguzjJ27hX1KdQlc52I9cxDnPfSgEbHRI0/W10WLbXyzVl4EF7zWC/m+
J8SSeh4YXMdbtKkQpu7gIgCDnxwNcUrCm3R3fecnSLpu5DUCj60vRIuKu+mYKdUBTIfSus3piU4G
gsfMhD4C2GkMaA6FCgWwnOr/HWaSR+kl40/sDkbmj2RFjGmbt/A+T208e03PCncYw09WU/p10uiw
aRfzFflta8mz02b4H8LTVjzyJDVaEer0JWuvomWxCDbfv81tT8B2KiMVqPUn5PX4oYAE1g8czJs6
7g7PxKdPzJTgYViVXdhBqAeggL3837M+F9vbeosBzfetwpf6ZvYXjV5TZBLc7vPmkQVCjcY/UE19
KZVhLd0LUMvTNrM5rwQqtWwQDcQfV9Yawoaxee81PThdgNypjh9Fl4nyMkrkSH0SsEZYEtGfB+ww
EwLTC6hFtc1Q4RLKPmP8GfobFK3v6bnhlJ4l42wWIOnEn3LP5zJK1e/ETw39lKEZvMgPzLgYRVq1
8hfFfzNVjSJ79UAdmDv0VGfoJVkMD1vN+idq+C3SgQlREXRygM7mFSao0gd+B1J26tgTqFm3lm70
U297Gyar43nfW5fANoO3TevaTCN36WTaJ8FB1za2pW9DyNWkwIITyFlmOAGmZPKeci4UlxXemB+E
eCCOe5hqwmvyQshaBJhzC7KTkbF5S+O6hbWn/Lfy2bteHFpKfbI4shWg2g2hHAd4TWYPuQDhmOCJ
bJsZQ7MXeWMu/oLYrjEiVrT3ioIOke2X3rOqqeFvCsIg8P4yQelpx1YXLEyC2Qnod4F88H1qtduB
r3ZnbCQ6J20qse1iwEGzjJQjdhZHJckt9fs1EfapuUHLUgdrmzXyeqbwZGv/yKpugy22VKB/X9H5
AJcm5TQNvGBfOXgiOFg2tx5r15A6SF/22LMvT08cj07s0lKcFARR0Ggsoyx4mWKyExtBf2EgbzWa
9zwOzwLuzqOBPRAUaXfhFNxxB3PwH1n6m9fQkw+F67/lev3UN2/xfVSQnEug8Qqbri6JbM4M09Js
ID1p8H3iKXaUu0RyuhKdw0tolqtnnbZxjEmgKnVI35feTRh9pFJjHFp89S0F6Xf1jOne0RF7X3Lh
eZtvSqZ07DqQwqjWawD4p9Gb/1xD4Ho/FWdNeCq/UzIdyWDblrH9uJAPL7Lln+aUvew3RixraK3h
EtBYZVEWRTzfhIWC4bYG69gg/R5HhH6xWQBJXE5Z+SRHlmf9OJRQrgwdGps33IcymIMZ2VSIInHu
Dw7jHHSbJ5mZzdpeS9YAR4tPIyzPyB2jV0WfSexqGRuACwUPzWHQAaeNMgaLlCuFK+5FrH9hi9zA
qVIwRvMHNV3Lye1j74NC3FyPw5gBG8KFYcUFJcvCGR8zcEi+ouggLwbYfZVOXGm54UCKs3m5zn2B
IFHDH87ZSrd9EkgnTLcv+o0uKtBAKTWvn6bOPtIBPOAyrjcC4XMCjvx/RppPAKq6ECSVsCQwVyWp
/or3NQIxvgaNCy8nzioEBVeYagbwAPuI4I3BUqp/9H3f23L4xqwRZ0ILEqAq0lfZd9QR6qMtCsHy
P8VfA+APtA/uMNWyxES/Xllq3AY4RTDLu+/5uVk94NkLxsN6JcedvxIDIAbDzgsRqh2o9sxpzVEl
JrHPw5tj5AqiMnU6qDNiFee0MGOiUYwIRC5NSSilGgt9a407sGv6SJUt+xdo4PFjukl5xADZHYfx
VGHoqOyyW0fHsYJ9TGo3hPIoxPypM4Xk5JOepnrr9TihUtYpbqM0H5bGR1XgUyO/niowJ3yREAvx
KxQ9ekPi8N/wG717E/htJsiMlDKBElwxv8rUUGvY2dKv/UNWzxl7ayWtcj2i0VhYSPVjbKXZ2x+j
9lbeNuP+FzKVOR7J8dLRZSKR8WOs5s7J9sZecMQpT9j1aZNgFA3HGQLgTHxEmeXBuULq4YRM96r/
qcgngwzZKT6avS70pIc7bYbWQXY+h4rW7PC7vK3d7e+3tPRRxU50SR/HpSXEbtCE62Gp71zCykN2
HeleYteJgRCv19fSRcpmIZyxvnzh++fjSJl62F06+YB3ijbrc3L/Rphd4lDU505/wbxrznw52eO7
FQYgwaZFGM14pSwhNi7A8TnM1d3CAgEkPEtrLFsaiq+Jf49cTejn9WZkMDGiyqLObwQvx+YbGnSs
0bhEp7H8XmcOHuyT/+sIpKPc4DMJq3HLJ0tV2NtZPCQLpIqzOZwKrbsk0DAXMT0/onuZXeRlqIVe
BP+Xq5sZ+zdZLMzHzjOdTBL1+l+56CIJX28x+DFNiC1gje3E8uPmymZTaoFASDkTTlu7iQNrWa9W
oNbwHmf2Y3oMnXdPS8flz7suqIUruahnlrIZXuqDpGe0YMcvTSojIM2oeSVHo+AAI04oKwLYX5gP
7VkgZQ/FGTEP63K6G+L+IqPfwN7UryLYqRqss6s6mPcx/6PLLhiJmhMmElyCSfdIqURNsS19A3Eu
EFyWMHC0aXkGyNTGogHuu5at0Axka/IVrLk4tUMjs/SmRpTDxva+rO9zK1OY5JO1VQOYjpHispHj
iJb7fqNr4zJSTibcr4QJ0+tjysAnveJwbRSKwrrOvPx8pcIYRAVpyxbrWHAVuOllh00b0WYWYmy4
K70J62rwlqWNdn5gcN2in6Dt3+8FbLHLG91iTosBkCwJuN56IuAGOky2Q6/FG7HQCLTpjfXQTx9d
ExHaT8JsQepNM07cAJOCwEX4xbpzS4gV4jxSmW64Xc5Q/9hehTazQgshf6NMgatjDvuKw7bw66P6
DDE7IYZv+zeXhjgLWcnastxGLuqdCXhxzKimZ7DzD5ATECOSJ78gW/heoVsNfuDqfFvEQgavS92I
aGaYKxy81zLnqnSzj2Hy8V4Tzrx3jmfgg55BxiTqANBJS0P0Bwsg4ZiJvbP9mmdaVobit07o/2g2
kzQWBaqlHaTYw5KslZPKllmjWAbgr89chpIrcYODi2ZMNyUt27CEGkclep/nw+Id5YkSgjl18OMb
zmrId1e1irXqP5XUHmJlat4T2MUJDwrWRDREsDZq/IPWN3S+ADDQ0f/YOT+zfM+GC5OZd8UPz2Sh
E+inohg8yWVyyntLDyotS0HGxRT0vRYaLFm9pTlf5CBYmHp0g36A3vATRRsoZaDQRoBVK/lM7dza
OxylGXyh8NW4KSobZg3LZ9vMCKq6Oq7uBZyr19JPfwHcgI32SYsJgysbQ5ax3XSifnm+eLLqlDHj
innAgIF7b0KBBXKWSTG4CGM6cL+JvnJ4hIzk13eHIRlSnXGlHt5yVKoTV6EMtl9GUK/bPkR0P6sm
Zg5E304wELakEY+q6RkJKFhy37f2NkBFF8N6/rsvvTxi4kf/E0cKLE/esheQX1LcgFAWi+AWbUje
WBKfM/fymDo33JFbeat+L8uDcRzlgxbl3ErI9a10mlf2NY/hhfmijIE3SMaDBaXWmAptckhDWx1S
dq75eehhCnXg3oSlY8jQ7alM+ZFVpryZ6hSZ7E4zzvJWVdQ/26TqnYg2zHO6RuVu+MrC9aboAVRL
LRImE8Tco0TnqqGkyTwf3kSGvwpvQnt9ohdMpAuvQHuZ6jL3//H/Gas5a+6ytc9hdWhJASa4JmZj
h9/si2PV2GQdDkJAiuhCIZLynLkXB5rgdRJ7MArT9n+44/OUzF8TgbOSnW6Re37TQlhl4TDxcGeX
xYUD5feCB4GWVEONQ8cPVR9GRYbRyOVRkz9gZ1gRCDywi2zJygmmo/rZnjR5KiiqnZhbgZqtssiI
KDP3S9VvxH4NDcJqNQy5HSzZsYXJRBUzt8zA8uRIZCwG/SwJMcn1LnXYdyr/JfyTrTQpeNaxq+ov
68JXkmq4KB5id6vs6HPc51jZLynM1EnWstcwJevF/H/HqNxw/4PFfV0/7PENMIlULvcNehFimDxH
s/FdnkYdg7/s+sQspzZrLLtOStoUyj4ws5ezKWmLflW4qLW//l2kWpHwDr2c+LVbKrK4f8J38BfE
aPiUsT/8ORRVl641ir03lLntt6SS5984axrzKQtMFYSDh5s1hdi8T5Xn6rPB39/X41DCj4Ubqa0T
RPFOC1RTIwaoY1AQH3OWppTjtzVXZo2RSWQJ4cJE5zLEuQjP8IV2+f2E1Ebpdkkhki+solYKXfR1
D/W52SAuH9pOxjM6MVQ2bUt+By3PZXn+dscZ40bgG87LTiGNCXexNN29YEu43cTDKNP6A7BKsVoe
eh7ElrffTAORWBF9miBumcjkQzmu4tKirL3ZhkCc/itmtLbL+NFm1TfgBYn1YqQiSs7bLTrggQzX
VnRaK6eltJoTn9Le23McvNbIAMjDfXEujHMvKbWRGfzCG944h11+QvTuwEEX9vy6Fia3pgcBtv3W
MP0JMnbQu5RHNRxarExtG/QmTeZ6oCp2Ntx1Vspsi8QRdWmMdS4MRvNLCyZdWZTolE8x4fq+n+4G
e3eP5a8TaVFguozFJFxtYNYuYsUw3Pjvcndy+4oHNHCywHcsFP1jmTO+tiIczpF/agKHFbCU1Uch
6VWIBuw5cEmT9SCLjvsTSTb82abT2jBFITVW/oHBhsCroDDGYt6qTITtn/rZ78Zq40xTYO5FCRFv
7IfOFgiU6RJt0xC0BuN5d4H28NhMfx4h9fPZ8XUYgUMIbPhlsM82JdXaPT7kpn1uAwHUm1ajNp+n
I872Ifgagx4d8x5S4q4tAH7vC0xF2ke0q2OoAdKMYCRbX7S+Eck9uODG2uL0SuXuH1asVzq/Rt05
OEvF1V8tm05Ic93t6zRbkkjV3l05MUZ+bTGVqJa+VaNtbqtLqubkvy0oSypQ4szL4rYgFwdqofFr
NOs6dT8S1epVNr0yS13t24//5ywfAYPy/bKdxwBTXoaIMjjhDv4h/X96Wp84rm51JvOT4K1ux3gB
g3zAw2JFkgAWPTXIoPxbJ5ZeRQSNjTfBM6q7LFuleIuqcS5oK5Z2VfCxt65GKVhBH5imOpVJFeNs
5byKRhf3vJbZb0tejg2eSxwEC4L0z43hY5UfdgIv0qp7A+tSimQUgWLUcUepkOqNd/2i7Ilj7aft
GDj4SZFCd2xvoBsC1mCwghJb4Gm0vPfaMZCJzTJhNG0HzLViICQb4SVhoaYAsBj4bGIswj7/VU6N
CF1OJR749/d3o8VK7rkXqgxUT5/oW1tDFA7z4qzZDh9TFusWSshjOh/YAfoiulohCcHId6gW1CjL
US4+032TXWNVV7pyDU2Yzbj8wFzqASuVs3i4h6Slh7diFqL1URcV5SiYmSKakBv68YX/ZqfnEETE
bITyfe3RlK/odAb1Vr0KUQUqmPD2vcHPJL27NHWLfI0t9ToiLHZVzvXbZyMBFMujUZH7wCEmiU7J
YIGn8VLwt1yqfR4Pl8Oz1z+5jeP0sFgAhdzAHDH+g4J8maJK3R+H9B7DlxljpYIrDc2cxMbouxzW
5L9p2HTfFV5Pq7fBVI1EKJZGGyjDYURtYoXF2fbDYYO7RqnzSYdt3oGVaYaguk5siVnKprdKr6sI
GX7hTbI9+TRJPfgPMoc/85PM5PVX6lEckfjq6YZNZEccQFc2m6WAXUCXQD5kJmfM9VeVdnombWIq
9kieP2nBN9PMCrR1xwxOBk7E9A1fYtbtqqo5paoHRdl65fOB6QAz5ELXsAFcxbor//q/lvxyygKE
Et3W3gJjS6zK3Q9EchTFq8qNTYOEacVxtccO1+3ll0Uz7LNgWhxEK6GM+Xsyupfd2Zb1g4gFiJOb
vwTCnL9DWW8sxLV7Y80ghRoLYQSCiaRwsR2PGUIANEduIDMpD13vx/yeIu9y6RG++71Bf3+4Wsnl
eFgjRV+u4Q3hUMuUZAWdMORQ3jPVLskq26RiZdKsTaGATQj8F1TMJ97hHP8jIMeiETtICVxpJgRj
iHww//m/TQawiKoeU03/UmWEp3W61euwAC6VkcnDgRktE0ivRlTNh00fNKUbn1OspRZYx3tT2Umh
Ahxc58zW9ZsC+HVNix4vjWncM29QG3fBmPdPDdtxvl0NzOOpzaT7tZySnWOS0RMzVXpZRM5Xopek
V0F/jJXRu7yLurbUeLKWLk0G6GDtlQOpvvcduWsnpTrvCUmWmTBFMGmeLz6b5GJzS0dvlZlt4U/F
9toeSijhs5EbMHl8wSjE4XtM0sQppjFUTU5DeYhssN0jIViyi2QcDj/WZq+W4R6M1/vZiB7qg9wG
NqJglQB69z0kL6Uts8uVlCXOMSd+y1m0U4DEwTCZyAdy1k3VMqguxbAdzrZ40aV+APGSKOOr1C3u
VNIz5rZ+gE8qVxPDNBIycwGnHhPIF3EluIDKA+y3XfgXzMFCuq3xmJriPbjsa9pQayEwhkMiPq0N
NTEXM3P2FZG5GyLoKsOryjCzsK1Kg49opMyPFeoEWcCDe76Ucl0IyeWW67IqfeHbjRbsnkC4MfyI
B9qCySlLzrf1wvGG4KRWwL8l6j6MPMegVa4EJooCOmZsu0uKzk3Sj0Kwpxvbw5Zc8qENpFhKUwY9
TW5vrAMAmfyTmZBrgYs9504P7+KJpJ+UMZIl+KHfHf2CJMGQkir55/uXLpi1v7mlMzWvIK6FbeDM
qSxdTt9+taod3Fi7Asm5LqIJW1fZHwR6oo/bfSvvvv0/6K6KlwASa/Sqj8jTzxM3sXkPsyUNlXKj
+/uAsyO8bLJB2fQ/iTW/rcWixMOGl5DP60qZtatlu+hGs4urfM2MRYjGXdfPy3xzvW19K/4QZA4V
WEkzGxHmehIhPYldAQ8IDjLmUR8QuOuy3B59+1h7BRYGDUJehbmZQ9TY3hcvwNWWf01E9GZ7F1v9
s9too8Iu9syLdXGoNiGd199/lDXxDMCgVlG5wckXGmN+fk/gWwZnDygcAwM5EW19BVIAXPuU3OGs
O5ze1bnQewb1ckRk50K/sKlcc+9MBtTPrA73S7pCaFPZpSzvsGl9XdQt9h17Heqzo+qt2z5sk0kK
M3G9MA5CmP6ZyETNdyLrC//CyjdkrUo+qONV9uzdyqrZLyRbLOFKqaYYLARoI1dYfqDBVQl4i8q6
jBEMEV6knr9TcmuxJeKqXMAZ6Q52mIASfGdPSKYCF7hrM1Dht6JOtkuU4w1CTEiRytZBId1g3CoA
q7d6to7kmma73rZ0fv+usC2d7H96CKQONKlpdEg9t0cEZVuaedfowrMVmSMwjeDXFpeAbC1cAe1o
QOuwXHPnyXuxrfaTcbxN01MTQeSJNRSu2wfUVeqqAoj/NZIC0P1OaWlMm+4yOxndxrBR6M+WjV4K
00yqEfVsns3LoMqJdZXHqZ4LCOwryKlgKL1UjjC7mOEsKAcTwwyXzvh32h0CfjV02LGhyRWmlMr8
o2Qtb0c9s2kiCs61+zLM93ekrzJ8b+st0Pwn+/STZMhrjbO1Kpk0uUzawcO+HygENmxroNWryONm
ThECWLiUvm/npYog4zydcv/8tsszgkxEz2CAR4J8p4pzuORgpkQ0vT6a0Icvf2F43Glgr2aH2Tu1
pON7LlTaQ5Y/L/wHDON0tAm4/hYI3qw/zWCyGSZD3LKo2TuikyJS1JN44Ipa8Qx5I3cIU90VIh/7
tkHUgjLo0xQSBh5raarCd+HeIAGebhd6LS/0lod/OHGoau+7S8T/YbrZK5tU5kNwgj4Fkom7NLDv
GIoAnqlKxcIna+a8ZKRZbqrznkgll55ZfLX/lR/GdQTIKS5Phi6qSN3Kemh/IyXyTBrzOJJqipKL
Fc3+bxW9ees6lK3aESbDVE7R7r9KVZni5aLnXULWd2dgbQz8WQppSS4btiL3bEF4C/XHNKhio4rc
/QHRH9jorScbCjXlzKd/GobeeFNfJ4x9M3nds8WmEN+v5531GSOEdsbNvRP3eD1Fq+9eYsSx866J
gRY8TN9FyRvD7Hf3FbJTf/1oYVylXpwGhSVUTG8Tpp2tcsCnr3mqHBKva10DH1h7QdyHIchLvB4X
3V5tKu29t9fgnIGhosGSLdjjQCZk5GF/4GcKr+8FQ0Sk27U8lfSasQfoQklbsO4ez9C8YO7OCGok
Xml/V1B4/lUOn5jISnM2EsII8bQ4Oj9uzNtZHIIMwCgxlHOoyP6QC01TGw7BcYoqZx7ChMc+895U
iLv9SFcV+gzo+qCrsUzG5xmln1zMEFBuI8hNgMOfChnUOvEptZyfIYlpyHp1gysUGDQhT+DPASIz
UrXe5OloMyUMY4GqIs58jAk8R1nsrRGGtBnbpgG9lCavVWrD2boRfIv3HIHRkYhy3b8dW89e9mtZ
traLgvOH9QI2z/2vumWJHiZAVkEgkBogX4IoHKYiAEu2aDcHtOBcef5AqOq8BCiod+YAMlPCiFmV
3i9hPIJW/vKQ5ZgffJGTY4m+A2aoJ4lWNDh33K6EzpeJ3hswTsoNa3siEeeNIZpuii/n637YSCQS
SowZ5rjQy1XX9JF9l5n9hJZwVRjoIIyEAyIc4BPNj9J/WvvYyOis+Z3btob5xGp07R1ecpVqj6t9
wvF7HgoEp4DAVS0dH+a6w+DP0VS/+3K9i6s/rYH/kjhjNtMz+WnoHF9+7UHtaTDc8FnMJz8A0GDQ
XPC8BwlgUOm3EmN81tr2qfm/8YZ9Kb4JfQ/xN70owvAw5GsKW/B7FrlkrjcEud9ENvg35QErtJEb
pKvF+/ZUc2/kv4OdUuQ9USstJXcAr//LN6KlcJPgO8CcPe1fmyzqn/73dN8imGxLhkVVMleoBWDb
ExRU5DiNlhkevDpxzqg5C7CJhKCbn5PEpROFM6SbRMyfS+JA/EHeQWASIjFU9rqub0CAkuzypATP
ycwOBEEyGdjpnjK6K7vo1E/DrsVF35W8i3Yzv2QnZiJqbaQSayBcBviUG/Y573ZJ0IzK0UpmQU7p
dlKRA0JZ2wFPybAhfrxIY+1mp6B6iNjbfGfB8BC4ySdXhvTRWfwrQ3wXBoXLnmsAxZZKeJSKIe97
R0rWAJSKG2Q/pMLtAsvr55tVIQClJEy54YKFG4EVj2QxyeuoFC8g5v071IOzU56wvpYgRVtOke4r
TYxk7FopqkjPjzptOXa8DAfLQVouPs8QcW1q1nbbB5q+2XXXwoo1BLZ7pMzxiHKEdCwUtSWqKF/a
gWrREaFwXBewPQvmxP8W3I0XLEYkyzg85NYUCx/2RbfqW0BR4sNSUT3DX0zqRoj9vxx1bEHSrILe
2cySaza2BBylb7Lo7vxzOaxxUNWPsoipv+FyMTAsK9mcXpwNtd+jEF/lsYBUMdhsUvhdvTHD6Zei
ufoTOqOnGe2foC70Jj2Yc7kbqWddCuRiCdDEyuDIMYv2rvnhtUnbFEQvrTPPK63ouWwghZMtbI/V
HxhIu6BxSjMTg0GevmZJnbGUJnMSlIbsdnifRrutEwg2yWGJgptRruMaJVHkQq/kdXGOp1tJ47IZ
TxcEI722kcPbePmBewT2jddRz+QjlW5MA5N/82YxS1ggOWXX7jwWAHUPTptgtkzEM6msFP1ENovy
FSc7YqhXumakgvDqeC24Ryr9CnZpey3Kasdn9vG324btb5sAIrPZiFfBFjtUFVaDK+dQcnb7vXvs
zY1BQ0ssQDesjjT5Xsq29ZUhr3uWHX1KZxMjM1oMew1EBvFyucyCIkA8bkvhFUokBD6lj1/Fw7Gs
Ptmnz1kq4deAmKWrhA3DxP3Pl5w55T55hW39C2GKHRe33YIDno+iXBJyNt8HNxVuBfPmL/B9K/zt
90k6bi4ezaNOTpFD43usqonwAZ5K93dYqHiyqsDWACL7H/mdHVGJsTjwpx5IoXnmulxSRh5sWLSf
YyLymhEwYeXru+LedcPSsE5dywmWwYo+esQoc4m4J89HaKjEf9AVtExaPe3d4q1n7wbEvZxY6y0c
BSHIMSw23TCehM5ya9yxyZFKrGaaxAXzCa6F9heXGflLEl1hqamWs5a8+g6bRuZO9FB9io8BJydB
BS6ym2ypBATiBNRYTOiqgAhDg1fBRi262SuuvRRs/uH7DXa3Y5pRk5COjjLEvzJI4nILkR7abwUv
qtIXYf120O1UE1wZCZRhUEGPeg/1vKftc3yLRc424d3hTzolRYSVAjKrJDrTntwvjd33yAVmQG2A
8IQJVhgEmqPD4KiItWOCL3oa7nPzgP8UuBi026XB0SalvtHbGuFFoBcyTwcSy/qNlfOC7OZ2VMl7
HapBuk4LRaOoS9fQGHgxHJSr6iWhhh5p3aWSZVUQFWoQkgc6v8BqsRLeTlV1Tcf04BFh8Y154WE9
p6ui9YPYy+0drqUlcQZMlCA2PdNAHOf4/bcDm8lbzFrUAKgWETfS3MRuVTWiEKAmYvyQIhJZpBJq
VgEIbeAsO+tsIeSITU+/ZAnjl4SvP5yguQC/0HEIsKMQZZgK0zgZKWZuqrbia4j1J7uSbsw8XGDu
fjIYTVehBHZvtQd6opZfZxf+uzDhHKP3IbOXJt2vEKWp9HhRitJyM7L7eL4+OtGTIusSim4OWxVR
Ke6hDHHQCWqfc3anRINhhcLxXH6JRbHvgJfoL0PsPzKBnN0iwisd/4vbsLd8PKPXpUtbWVcJONaM
cFaWiguXGWW9DatMr9rJnWcrwnkGWtqvWfj6++ZpE/Kqh6d3kLrJYnKeJtT8xnCuBw9AdeWq+Ymb
GXwuxGRHou18zTVUcxoyL1DNuNqK2Qj+eYZAZAQwTtG5V24A8Ogvz3Buvm/nBMxB6eaf/28hu757
GqKKN5ocBc9jDBxPr4bO9oESrkAHvcFtASNPLGiIhsOWsNHdmwHwDM2U29YRWLMpSVv1oYzQTX8W
D5fnkKq1Vjnn43Me/HMz7jqc0xk5G3P1Dup2MM63oTy+0sjXgUhYwAg/t7GeQ3hTtnc7pOSNDT/t
SuuOYVTUZR+e37Ko82LGEKitZ+l2HhPx0QnrmroAuDUK49HV7x++OjGHBkc7901LdH6NA6oTXaVX
dQISPURYnx0fj7rx8HEK9BvmYpllJNIbMm+TyWGcwodeuB+s98qwTVBsbQPbksaIrynBcP+7LzH2
wiA3YX5MsYwowS4qu925oA7nRbKL8qEO5J8/+V5Og8IAm8lbOz1crST0F6SSnffXau8JsqvfNGiG
8pFvqPMj44ZdM5xmmzdLAnJmoL8jyCxEt9kayEPi3dPM7r8nnlRz1LMRNqLTHItp1cFXftyGRgv7
uKnSi7E6cJaf4D7ev23WTGXL23ha/W/6V4LB8wFVCp46Yvqa6Qnn/Vc5yeu1/lZ5mxsTcLrhlin/
hCZ2gt/Rh6R6KaTQUoYfyee8l8C62vf9cRjOqLTmVUTk9A/RWMfyg1yDbnIlMfNKdfZqYrbwaYfd
OVQHc9cLFL34xtK66SS0F7XFo+IYgWeBD8XDKNHUu++mJQguhq8WwGCIDoiV3mAL096EW4Aoxhch
chBS2L9gekxQ4rmiutXjYPBzi3GQv9wSTUg26ZRm2yn6MuFMB2JyBNDHs3Tpb3dtrgz5zGlHzpVb
5SWLxRd5/IBjbs3bLFvLRlKiX8pcVlKszH1sVAzreu7mhDv/gnP1NfUBJUwH8+I9+mjKUPvWZpJo
PPElumxB8PSfkyH5V0xTvOAzqWzNo4btmAgA05cfHrNZZWLMYN4hXXTbSycsDpqwFeWlWPmcblVh
SoMIJxSdL9b4+BQq58ZUKHBnOo9408T5anihw9CdjYBBKccF6LbJPFrxG9k/omJh/ow95/NUIgFY
2XS833ajOzFIo9f4EZR5rHH1q17a9e+45ATtuoHfOMbjYVdDPeOKtwjdtLt2PPEJB/3veoKYSkPt
Gw43058IbECWCD/ESMohYV6QIA8uQCPiMnFAWkMtdxMMtsa9zBGhQwbqsBsFeOpzv3v2iky8P79D
h7EWToQgOeUEzUrkHOHZwJs7R//BYVQUS1+Y0P2kGN06Rq09+oUQOCuqXYrMyzy1xs6HCzxqHSFk
9o/WiiVRXClPzncX4xIW/j8Wj7HVrphh8upM/Wg8THxl2Hu1ndFxAUVFaouKVgrYcD1BnNgsHgQS
Fb54RD1N1QCss4L5rJVue95ueJg+S5YJ2FUZHrx7hcwDm2T/f6NihmcZkKTc5nukhRyKGVSk8eMn
bf3IEaXLqM3fuw6ty56nJd9Ti1z3jq6XJeQYlMUuWptD6BEJ3E/S8sBSwudXLyleP9NHFT7G1vnm
J+oCoH7TcrlCX9ilGkCMaMVoRCqbkntuXXmbqBjHknMwWiGYvKD5zQX8GBfIRUoYgq+f6/wSVQoi
njFLs5v4RLhJ4h9yUmPYHo43tFGFRlYlh2PxhI3DO8Hct0bKm2ZRvfJkmczgtJn7SbYCwWPT/NtY
TojhP48WrewbH3/n9oMKq+Zyy/2p9OkdycLp1zvimHFkD5oUcXrHusqB7bohsmNZPYdJPOiAEcnq
fFSvqu01S2DWAvSeULPB55WZlER36X4FStr9XK/WjdYMmPpH15zRTTSi0BpQ5dZeMxTWtXdstm/Z
axAsMvygS7+e3BeYtkFkfWEwL7KfAh3LpexGm8QqrHEwzkMh+USvvLSIExcPhNGrIf+1dZGBg0Z0
NnCnYc1PDsOPM+6KNvQd9BJ8bYEaNYv3aCJpqjj5WbRIgCs7QWHLj+CxvKAN837vyaT4A6NK/dTK
ygNIg7rPx4dnDiUQa3f2fMflDydeL/Gm7XpoT7ypJHNcClycVbsDNCjAeHzEuUr2eB2OTufehil7
4LonLgA1JRZIv7Hntl9DOQZh3bZrYw7Tm9F4pwzT+4iYSmrYyx1i/03cjane1dTy0zowi7IIl4kP
SOxZLtdJnrOUM3TQhcpzcQbrgvyyHHOwBCmOFt5DUgTaV0tbaxVjahEIYhh25PeDff4eNAAj7hXa
MmuCl766Xtff3JPIWqNgaWK02/ktS8SDj97EY8HBS8LOMpUhEaSbBQntZY6hQGnm36HETOgeIxH0
WxBR2gwhPAggRwNuN1roffohtDmXL2ZA78Bz35u0ZZjzQWxsIqJIbK0OgnN9ayLmr9OL7WxR7GbC
wxCybBVcS5eL7C9F/qtk/NG3R8K4uROQLv7Ab8FIn5fm3V7+2E2Kdgf+AeHfoMBNYw+R0Ptg2uIN
SEcLb2JET/69fxVPoq1uhYVUFzZkHYGOFLv96df0jQKm68+qbfGCz0AV8I4TJlFn1udgLC3qZ32+
k+3QKyxXVFwFRuO2PVhqtOA2JJExwrnbbM7gAYoNw+QA4zQpAfehRrPPbRyTCQFqzUIz38wI+/pP
7yFiZ6vrXlW+R5KfhLPE8UqAOVk/bQnxTQumWMZpXuuHG6BN8+G2MW9hYNgr4fzFbvJQvijvogWL
X7rI4uC1hGsGqdewIq9YmipAKxrU6VYI3BzYvG10kuOr795wDtJUe8yv41w8PbYv4EEouFU2zUna
pMG5GXAuDFRt6vEkzKVotFLOsRFxoyHMFA+f+k9kBqrHB4qMvJWwJ0s28SPdiaB7DCzKIH4qjM58
6wr0bhnBpjy7XsC4FsNA/KgaOFEnv0UHQYUZGj50OBlFTT4tsV1z2FBMyDcnvaNtGPgiOzDuTtTY
tFDCUnN6jm+tqI6MgHD0RPtHE/U2CyjkKaMlfK0J+vB4aRIbfPtaX6nSn1hcO504abeRdzumc+Op
fA7Ec6kMWYIqhQmGlhCcpjW4sp0YC8qkttX/ZXe9rqvttKaGU5CxjWXFzJAyS159bxb8uHjJtXvH
+bSLTGdfoObyo8s1WEdKbw94s0qiARPG39UGSJqH8eqypfwG1cooACF24ZKxDlWb4kKDm/6ut18f
noCQmVyog4nxA1IbCQPckp4pU9RUMb4IMf8yo1SvGBMHUpkaXVLu4VWLAn+Acz4NKd8ANnwRpPNN
DGAGdcjnLmGUtdSElnvLa8A2mUaZ5dPQZw5IX3nG6rBWpdFhEifIHcqPr8xlS92+dXnZYWkQO6Ck
WEn9IlTfNtkhf6BIa68VkIsMra64UtGvRVzWL8UkalGPo/UMCZrjkeVJCylmRLFldUrRJA55311k
qoeRekP1uqWDnxWW7UxLAzNejmxZKFEF2wrm+4HrhkgfaU7zTtefIn4kHiv/Eq60dkMUzxILYpCv
ht2TnlcxIq1F8GibYQaYrHsqU4vvbAoiyDE2l8PUeLdlnwsUxD8PIms2WWBkvkLpdy8y4MnEFFHX
TV2sJ7n01PNjNq8q5fEgk5a5yAq+eAT1w/LQamxzQAq+e9OhBXAACHYb+TBVL/wn5SWVVchN/TaV
q+7XZqvpMKE4jKMRZ1+04pXZZd+cdSSq07PoHpdqrojsGgpMNWPHGBKjyuJGCOdNrPNuiwjasVW4
6YM1k9PFtrLHa3+RR6gXPTwhJ8YIjnees/9ScWuGV5wrRdZhXonpFZCrW7rTduIChScq4KHG1g1y
yA2JaIeABx+xRU/yLw1dYm/TI06hjBGOfAewv933ZkdyyY4yppSKwRnmbHHQPVW+KbmZpEMs07vO
u8OeEsi8YGsEtcleGChQ2cynNbyoQwGuco3ZQKtk635B3QVp5YC3D76lielS7bUx87iIW6qJeEre
ik/2E85xtyi3UvWzmLF6zRpSwbXSxbw+FpXEUo77IIeev95jks1jgbYMhqxzQdpNb2EvE7xIZ+Xg
FnUHADskoyBooBOIHq3YlrDck/KyFF3WE2TvJDxMSYF7Sp7D0qJd9KT7SKGIznd1EkPdgHDSc3MV
4fS1d9pbQeDomDhcP8WsSfZKathxipyyqZq2+8G9UCjQGbXSCyPO1BN2S7uJ+ochlBn1Ti4LSLQh
k1NPcnzkK/0lo643t6AqIiTTYRP9UPri8AWrnkhscGuXWvAFwMjZ01n1tOiQDyYM0/Nu/9ng7b6L
j1znNDBw62EAI/7f91vP9PQMo1vfVgeCLPDfiPdlmH4Mwp52dPVPsbVBQd9wjX4sxl6tSCMq5uqR
eNn83zk5MqTmeVFtHLS+9zoNRIHiVu8/NwNHNVJiH/62K2NpgfKseSKHZFjTIHERUT9x7gZpkN8S
KsciBD/x2N8a+QPW3XDmE7LUxumkb2Yao+ZzAxRvbyCH3MrRnp6XJwToNOQE+wn0rbhBcrQarXhv
Ij3rN32UKHxzUZB206Jfw57Tz77XR0edtjw1kAIjf92x5ur7J3AoZ0jkNj2xvAtEQ+yW0d5ecf+E
HKSS6KBfGTOJkBtLFbP7GWHgpTyCyAGb5ekScFJrVvIEHat/VVOp+Ua6u0RBadBkFYdtBmKYryQV
DGjtahJEY/nTjukEMPzKhxS0Q7FaczUQppy/F13DBoZ3HEcHf9AvPFRI50/NlskhzPJh+EFTEds6
0Uzgq+gmZNKtMz/ge8p1LSgl1LzPjar6K55ZnPHTsQ5X5zzJoTjYfh9EM4Fc8MJ4hnKA/Y7Bnq9p
RqkvgbRK1vTafSj9jS/ap+anx8A6J7uQwTG09lmLQVsQQ+KY5AEoEqktl+L1+2QwKdcqP5qNXR7K
pxZdEgBWjOKDPXXU9fyn/5qW4y1QYeeZe/KE0YWBYmRKU5CDlD+YRtYSURugCI1B3EyZRcoG9DlX
fAJ0p+LPVG8bnGWyCp6L5WeYSjEtXZGc1OX39yLKXojrC5/0RZYbvbYJsam+02uShPIkVftQ7DIP
eNAUHSAr0MZtanHcTnG0rKAhMLshvq+W2vKY5xDa3dBTHBsmw8dwqSNKSdoAkhs/JARi0c0BZyqe
fsXOzbvmBHSew6J/7t2pj9Zein57S2uZlrEhf/d9gti42vmoYMro/UUahcW3Q8BoJKhuwqwdepB9
QnduR1b8rvVQuR8pjMyX033sMpV/qAronZfvbaxRUrTTsgbOTha6Geylurkvioup5eGMLqSQvYSI
wFkDLbveP+gW2O3k1AQZ/PVCvsmS1lkE5QKOfUaA4l7ZGTt2KwGjVTukn/10haQ7RVZysuQaEX3p
ySVwWL+wsahDRjRI1809ddTVZv45cimcknWEOOmUng8sNliB5kv7ej5ahRaZspIEMQ9UsSPWaJb6
4mzcKqZuJEfo2gBSH6/kyTC+iUnvQjZqlE7bXIIml8ESYcs/3uHYajcU8wN8o5oCo/b29gywQsqG
PwLIeyLyTGU+ZDhwuoGLt4PAIzcmUa42gBLVdPt/WAFdVUQw5TFNyFd8YY7ESqrk3B7czltksNCW
Vu27jSsGmHtdguZFID0f8IiBp/35tzJ+Neo5QL/Y28DNncCF7z9dQAJMPaNbsr2XgKQSQDSvGl5u
29HatqkkbeWpGZwsrgEYBMzA21wilgwFEzi5hPOz/Geg1hmqH+L71fa17Z9usHYkHoE7aogGxEcD
u+mRAKpa2Gx56hJzyBqHCrE/9WyWVFmEzOAnLb6zBPRN2gxwm3rnXmV/6+5gYVGIQUyRU7p9Y3of
UlkJjcGwgrMZ7DYEtnkcKfOouqzE2b3CDh/3W0Z9y3/jXqt6+F6J0U96oihRu69daTRzYMCOLAEa
qHZHrDwFAyXL6mPX+/5Ntfaqqr8gxzuMrUdNTeeemEHF3VPd68hT5V3e//a3obDMhq9A9cu97ula
W9piehQT1ZbXTEizIsJqvt31EOjbqhucLeOWXB8qpve20I7ma52q7+KZw6fITBNCoThAYKrUXbGb
37Nju0kE5hlu63G3Cex59wD4byFbVQKp0Qxz8FkDc963XeWukTRGdNa5jTGkcV4Y4XsURC68VZLZ
cLSbQIXq4/a1rRHWflvXAI+B3UJpVt827Oyi1izZsCL2aglRppaWe6uYOdGtx6jbUtBeBPygRG8X
Gn5SD8JwFv4u1sA4Ung5p+91ZOOWocE5+F5vxSNOCwGzmNoRdsrZAnmXzUdGywec0FdC6ZTCsAdQ
RqKbKp8CMpZDER8SoHmflkSnKRqFXWqtSKM3LJ3sK4bI/JldtIIrOtGXyeft0tHWrXf5U4q7323R
107xoMgHkWaoY3xb6OSSuKSTafZ6I4PhFauU/ZNlfNPvnuo4Ba6qyon+XhL2Hfo7L4ewa17LlOgy
o0SyR3JqNGwKOzilrgCcfBCYyjUQbXEDhqtIh09gL8xBLR1LRY2m+ZWS6prbJa9O4ge5LD25958o
obf2r0dj1knreHOqfIsH1+Tqp/aVs3mvfOcOj6LlLwHHCy0ycVWsvzg9lpRAjgiUWnS1pGKxRgkr
79twshJKuQvSYh54TQvb3596sHwj4C6QTMo1EF4jr12VjzSZWuaxK1fs6YD3XHDJ+1JC7QBR3E8C
HuckybN3AqEZ9rHGxRBdtuRz1fG26T70Aieb+9HFQRhIzhsavivcExXLGv/VIi8IfRcGxKMV+Kc/
/RxoFitR4n2D3YUXu2EwPWDyVxZcQmMwFtGakYVeg5BrIuexXbQLKJkUao27V8M2V2rcAy0Ygi44
FQMFysAlL7MZGxl4CmYtl2Nbo5IDlIlK4q/txMWA8flcZyzRGMJziNbmiWDsiRZZYx3xnwmnD/h1
K7J4Q+lyGviIkCsXFjzdlS9ltbgAx/fiXam6vfY92+YjceJ/ZvbpmbhsarunwP7YwQsmxzke7z3e
LZvh3XpMC4i70djKNfQuB/imk163cWKVlCpDkZquYwLsucBGixXkR4ck5CfPEKhRCUNqQSevUrPg
nS1hdx/NNxaoONmrZ+/iDucBDBCZNYp8hq+G+mn0Jq7S83w47IfD/laoZkmDN/lR0Q9CQxkBuct3
kRlnm6eFhgnS4/S1wKESAb7hyJ8Z8ST0ObInOtk0vaLoqETYjUwkJYmBVAZgU0wnQuT4Q3h3NS+c
gIEgsRVTUp5vIvKTZo6cJxRQ2xMCnvi19lhsOaU7iVerb8TPnd3wPHItBYspwS+6JOHcXbOx6FtY
LqXNYG/1eAJ5eHSHiJMG7JSV2P/YELWQyujG/Qlsxmixzkttl6+mjTO0Opk3HSgTBZXNFL1Nz86s
FPshAKr0PCg5Q6+nv6RL0DhLfDONZX0maAcXB5dRH1KBQGkeMoOdFbC/cxT8IvQf+5yJmt9tEH9U
++xfCU41Ua/Z7guH9i2rTYecRE2w4GSAyezsUlQTZ6Ro+Ja8fB0lIOzprk5X3kW+UkpqOQmbiwCx
Q8TjqI8ACCgk+6FluR5VvkzZaPyD6ove9x1YrWV+Ga8dPp8AStNK4jUMipTlaDDspUPhKQaGHRgd
uIHl8Iu8DK1y6IyD9fTyfz3n4JxweTKzt6nUVmsDqblxFHpC7S1E4tpfffhBqaKCTc2m8hBIVro6
55w/zPi3IS//w1ovwQeImZqTpwoi4kJwo/9LCohV1i+RL3mlgJTeE8xqwZIRpTE5OiFBxPvwbGjO
ftzIdX+L23EJSi5TOp7zhqcKrmGMOuwmowmuurikEvnb7Im1Fu9oyT6v/5veZVQeWcQe3YEIySP+
hPat5s1v/sAcGlEIKtNyG932sW/8pC9HGcHZI4zYPt1055vV4uV8qNzfknAMgHcaQKFZyBdqKB5Y
ELMTRs8/cl85VtJo1wJMaAPjYwjKuSte1ik1G46Jgbwm6fRJuzkd7uAyS4J0g3Oo/n8m5LxSXSK2
XV5iYECuldThsANtEHNYhkAwRQ/rMx1yGIkvIMKv4G+3LhgbTB1J5/tDdWGYgO1iNcXOdk96JPka
7Rfl2joImS4pUhgLxXLSNZtJVx/Hjpaaje9FmxKs86r/Dv5NbWmQ2qwvA5zdQx2APlnnPQPn+pnR
OyOXNBvdGjWLk5DhP88sZr+HUmQOK5CiRzYAq+NaqAIHgyyOkmxBNvN+YA2zLJcQhjDhfyX3IXC/
aY7mpwg7EL+8nTwts/41X8tgIwcVpDxYu54HyRRQhkwlqLvjKfmODbgTlbhHeQNGrH3DoUERJzbN
PVgjVBMzFRoKyty6zmyAwt2vCO09WFqgOoQtqK/EGMLFfGJQT7GOhywX27Ea5Pgk3sf9PM42VBPE
5nvv+isaRgDGQo4ym2nnOhlyKrMEw7r017tMuhNaH0UXi82+BJV+unEqOtujzFuKbeNSZoqOyc0S
bp0Ppo89LSSFkrLYgWl4fXo8bvt5Eq9Zs5ear5sTL3jfps5Nnrzd82xSNOS9gUl9xt+HREPH+ZZe
TIkJ+UvS0/xS9OMKMtkxwx2ZIVEzAhNl2h4D1/BwhwygsFdMh/aIMmfFu2yH6PuZz7G46DmsS45D
Axbdg6M7xlyaCqdcf8DR3p3cprGowoAnD7uvGGwJEa0ulfQe4mLbDwKOcphNGOA4q9QAsjkdKHs4
99QB4sNUMuk7ulXMBMucQ7hOKSwgkA9N3MBIwvqbMvcwS/tY89rH62yT/JrUGTChpSOZnfNW1ugv
ZIWs1XiZOWQSc+znK14e9m26HttWzqh73N636PcbO/rW7MfEWOSF5WI7uGcYqy0BAdOaIL3NjwM1
7qBQ/K5z13lWhscdFdlTQFYxhteWOokVHQb4H1OEGNdAKblECL9bg6JBzierFN2i+HKp6qnaduL4
KwpUw2v02sennxyjymxKgw9CN/SC20JSbD6sp6C+pC3DlH7j2dnNFAFWVR1/JLoaI6/Hcllsz0Na
OVcAlcsO4cqNQuMj56lKoZPllLs/VheF124pXGMmc/FJMO96UBFH9KlLHooffr7loWOehK6BSiCb
5nXK82GGuSj1uXqTiLVTRWZ7uEUW5AI6NRzQjep/kebkNRa9cch2e7Zov5YSdyZkH9MCIUYoer4m
FCi0tlX04hyEKrwizkmwsQCYHpiMbJBYpkXOJxoskc6Wf7uq2qps+dJ/K8f5NOIrgKdY4A3dcTmb
2plC40Udq9q9wcKufLj8ifyYuWnLpVtlI/aVsvAasTZyqJX3945NhzQiZpGBicRDNmgHzBe1V2gz
4yqK4sQ3oZbaQWlhdI+jTAHGNNfMgeglnjxT8d2+7VNwOJ4cwMBebHiayOgWLg4Sx300rt+cLPbl
OUEdVJHoHO4bXqxQhElgx15pvQxLz276PyN7Gk/sAXnf1bJOvTR7pQCN6WANxJFX5Hee4RhY+vQi
IyGu6Kg1R0O2ZJPXiXRLWjG4ayhzuraNu5ZGrchMpC6JW8345Q6GZxzqED9sPgwZZ7pceEyMc1OY
LkIFEt9UsTpwaxF40+9G8fpVw70PokM9KE133HH7PsrRxIfR/5nGbnyEeuRqfEF/1Rg5t2eK4CUk
twvzp2+QKqM5kW3j5tVa4tgYZKdHRjmw5G8lcLR41dJZu1lw2h1YkmslbVwKpdRZ59p6KCJHjQTe
j6NEJSLJKbQFNyKX8dR4DavZWM+pz+B83dv5qP6nxo7QYwOmm7T98+yG++OTJw8IzY2tXLIehho+
/1WZJBVhcsZLj0Yj0iNfuZdBrjG9suIEIRPrMKQKgj7OlQpeONhiP1F6gSx66l4wO9pMfNfVLz+m
QiFaLVWBTUtVuYrd4uCUFt/mtXt+HH2kwxj/lCVvPMbkmXILwKsxNxFzAO5OZCGZsS8ske70R+HI
vuoSlvTocs9whucGMYQuwIQj5sPcRzeslzrIu22bS3f7Wc9/TCimSGOkEzMlcjjT9lftq24ClKBb
sqB8sFuJ9xbpB/vf6MRHX3QPRYsA/ScAGmSqS6laLlpxBTmsmTsUUVmhK3Q0y7d2u/Qv7fqp4Kll
Eshr0pmdlnWi0ESsPQdzkYzUcIGPr+axDKR2l6ts+ClhPEaXnKJFqgCHqvlm6v4668QPuZ0twXHg
y3+bLJ+ABZCxwClWofidJe5eSrT0hQpfLEj+kwOl5Kd8jjvVhxFq6a/GSjh52rTCpBlu2YBUh00W
y55LcglgRy37BohCmeAxpYxaW0/eukOdYhSbUZVgtp5FHFK1NFVHx4ksGRzs2DQr8SBBHu0LaALf
h2dmcULiB6ljy54z+tMNprodP5+C5nrsk4VmpGUwVOnBkhTwXhXZV2S0QEy237aRMMUdkZUf7ZYS
V7DMvhX44CyMPO7q03lPulBVlP9HpTCGG2EkfKIviMt8N3yllPzXifkMu6fevBNr8e5uJfz4/exx
JDu4EIYeA7YtQbIm1rVzfr4XDnAFKi1mvpdG4kej013U9PrkmyiDhryhQhdkeyzgOvl0jOUm9Ofb
L+qQg+qhA3ULQglaxWZsLy7FXzqlteMGnY8seqt5dj/0020mYeqiupdqX9o50fdmu0nrCOm4ciKC
vOqqm/lk+LXGtvndyU8b0xC9EpKUmBBO25eSSsD0prBomSG1L7puxxkC2p5zAPeggOMM2lCrEMmc
3XBk2/M31c45ICjEVJ0rWNNRMcpGD6C0K2LJb1xJGJIwsFvarEyslbCzKFA7vVs9t5aZhklCyXpS
FhIw2GVzYLsAOVrOG9lrOnR0g5ELVh4aU+RhuyHP+NKGaFbWQV0QGecAbKVZakF3BFK/cwiJADJA
jwkx/ljX+ryiZvsPriGFdb5cxdg29T0UQzdBQyIzt4te6zGEfyRMVXoXDNL2fRSAEqphRXKYylMZ
1OmpjOH+iY6R5gxDDRD3slnkFrhEvu/Hh+qlDGoDUyr1uJ+RXJdFA1LwPKzsq9mctrsZjhENCcQ2
6RniwxmN5WhuFHv+ZJpqSWYcPScpHDZ4WUyLh6IQzHToMYT22UoDnMQubuufZX2A4Ceb8Ndw8qJH
kOu8Ipz8gWegl9kvomuoazGzB/4A8Y9iTZ1SD+1HgKOT3OBOOOWgKd4pQ9ZnDgbWL+Yr4NSZArBH
/nkC/2o7OLgbCza9aJ9vggQZ7KHln6eBMEcjMhS0pW9/r7LZ9WUTWIwSMaKYjBggszpGJ197k35k
tjTS+5zFIquBjSUEfWVZ8y/fxD/GLrlhAf5PJec/bLzMEA++n/9p1Z4dFw8wXyrmdouImG9FR0MO
75+Lm0zO6PhUUavoTpeYsh5ojzkD1v/2jWopW/z+xd8s9M3Hx81Q1aCuRiEolFBqmezKBXpBjaU3
YliQ80ZAn0Iklin5BFwKGvEC3QHnD2M869sun3U2dZxmYIYKxUdV5tsJb9NvKneKsuI43VfwlGdS
DHGzXNcH4npqSVwe+43Eb+1nddNM6kiYIypOV/PuzcqiCloSjlGeykvtZocK25HlIrdDiCmH+1UP
mqLKh5EuJQCPLw9O/eNzqwU5s9XXCmr6KUkcwY2/qZRURwdPp4vjcYqxF7BK4eXDrRGdGxqoyj6P
o1LlbOGUxEpzTjNU2T3rH0lL7+lLa6NKjEnos10ajsHodMon5TKGw1P1PQRluY4ZbIx6CAFicWwv
/8WPk/x2eWfJH6goNnBmnD8heOuJQgzzift2v+CRZz9Ln4THXxOkSZB0B6WmhfasoY6ccyF4AuSc
suZacWKg6/CQfTF4o3rvkEI65pukNF7DvY83tHbQV4U9dAXnk/xpqZ0jzg1g2i4hT3Z+iZ6G7c93
pYtGUUGg3m01BdEyGcPcEFE5OeBCB6ahIHX+nj5Ow7BezvdFi48vOtO9tc0YQLqfjipMYb5Lklr5
sj9yocFPWyJhdjPy+2XOKatCqWqFGcUCdcebF4gFJbRAxqpKkTuS9687WW9rj768LMe9PKxwALL8
h6oX8bndQfvy1EGvKQ7/pdzT07c40xsd9QB6QkA+H4U9lZIZ+4yr7GPdbLlzl74sFXE6ksAehlGv
XqH7golimsxXTAvgXYTOyhgCp87aGCxUarcecm/dxiy8LRF0n1DPr1E3N51P9DRh+rxXMWGixG7I
eNolurGUrHzDqKgHGeyhCC7J2y1AqiwPIbD0OGaBYkiiuTqAzGh+35ZKIVYaoHXd/20GbUzYIJzi
4+UIzNl8whnwDNEoIdBOEXzqkgydL4qh4UjEz3pjsHRxqLobms/zOlHtWIokag/AYQ5KnmC0ASRc
zZunqOBW5oJXDKO0Slpqb1IDb8E41yDhkaeSNHH3je5d5GK2cd7AxRqw0C1Hks+UIyZrRLoRO35D
HdUsf4eaBVuXZeRjTTMprkGigHcpNezkqFkixsTyaASLWbdQzzbnbH0Nf9ifR2sJCUm4j7GWPF9F
gbeQZQ/OV/m6Va13L4lqJw9xEYsTmSaSjqkXlr8kQjtbfpQdQM71bfXBwiaqxp0KVkIIKnpt1KHd
c74P1K0Nq4ro3N47zBTY5sHZf16LvbOhlOmIgUlna0WXUhLXHeaz2w47Sw8UcZ2PGIpyAzNmDXgU
Jc9OArbTkcN32Cq+lrw7+hbH5fWyfvT3DdnmMpLKeF8MT6T56Dh0YrUL2aI3EyW48Z/bSw14khPH
tExqPJYdgaHGrTqOXyymIJZ6+9wPUNnAaRqX6c5fEd/Us16cFYsYCUdGWeBN1nwrQb4C5oq4d6wp
InVcje/deojXhJpo1g0bGbJdrZkc0trB5tODpDIAeykir1nA5jiXqqQiGWlmSpoP0ULz4EMXokyT
mWWvkKf9WXJH43OK/LruT0/q14k4t92H8MX5991UofbaNb0XxQhuzVVXHvDamKJKpLEHiNXbmtfC
oqS4hs+ibk8aehVE1RBwbNNU1JgBlUgGxFNcSDs28huNyzbsszPHb3Gvl4feZT5Z76r2lpVu60qG
ZX4yc9Hm/VMuTinvgFbik7I+QkW7QBR1wNtKUayVq7K8my7RR6g4bx2nFXjfCBpvhKrPSlw731dt
VIjWZ25sUx87BL7PC/2oeFXHnADYafkH6SLx4pf0+umF4Vc3jt0qg51NM6N6WzqS1ojgBNpI1IYe
xowdmUCXeJNIqIFrmYpx/xUXsmWot1gurM695xoGwnS/qnhAb2LqPCu74x6Qshcm1b0QiqFurDm3
3tLiZ6cIIWr1orxA2oqzRfeKXrGE9JjCZuxk0G51kCA3NbBd5U1nsV1kDsd1cqRikTpMUzlzIj6b
akgLaevDmuq7TPXqQPBc9QqN8m7DcVK9DyzOZKoTSw+GbntvsoTyhM6BWAxA60Wiex8l0DPkgoRJ
pu/BPRquFen46fqK0MOuwb1bisKFtAl6jI1+NIbnD0m/YrqtR0amaJB6yE0AcYfNndKzavKomuXY
mW6OTY5DpqawsY+z/gkQlOeIVL50B9s2bbPBrmzULeeJwIs38RyYqiuh6pbhiMRBp4QDSAP7InLm
lP9WiyUC8NSkk52yuRq0Vu43DyFZET2CXfbtm3YLsZTtLjbiXNVCtQNX4t8na6lWdcO2xSRR+o/3
5OnOJz/j+t+BZGsiypQfBree51YAbT/v/Vb6GPsGP68cRDdIQ2oN3jL7RlnWF3a//iUiOo0gEAU0
xPTj3BZ9BBXnqsLfpIJarQf9npN+c5ca8/vSQs1wfWQPzA3QFxuf0uKEd2F3+ZHpCifPg8HQP1wQ
Bj+c+Zl8PzTncEtkD7tBnxuLUgY8m3q6A5Synwogz0LsZpOWrxzF2vystsgtIWK3KEGmpa21e9Ce
zJdpZ+LvKuoo+5K4TashN7y66tazDnK+XLekhDXswYMzLLeVK9TZczyo5LYW4JfszjBST5Aq+3tz
Sf+4LN8BwHDKwlZ6xfUKG0+SlNwBAQjBSWvmm+PbPJC1ssKivknn/bWR0ufirEeQ1LCUv2uZtm1e
LgH7susj4uzXSgGSTf/FkivWvK19miQgMeaGp+R3HzrhIeVFrH+M3fO1y8l+MFSRC0g3YN3e4EGG
2gTJfq+6bki+LysxlFW/kinqSK2OnKmzEKU6NT9TNStiKLRgoqqh9OJslA25qahkE1oA2ZX56vbo
X5QE8EA935XuyHpsHhiRyFkPV+Fq4INPVPhHyPG58N8Jt+EoNYmmlrD2pYK/XkGNfjamDVKGNw1U
x9GlxOzseW1sEDYHSPjCbGqG47rd8DtAeJF/BA/Wt/riEzXt6kU2lm11d0cdh/Kaqo+enVy7gtSG
UNyh7XPSX9KlHbCZQ8UuHbrfPEwFZC4RPjUvQZnsLSLcahHv4wlQVeLxd722KcE7IXfo5UO/M2yr
cuSRq2doJfuNtQoxeEcsz2RCZWHhkIZLwfH8uLF3R6SdiSifDh5NlISKL9QOzvIU6WC/UOc7QMQ8
Mn4xX5hrIhtKy37ZoBhgKpRyHGNGsON+xUJ/whLty1vR7lMXFRpZUUkdAmLMXZ7GXwcsgKEBWKxR
qmM7exdB/MpaFOR6EDplXPNSdb1xDBcn/Ykw+w3z+50TtAap6gxIUFQn4pzy0938EGDJBYClyY/2
fnhVPXCbjI5oYxp/qOYWjaWI67MjeVGQOGIDkyJDdXVA7ihHPM3ZO8yj3cbqrBQJsN88KLYEOTJx
jrd80qJUa8SRlU8gcIBDnmtJz3UxGe+xa3Mh4oWJnTR9Rt34OR0cvQtwAdUzV5ixAO1O+xZVzm8W
+OhpCzlXtstIvmEuMcfHK5RS37Eb0G0PbxoSoEwcxjtAKbAWFoO5KjYoW1AMyiYAkuTkIJKYCA1/
nM0VEB3zDu4+VT2uG2xWtS3xhh56GO3g+pABg+HvGKlMKe0zkh/A/EGGD3UTtQ6TtEgejeP4YFel
ujqh0clmp0uwNzgbGXWxYMUT2EqYvOp6A/kuVgU5v8YR2Liajx+4obxLf4/EEf36+n7gluW4CKOk
sWj53/ASr3OJnrfqkj+OnD6cpsDd25Y41An4zOOgSDc0Rrxa6ZnYbAV231Rt6A5BCYnDKHZm8bcK
nmlIKPmjhUdTBxoCMnwrnzWQYzJKosOrwSXQKDNYJHnLyekd52WMmj2E9yZki4G1YdVDnSLfuYM1
19t5+55H2ijEyHXGlK1cFFo4vPncO5DHbXQGjvVtSB7rlIVdIHC979CvSSaD3DdzX+dkUeU8QJN5
IYrg7+EXsdrO1NT8Kmb90EVjxf3z1Sm49hy6x9gaU0Y//pXmrw8o1lj8tMI23Lzs2EEk+PrPhM+K
o0eX9/jmWYYkkiTvBRuSg4+mFABP9/T9LVCF208MdcqN+c2f6xA+WK6yPiZm180svYs+UcqADeuc
nPvhhATkZB9+tPFkw580818dV9pJqaNRZwrnF3EFMfw93fKdGh59ttOzvmBLzuE/KAdeFeIpUPcV
vdGDfyI4qbjtp1E1Pl1IAA8RqiOdLOeWsT5BXKFokNXIxUVTTYxPTja9QMipmFVlsEtYJqmuRNPO
Aius+xDMwc2VHLCJnbX+aKH05MBVomdhX/mu+0jYIhe+mzHsgmqTlbaltW0T1UFl8Wo9RsjwgIXe
+rLAqpu4smL1IfJgAJL4TCWdPGLI00j2gEKviW0+mlKNbjebRApRa4EqjZJAcfxAedLgpX9c6MAi
dAcrNVH2YzivLwq7nsOGw3vqZdY9xsUzBTiptjNtrPER4BIzZ1uZjz3OHks7VuxHQNA73lefQZkF
DBB6c6YniRS30wl4s9wLZszd7zIC2cee3gKwbECHw8ldLBbYeia3ZuX13Ofigx4OQzjKuVHuSIfa
jeOYa4doECQ8IA/igfPApVcrONGSp5nO+ay3WTlgjJq/FoSSyrKpdvL8+dPt5DuCPr2IcL9lxbMw
sTD65i6dmL+WByx63WIj8zXcrHToJintD2zxE+JKYUXMTlAZ67RccWim+pQz0K8Av62674wiVsE4
rqOeH1jSBj8QfoBTMSYmKlV/BBsbOHcHcF+uU4RaWhLsp5O4qru0oBHbzh9TovH4GIQR/4auFSFB
4SWgx2utiBnCxUfDFjXluKH/WC6a5BrgUzoHX7xhH8h1Af/MSd/27tnJGV3VUgV1wYzNMfgjnRpe
LCi0z63rE/gNoDkU1ZXS7UyQ+6Ca7oBDOPhyTQkijYXWnQRxqsgTxRH3TsPVXK10f5FzqHenD+VC
lGYWJ2v1tpYS9UtCMKbgomwnFUQxmtpz7aDjaBWbLv0/JXoeE+2RjgUUsfwNRXN4Lcp37liBm7ZD
PgPp6Q/ZCQLmdho4Vc2Iag/dknwi0/X9lYaaRcMsMaR8o+m0ztFAyvfEf0tHh/nvpjRJBC02DG7Y
UeVBCrmj45FcDM7Xg3hoJRQLaZiXWnIP56KC6XMfgYkUh1DZ9ZsK2IoT09wHKwCevvdlYvs8F2E9
AKXMZFM/4c8ztKYnX+P1IEc66yLM61tRrX6COgxyihYvEmRQ2ABzl5dCmLH7i+UoXMgdoU0QSFf9
26Hr45ZSN6cI+eAsWW1p9pDEGWLrekgJFsdoEmTAOpMmmQKTgWAwRfy2PM+t7cXHmuPMHANpcOll
qyyNs+lOYukROAPvB3mnhChPGI+P1MgYLA30upWPcS4sXHZSz4rla7o+avWJLdyIUriNhhlBr3FM
UEC1DAOrUN/y4ZzkiOfN+hK5NqGxJLvpWyfKPb7yXAz/3TWmOqW/Z8TbNHaXvXGpECiaH4wmOeHD
IFEAqaeOvPM0R+zq3u36PVg0DGW+yWSW0L9USJVsDuNk1+POPXxbi+2vV+S61MWVETIk/GDbi3xv
2wtrLCey487oSn/VZCmlf8CvxlQXPKG2jF9KgcLVT42w44pR/JGp3I01iUlCFP26BIUn9qTuTut3
NmT/z1Z3Xv4n9psuuCSgpZuFrQrgQrBAuVKfV9ZyK5r2v2IrxP3Q/fLJigGr+EWnxf3BqQ1MGSMH
KVDCbRIOtX1sS7gFHpFuNaRlreP1HCpNggtqYJkxDBB1QxD1vffgBN3QLmVWMo6BJ+jkN+xnW07s
Isl3QoZ2WGIAceRb7OBZVFKnHbJHfVhI5ZlCpQm4bmMSdxPrAFRflqN4yDrsJL2AAhmeu58KaBoF
9z7cViwl3TBcWWK7QgT4UKIcnO/y2nkdju3quyOLRLKeRgt6P6P7NFFxlDEEIw7xflJpGaPVw6bk
u0Bf0o3zvebSlR7HNjVusPyqZKmAFaS8Rs9YTJEtoy2M7O1QUozVz4T9iYVVzBMEsb29VHZjeUW+
MhkfRm1iydQ/KeSS/UF6zjT1Q8YWlnZyeHB0nxRCGrTCDqidRAtWfRBZ++Zc4FNzYTXQvH0bjvW1
G7Q8aDXmhUnSJzex2PSR3JreqOVBv6DJC4bzVW6dhPcvkfPcl6eWQFHmxpQ48XKOD9mOXONpR4uj
fY6rcAAEeBphQzfeOOf8r8xDuM91BjpvWhmJ3WnBNYNlvhRMmJztMQD1Jx5lxKrRT/JfhT/hwzjy
GGi/a2b6bV7qckNvJuAxMPxOgIvAwnZfzWy5X9REnS5dT38VJJU7vQnOJrKGav0At06WiZgbL2OS
BjFb424M85iOG+Ko54tOqfZiTJH1WXuL/GMzWubnaFjnLdcTzHMsv9IiaxdtGcjuwdrtkcUI32i2
JAGcYOOi1VwDPz2S1l3O8+mm4PEXqJU/62b+TSraB6lYT7o+5CgL5RUPXITRwE1RUTXJfhFxiKW9
Pb1kkcJRkkFNr83eOCwxKJ8vWAanMbunuyxrjvMiik8k8+Bkmc8olPUyBq0pbBwGuQBegiIASV3v
zw54XFiZ/5RiBEKPz+lF/6ONN50jBv5CjwREvPSj8c1Y3idtAkATyEPv72dngwSkH9Z7JVqfOlnK
M83UFe0DR/14cM0ncvajDW9jNoscBcxLGU3y2mNMlDGyW0GFtmrqCy63NWG9oqrobq25Zo7JuTlD
iAl8OF9kcundfztpCj4AU/MNhz+wm/1LEQpvmFPvofsj1KmdFHdjPMPPlNqe0UzcF7JT4kjTDXFE
1TJAdMAzWdhpZ6E+sXoM9DY+x0Ekcz1rDth+GJvfbqWVf0Kvxh+Fuc8IyQhUi/HDKXnbPh+cBIrJ
A7snudA6/39/8673lv4AjCko0db40cBByS4gQm9oW4GZHUkKeEnrD4c3x910x9QyyL1nRUeAdtrG
Q2UFtvIg2b1gd/gbpiTF+eacTjkR/3hPjzQiBK9TPj8rppeaWjSvGxtdnjIIxysfEG9OIYPNO1AZ
bK7xKBs/leu0k/gTrbudBEXIQJ9pW4V04WDQ6Ezg4gzaDtU/uOb3DUDjcGJJAuis/zTCMNML+7Kk
E809eeD/fF3gy+X+hQhx2AmyWeVC0qqpsGQEvImNNoIwl1Aj2V0lOhu6kQ/CcUV0m7+sT+VxzT3b
lyjo+Yg0299+xchkiwjAmjg2QxQDJi/exwKM2srVNhocoTBXbXxGqYIxw+ntIB8btIy0vroUH5Gu
AiXV0m0GsK31Zws3neegCToouLSa/uxiL/Dh6SoAamYF/iE+SKhfLMSD4IovorbtxDa6T9RPbub/
AnQnNYTWDhwCU8HHxvhB6qzL2fZhquu7qcNVg9MKtr0i1BLlPWXeGUeU1mZmkrOysk+EAh8m6Gfx
L8X82YjuqwwFZIQ4owa9uFESZzhKkOWxwmGp9qo7scn7+xctYwPY5qnYdSdCdUR9FFp1YtQYGjN7
hzl1qAbvm2BkCHa4kxKSz4lberiXwyDEbgU01bcztdSm6rth/wAo9t8Hwfd89MsfwRGKudH05kuy
NEVQpEthpK7/A0XXQy58NX/NkWDTnJNdNMLSK282v4npoNvhMZBCmiA++oe00zjnRf+kJAlX0VYw
LyDsa3CDuE6X8G5Tdbq9ABHmP7r/9lexw6zvxYXjFH8IOhqwr27/eT9V4C0qWYOsjKYNVxe0Tu+X
A7WBbVgU2Wp3gC8Z8Oi44OayYzQW2xzpQ78dVriPzgjP9kSRPfnKWzIfJKrNVSlpkvThPXez8gZX
yV0QAk4ge62mn9fidp5aJoBsMe7kiRLmcGJK1NXKAcOI7cktGZ5whsPNy1BlKjoKKKr63yxxBxjb
9XFps6rs8M+foFp0o0qysfE90SO8GD6RvgVK29kIqC9wOloBoAH0E/FO4Af0gia16qGlPJKr3PXM
gBG0u4JaRhelzPLq8ajuO0oPaRih3pMxxtXobx7jYALrimwNEZF+jxiu7OriPPdPIdkLC/X7Mt/P
CStg4MkTycpAEWpqr3d0xrzTgusyJlQgkQgZNMHxLZh+V2BAfADEyCaRwMgvmTeaYzf69TtM3QVb
XEfQai8rm77GkzBxm1rAUykdFjs0Som23tm6s0kww6GBujpwHq0SMgiv/9/6sAxCovdRrBiR3FRS
10z/7Lw9h6vINpTeV0BCIfMlnb/n2SKaXpYGgn4udNVPou8eK8A92uArT9oW9S31c1iqmSBlXtap
Gipg0GXVgFeK2Uqpm/gdSFm8Md06yJIgIG/jpRHEwn7z5z8qOmk2mhE+g1SzB7Ux/OxS9XxLWv1z
OpbjVz5PP2ScqGKhrK2J3EHh+B6RzR1aGkt9kb5kKGfloyP+M/IAqmsSc/XgovG1dT5BMllXzkcU
hR5SxuhYBNuitqkNvbQYoU4ihnbYqgnO1fP5Tjdv0RpQQstVMGAT4/g7qY8Hd7/Qay/RvqaSSh3w
TnwjAz/0c6WF4hALQRdrp/s49hUQGbkqTD2eVr9WEEMNlc1pRCFLeHX+kIvRNH5Q6MzVLe47wPi4
am8qnuk1QKPhIKLQuocUzZLNdZpdXddYFdnxGc3RKoh1mBSbPVdkFS+3NarP1tvaGkWS2ONvFV45
1Zc4VFTM/bemaobdP9Iaag3cRU0cmH0EpjuuqZ3r2Q0s0l42I45cC0GS1YwlsBb9phJjXGD2EZO4
GsMJ26KV4srcjDwemU76ETbrakzNhoZ7OYHcxgP8+KjVpUM4ezSIdDzdkwp93vGXfiNCkU2f1vuZ
1ISC+qMiJ0HrkNhCpskLm7P0dL4k8zGSenmzaSD1Q2NBWEkXZfdTbCbqG7wQ6xCiE+SEwDXKL2zv
lq2Q6J3V3zIgqSw0wuPyv9GNdmFPSCvIhXNkYzysIDeK78J/6/LAFz1StdRqO3WY0Ko3uRHPfQKK
R/rZ5/p67qIwd0AJa/eX/2QwCvbgzuoOlgo4UPOCz9ahCl+T56MnD8igl0/hiOyP42OSVRXu4enH
aVAOSefShvuGCnuvA7lQLvRSt86fFVxSfMQzUMvGOHSckSvU3L+oQsLenqwrsDoGOxYoD4gOq7iP
ooRgAuzWYa9Q6QMeCCbpKot+8lJpnQ9KmtjIx+QDnHzgNoV5u5exkPHBMV5mHwZnaYM4atzIQDW4
gcTFPa7hy74MhEojlt5ii6weeOrN+hmy+lHC+KnfVhzMjHhXzwEVoATT5F7BtI8xwM70TiE0bS2V
zdJXD8GD+KTdzLs/GZn49Zw4R8a8zYrEJvJXUmICo/LXlXifCC/XhHJ/Ppzf8XxFiBGKPFyR5kMG
O4noha3gHsC+6SdiS4tY8iB/9KfKdfzFyzYl316qeF8Ja2pILuQhsRtWEWjoXrOtqxEu0llPxXxV
Vc/twJI2WE+LxJBik/TLUsVcN3qEeWw21gzy/kmDOJctkuVdhdChwWM2h6yzRWbp9LhyZshmxh6T
BVMWJdo9pprKO/d8q/os4hPebiWYWIfdLL+uezyXGAdTGZ8vhKijGO1CKs/JlMF79cGD8l+1bnow
UTn0uOqnHRyXrf/jJuNsdeFonVHCzAf2OSVVXjaJeLWjRFV3056UlgJLmvU6M+bpjgstFyaC9iyT
wpJZh2votyojWvkd3BXD4xV66EPguPYmZB7qkczsuSi/pZmNLQDtgg/QYH/nWaCCrHIuEWac3B5k
jfRGkPwLcM+G0Wm+dKlXXqVyzfLZa5CRRnr2NL2H1orVE6uCvJqOVzqezhgHqrQ0wLlAyp+dU+vV
9qwfrUF6L7S27IHAlR4TD5WSBfl6psCNNij2F2rZTIxEpQu06GYH4OYk8u9MeD1QNsilwCKbr5nc
5DlFt9IAoti5F9pJT/nqQQgmzq/omLVpwVgDRqgOkI9OqTvJ4c9ue3htcZ4s+L/fvMZDIFIoIwDz
Z29U+qiEkfHUQ/vA88OZV6jByNEd5a4zERuZNeYDD2abFl51oHnHvekb5nbTW2hzb5jn/kYaHmir
LYDcsWWvWL/L7u2fYRfOhrOqjVSVw1QvddFVChQg2tKRzMPSmhj5WZgYB9Q3nVg+pvSTs3aoGo+h
9KnrNUGCqbgaVJWaW33mI9iTRmWjzq6KJ+cDDKZSXaAkMhWt/kJ+aITYcGQVPuc+YuSPZrksZoDW
r7YJ5Lj6uYDoxLc2nYsN9InZ3tBfjaH5492uWqb3qTwTqDVs6ZXnL3SDPCGNoqsYfnBcTWazsBlf
vOJ3rZrUnTo4gg8+Knrd8RsChfWcIior0c4RB5MK+K/0uPBWOYC/uF/YckmXIDm5Sw2FvD0qtyPz
h36dDQLS3ogplrq4A/uqveJcwgdtxZl3yKf4z0W3qgh5Q758Ch9AYpWR5j4oNHFFFTTdWhiGWsvF
0AkmzZZf4ZKFNa/hvfyzbMbqKHnz/tx5nzQgh7k8+R6z0aRNvNUldDHkJeVNQDiKMb1olN4FBPFl
Gby5rn5qy7i9JSha7qee84cwFywVV/+D0nmQu57d9vY/dS9fIdT8mDHbY4FsNdoAQcCh3nsXCx99
+JlMR/KjGJFfcSzn6AKu2qmsbvUJCIJ8wTxNL2UdFzkesqakAX1AoTdtYoAp0GCzkrEYxunPI8lC
oBztRVvqq5f0TeBtfoueLBs1Ss3t1Cow+5UzuRlwQuomZ/vxG0pm8ksKBb+ffgEGn5mb4LDbYqtU
UQ+QoeWWgevIOBl1tc3nigbDq07CF7FBPcbP3mvpIZcYugtVpnQdkEPLZaeJrcUSd5RcDE+rD7x2
q5sSG0f+8ghieIZKP7meNao/3kcrbIFWWaSrnzGTM6fIqYtVmDf28vKxmW7jSAcbp0OmKwf1BhFT
dozD2jx0NoYlTeDVuD2c4Kzkb1aNeB5kYkk0UXGNSYr66dkjqZ4FLy8Vqthjj9o876+JcC9TiAY2
w2djKEKiyLNfcpOiUE+ItVtdDJRhtqhFvmMZgz/j+lfO9LUqGGO4sekfQmKx7CDKgHqPYf+53ceM
k5x2B6wBfy+JktRJrDiIHBd8weWKUNfK6nizqWvV3JSmweXci1HQXNxMWyYWDDH4A7onzb7x7sYO
+3uT1aW7u19tbqaOinXw0RRm5gbRpF8xeajQobn04zclfEj5bX7iwFi6I+9GezNxxah/gN9g4Tgi
TU2B2rUr6Gw1KFQuURr7dTDZv0dGeU90YbbQU8OXk8B5kuwZ7R9+7sVmGinSogvtQkigsuHpovIz
4S2zJ9li2zNvZ2dAlgqEA6Uu0icOVsHsWqqGvInWGAMY5qJUCJfkA7/rRzoU918wcsHOh0QeDuDQ
9+2FraAWW67a1iQamDf9avxKr+zoxSUs7W7NVDoOQMd6avUuOBBM9f5Js1S7HIA3b3pNn8PyY2Hu
D50IKESsQNYsU5sxaKXUHkmXsuH6H6IF0gUVTn2NOdvgfZSkPE+BQdd4NBPdIRwhvYxtThGG0MzT
Y1AkaSTBJTQyAPBMiyq/GOZFFajkP/ttkaPLuLhZw05WEss0qpfp7b+3CnC5r3Szj9ujv9n+V2Ng
uECzy4jBaSG13/KGzlZGEIjjfz+w33mlLeuTI/70FcJkqbEEe+j+8R1BYVJbz/FpikA3LGAIPQVD
+Uf2hkzBL8LRV7NQC+mtcfgh9BFzqCC2vj7n4Np+8lCVzHBOgI6HWvxKje3+movb9GlJn1tOG/9M
eeRuEUNWcv/Ebk4frxz1mG/5byAPHfN52huIQMuvumrDqXw0Hvq2K/murhzArqa7PTW9lDYaptMn
4e1WvJsldTZvyOCMUWo7Y1yVhB0H62t4VM5HJ2EMrItR4lewH4bSLv26g3CjThXouoOoYKwZiGsj
ATkhhWvODyEOQrDVQd1+1Nyexx1CovM4FfxdjWDbhaiaXjDiBfT18uANJQoTGRgcjciieL0L7BZz
bvIkeGiKnedYNYqIW84dcIpTTNtUJELgOZBSPJUPgMUvmZ5PtxfqEyV9Ic4ZpMgbePJ/wSmbX6q0
wWg/XboBfW0VvajHdE7DhGCtFuB4FbrcrPITtl/YzBeAroP6qsqFN8c+HD3CguR+4VnIaR2xS3z5
YgWvGioE/6cHS+ZVOC+m2XrvrW+JGkA/OsveHhAB8Z3tJa3vEYjmjUr8E569ZYFdz9Z3lT3oOVli
hOVdih4uxoYBTT1axwkRDLMBsFcC1+T6ejfJ0cd7YgkIlKCalZ29CO7/VRoLOIz5rZ38v6dtmksD
5u8fjKJTesQaBhqfGlENf8cmiGdneIwUs1CUK90/TaEBQFgp7Hiuo8lIT0AbpWqoOk5evVD9m21b
abEwZ6B0pasUqCCEbz/3ufpc3NR9q69XOQFBbG1jozMOEgrjJsmqU2BlX/tIhiTAc+SyK1AiieZS
A9HzJsAvzqoZfOA/CKDFocHxcaZtSpJbhAOCDFblxX9WNK6Z3RPZQN8yolzwdRuqCZWfJaEN4S2t
WAsDU8tzAfry0LDMPYAB0rq92Ddpn9N/eYYWI7I+uEQEmn7N+8AMU/3BOwt3EH5Nped7MspcHo1p
dgKwVN/453QGfRMGbdkzo6QnTNaD8DG2PjtfniFnFNXF27LmKF6ebFeXm+v7Jd5BgbpVR+dCCXK5
uswyNC88W+iPPm8qab+PWML+d4lzxzAHyv54v8JTWwbDhRkgLV8lyKq5KdHQf0yt4S/L6gycTFuq
8Y5LclKk8Vv0uFoIf0XWJKhyJ922Wys+AuxYyEVRIVDkTZrNHN2Q6SbTMqNvqjsL1xsXMYCiOs9B
2SdJqVy/7+8d5OWq+o5yFduY1TR5wwVJmxrJGF+sMMWlNZHcqlNNTO3rAYypOCnfaB843MUkhE6w
xx6E4TZ4c9moQh/RPEUUbO1mHExJI2sW/+srvfNz7FAL93nT1KHp1nKY/Si99tN8vpkzsBPGC5Mc
hLCCdTQ70PTgORLnYixEwVL9Jwl4YSJZNzvBeqvRXoN+Mju0g56ZG1iT2ruuDDdDCgpmXeaGEMO2
47zLFXbYqE3tYePnJy3IHf8+eV6PBuSHN8qYw2xMtbhx+1d3xIyVRyRb13H6ohFB5EXK7I4Fa8y/
EIKHB3MwUtRPG17rfcCieXsfI91ij1kyGqOKgfduZ73hTooDm70mf3tCREruQ87oY3IZTScO7EVW
k9rV1TvLEz7gZj6q30BEQpaT8j19lEZnWvVQf46yA9qu5w4Ayehhkt7IwE7QGGQRhqCweUb99ToO
zA2n1xe8GZL0kQkss/C4p2Cpu+LUQB95QkMRCY1YHV2M9W1aqd1e5Ry1bvopAWxsKn26g7hnk8h6
/IO8e0RcH7n8dGw7KB+lyWACVq/8QjJJYwHyLGX1tBW0cnPwFPspnYhOGNU8GosZ+d8iGfHTsLGn
WaFLhGgFNfzF8X78F6WqxNu9ne8D7Inkm7Kezdq8Tfloz6Qzb9zfyrXtLuDNMFgndjHvdJ+D+c8c
69OzRSfUUniXEweaXH1WVcoj8c/zUgjR42PGoH0jluSIZtlT7lat0qSp3zhl/viSKGRyPOPlH7xD
dOlOH7kQ7dPptyZXkItGt/ukiFaMD+QEd8xUaSxN9kTJfp8L9GeIwB5aSVMtJfcjcIHm/XEAGsas
BU5eLiRBEltrElBTCIbi8Fg7bFys5A8qNTVfn6G6b6KReovEPVnCWtMc2/TB+D0aUuhkJrVBLumY
oaVWglDUUpQv8NeIQm+1poIYQhTlj6+fCM0ixuA6PJJAHeBhQbkrwEL5zjP/n//NIx4S5M/Ow5bZ
EFXmVHCldEaxlz/spXFYoRgJYmYkNAojys5tRr9r1RRsUU+TPNwJOjw839SknKaXM8X7jwaQ1LJj
/G11i4k6u+T3uf5+tJwDg38XArDJhlwScewtOnr1Nf1kTL6LmWubcZscFZdPYUgADRs0J1yvQ7kD
YDQXFfNxXTJH8h5sOhanXRzwZ7HVBlwSqhB6o2ODNABkcNZ6FGA041zDte7leYcGQda9fK9rqWfB
d35AQnShD0frUeQu9CrA0opdMPFi8pyQYp65t77F5xA2nDoRAdr771HAIyr3ipUuhUG7x7vKrNGa
9IkjrxZY+VvtWXjODSXl/53DZJQ4IAMYGp45MTom0eLP56dvroIbyr+qvQ8TUmumUFLXR46zCIxs
jYPqJmojQ19W35zQxpcez2+BivJ0VsEV58MMraApiIKoJDqtuzyWH9LFvZ9BaWVGkyGpeQgJlXQg
RR/NNOZ9jr3V783wt4I6+C3j1rr3pWRwVGNeyHjpydiU8jULvLNm2ON1RF9BjKZOgQUOmHWV35km
Vv2WIUQ2YKRVa8CD1HWFP+3LuQmBAJTNddnVqTUw8BgkRAlJrv0bOuYRvRZSxm9XdKTiIkPZdpeJ
0sIr9hQ4A+0nb6NSjHafxl52KX2ecgdjhmC+3Eq/Nk3hN0fGyphzLdSEs/JyEBQ26mZ/LTnOb4ui
L6vIki7z53Z+DIffTvuAZMzBntpcp1NltSVjnHgy2tiQ6e+7wFlS5kj7QxVuI1dLFbZjvu7mi9/5
CHef3SCbdob3A2UGJyvYgoAbuVDydUIiq3ap+IsCljMW+5Gcl6KcBvyxizWdMYu+Xdomi8cRx4Pd
QeYxy99HscRzSXkPw3g/3RfBh4cq0SStbMvBD+w/07YRrsRQpu2FQYJfgHRzcJEnei5/8BSHRR/z
otfDTTPhEHvbi+erx6XcevRj29ItBkd8UJWVPdzWcPlBgCZDCrqT0B/Z+IzkHAWld7mvhtdCYHu/
F9gnfvOYxUcQfGeXQsXPrZuFktn8qCJ9SN+uHwYtR9zpfAsG9uYlx3S3xhrBJ7TxHhjbH9zhLNEh
wVGsUIUJyimhPbBEMVSGFFthv7FUyMyQCrYkYc3pJLXziRRPIzLBXGQSiCw+Ed0YHAHiFFy0gQHK
j1LfmnrilCriHo1T0SqmY5gyKVPLlgYOqFc5OtHDqiShaHoQNLiK2j2/d7UaTTNDKCYH4ihEJLAI
bq9c0QetAZQvLZx3AStE8pXsnBSU4VPfjaFQuKKoTvQn9RTZQOL8lRTNLAEOy4rkkelMp65swtaO
djdcyUzms1WmEX3UpVaVgIdR4x0tbIJyBgCQ2OdZiBTv+yVzPwSq3SNTwqFUdrJSBgMf+SGhiO7u
Lw0pLbAah++k24IJXytgO02eXyIMj1HclQYg9YUx8hXP4kvdtDlp/E6ZQBGAjEwl2et9IpjSADfE
/CFyH0MEYvKbfkLmW4OEB4w3jy82m2jxzvedUBpDUBW7pRA4WvsAu+6EU3Jp62itj2Jj2YhCWZCu
kyWMmOxamenz2ufVHcD4gARG7+zRYSpukn7CqYXWVd0HSOShWESLCD0ooTjGImrOOB84n+ZS8dPy
OUZUGRdSIF+Nd3qpfRz5GVZ6/YJa7PI8HKTQiAwkoxc/HK5FwVKe6Z96Tle8H7TJXQB3UIcoEiYu
4lqsDlf1Uca3E/XR7flGpe3yLXDCsgwC+Fu2S3sAT9jr5dx2eD0/tDh8ZHO5ALqNblB7sw0SxYpn
1oi37WArfD7Ce9USL9i9NqouqYwXPZ7FjAFSIbGGmdmgSGxW1QAXQt2xVzIRGxcKu9qV6NN3Pw0w
+ssxO2R1HaOfzafc8eqnv+CjUSU8QJnsyB09XbHxXEejwEojqYosupW5lJZLSP+PpHKDUM+Nb8Bf
8sq9Li7akhaq6xg8S/TsiGP4WfpUlJlxs+amZlhZQanPY98WNLoG+/1vWjONU2cOLKlv5T5pDSzt
MDTPy1IhOltGsda+cdvwDd7MHoVe/ZXqO0AZBHO45QlE1HLbOq8AUFyXNkL9EP4PbJvKkK4hKu7K
wmYYt9FIm97tcFTpWkdrUD5V3dbqX7XYstyqGTS2dzkokkntTFyWV1rUywqqT8Yl8RTB4r88Kkkx
jqYcZE+QpWfPtHcBnZE35pXPWSx3EDjHtbhoxN84RfimB257N1mtym4CTyP7Vxqdwi/5pPJfFtVD
FXSBhe3NOojTvHNUebNpySKFj1/tiJYj7rziB2w0UWUTLmyFIOayUjHFE5inUnjhXNlyxJT+qeAo
+wXr8O5g3d5udHQSedUm4BLrLbETr1/s/RN6Fm7TSpFV3q+rc6diH7hhWBjkVLBZS6NN6nLStxyG
snksA9CEtdXmaTPRSJRwzifsTXj6ot2O4A6X1jkwiQP00NtOMxUmReY0fPJsXLANQiimTJ6JfhA7
lCudPcBKcTuDBtN05wFvBmZwR2kRhNcqdmm8evpzLCCJXLHlWsC7fw4WN7cq/PKkWrp8PqztY6TC
HxP/c9QaAASrhiuSiEk+DHxDXDkqkbV2iS05YY2X0kO/G/Jsjc1j1ohIEC97N5fV2Itaod8Lkhy+
uJAXw5pkypDtTES77kPYPScQUNohwD9i9QxWlYXGRqOH26U116cB5rzPCfmgGyGLvzVhe3173wlx
m7YQPyftMmCn+8xZKMHJAk26lVoDUvUeGVaGrfTavaMZYTgyu5nPIfJLTjpI100yC5dXUDoye+cL
iwldfi/phbBiFiXA/tXV+G61VtC9sGxQaWENqn8K8TVp/khgxN3AaMTaN8MoWIZ3l0YfwRQrqOSj
/WV0COdwQXKSD3/OqeYunvYT3+Ai18TIydrvi5+FoqDUJ0z2yAmgJllKHG3rhtuoZaOqqyL5IBdk
EMqgdq2Fy+jNQV60BkxwT0OC4YYo2YCekSgRawsGKsxP8t58auzAs30Av+ye1qVluVOnjUueBdha
SEQ1GRawEK7o0MQXXUS/Yd9v+mois9fBl6mg4nqHZp5D/wEtP6Fjspykek7MhBFDGdnIYqATR6Lx
BZc4fh7h9lhP3Stwuv6IutPgQ+YZERO6Yf5e6CR3OJlLAORHUv6YKN4zYABgis/jJ+KHB7/WKuRD
8KDR+cx726aFoNTQLZHEPapF59pdbBJTOh+ElnYgKGXYe0IYo03hrt1gmfYryIH/qLF+NgbYJq4v
kSkWF8Sycp1s/0S6vKhljd7nGkLrW7lvzBpKFdLOGgDeV19Nc5QwNeb36iygEzIv1o7g8v2x49Az
mIhyEvPRVrXFiFv67A7Oqx712+iPh/4E/KEH3GHwNDFCb+UwlJuGYAv3UkC02tc3lCYOpUwIIBkI
v59aDeMT3vpdsu8gkiWU4I3uj9tlYUpUN4zEL9FS4PqM/rPAyV4753ce4Poy+BK6KXPvktgU++3a
7beeIdTMcwESyazxf8E60x/f+LulvEA/l5LDsEA5jal6nCDw3iDtKs0cREGypFf04xjcN2D18+MV
q8tfFU8Re9ZZMQF3qnmM9ltj0J/xcLbcWPcEMEFSGXsTo8Xwy99FUO2cw2Mh3/a7tHScMFPQSi69
PePNMdj+rzVVrwwFpz/CzPx/Vd0khx+3au5xf5Gs5raTxjwoWAh0vCHa8OU4R9MFmgUfMIZpx33R
Nw/ORoIJPiqqyVfHZfFMFkKEWCrG/79QrCFxC7XoEkgmEAaPf1bueEqLoAtdC8s89M4XBSasmaZF
w/5iS7nQKNt99QuKIVKPzlaiv4T3Q/+RkOT0en+WUxCL1Pn2/VUveD8IMn+8Uwfv/32Ntffx4LYp
SvUa7wuSMS7dQFn7VYF5jLgX5n+VB19djPEmh7eEfZaG+kkWTmDtNyuEQAgfhwY5Q+KoMXBFxThX
3QO/cynI7+Jl9OVrYPhouQM8SNqAHHlbSPCLVNVKamBWg1VFHDE4DUkjVQgAttrbj1utwsAjn/4l
F97/1djsKfJEIHmTZzLan7GjABkzUNgrbDFiKp6hGIqh+MikYHfmrZKTNhGgfCBB/EvV16zn+Hrf
zFGuTX10FqkVUvPET6eh62sEArbO7WUMs/3+iuklbGfjYt67HxiGz+IUzXjfSgf11Rr3IT+lYnHu
9vdFIequnKbJB3+uJ1gg8M+nMmb1magFJDWCcmWbTC5VU25BH3q2r985nemr1rFRj4DKgg4ijngp
gGxqHNF25reVOdgDaHgrGpJggLUU9zeqG/9m+S7Z0k1oNUcwsGZQqd70BUM0EfpjxjdVBn39s+6D
FCgLxMILJT5w7h6+GsWIlzG9NxBYMQFjAyPhGCJ05L7qxJtislK9BvfgGCRGPKkNhAfSq2VRdfTM
i+5fPISB2pEEzLnDScpvRpbqZmsmY1FbSQmZbm9n/x3MwV9+n042G28pRvRdNlamfNrTGoMGPkyW
EZxOyIyT8uN1v4cjDsTsCywuGLSqfSKn0kWgfY5WLtLObeeA0Cc80lr5pzH9MxZhZQyDyzgn579e
WggueSlCGU9t/AG1mjm5CgYxiO5PXuX60w/h54iqpG7A1ymszjK+V5A38mmjGdQC6ShwSUlXihzj
RA4Zoh8Yu1dst5FmXqwfQHcJbuaWR8urtW3rLGDhuTt7Pl6C/Shls2Ewjz4niJzFdFjeSxP+SVWZ
iF7bs/6Rid9bWMjHJqtv9LhAOneGJrjq60PkqY8ShKJBAXTP4/Bn9epX2Xs0TuXfrqEvPm3PAyFt
LloP+xL/mC2+YRU8PQWxzpiFHZ5TsWIkbgVucjxtlkuJLRtkjaAWVtsN2I264KzHHaN6lVTbQL2F
w2gjiR0Bq9kR6o50FqM4je6pQQQPKbF2IHspnMbYZBvPO9sUXMD+vTWHvLxUxr66yNq3gGhNxsAg
Tj+mB4QQzksFHwO9xQoaqSZzw4F14t21GE+vAqSa8QQfxBxnMsUzttUcuDB1wcKC3Bdm4lk6KX9a
HwDv2iWZcV1KzUq770tqvymoKHgr0dGW+KKm1VSFIKQWrlSqRQOua3cDltIX9bAOEXhKw3Mc/0Nb
jSHd8avIeX/g1W9x6y/WIjHkxQ7ECIErwHM8V42jr917AqxjgCRn8VK8UrDFMNjMiE8/5d/3dxwD
2aqKaEVWmOQFZWsfCeXq76qYKxO6nsRGeYqr224TkZPvApC/ChQ/WXbQ65N75j9p1yoEzcyfRQNd
fKwQ0uN0mp3jf4z2wgb5gYkVhugZKylxGegGUA1f/0aj5jgewRICb/hWr97fxfMha5DFmMFXfy4o
WTlqV0RJ/99h0ocvmSAoEgcC9hKt4ZMbS9antGiwtlATg1L6MUSeM1Zi9QxkdIyZq4juYwkZjRMS
Qb/d0OdCutucEWfyoci9asDTv3Q3E+Mv5341Az37ABpw+DMpEEs4SI7dkeGiTxGLzJPQLzbZU4I2
rz7M0Bg66lJ5BYJdXi5HXqzRH7V9nGmkDsMH6PQASKc3hokwuQ0EGRSY/M/ueZgUErVhMPokMfF+
e5r6otwEharseW0pE1pfaBWztMoF7BV9KyGlEPZ/LYsmCHqoxRKiCx41qqb3wPJ9f1WYRU8QPqME
Y4mun9Z28Tw9KFdOuva3QSPIpWuIMMl7+P+LS85dkXUGdYpRr2DsIkyjcx/x80O7ua/DVzaemBwE
eEbUBsJuZiNeg1By022JkQfOVdXfMmGXeaOBknWurTBjDU00hBmA6uL4cdnXhR3jEyTCXLHJ3H9c
Z1npEoiLNTpZEfSqR+CeTAY2FylNsGFuR5oMjvveSA8sZEXuKtE+3iOZI082O++hVnMLX02mU7Qv
lDbUlr0Qx1OuXPfZ/l9zaWtHbj2EkLtl7Kg8kb5Mvz8VMAvX0EXUNODgz/QmJ0SU7STXKOTeJC3P
fhxnoQCeKiwxWlllQJ75x9AVRYEujw/TPHrkhxcVsv2u/RQ2WGf75axrItbtY5qoBcJfQklp1I7E
S/URz2ok6EczohJ92mhMs3aQHgCj2hp7jDT6q74kTUCjSYiBdUyQiDoXWB+J2JOBGKUNuVVrcBvS
jIWo8B9z6aedeR6V81knq0yREEcgXj5wCp6l93EIF0KZ+sWGO0gIMY0w0w6//yOoMgp3u+sZfnzT
dsw8VfGf8q/ISa0q3fRiKKe+2GSHXXLA655pLn9GRYQpZPLtvYDStQVpjpHOc8p1O+24uA9vCjf8
RdL7wOYd3pQnKhB4EFfiVhte2mZyT3v5KNhrlBvN/Xl1S3plFVxtzc4cLi/gRf9/j1xBzfENII+Q
wIfZyBY+1UNsU8dOeX5t+nayiH1gwbygYkYv4UH/aYbtx6qqRFpiivZzDAdtcVmPgH/Nkoz9IBl8
HzmQ2je9UcrhRzn4iIQLBoi+ZXPIrk6Gn/6cdSDROSTVtwRawvYcsveOPIOJWFP20sS18sveLK0u
fAJUbPsR0M662/spYgPE9NCaR7HnGTfFS3qgP2IQ6SgcJTcZ7cQYSBdHK9eWWGly5JRmlfY8vwwm
3sdCVu11N5RDgF8kq7bHE4C2rbIu+I1X8sig26Ab7rLUo1FdBt66QjNQvgBn96FTyPz3IzVbQXKw
i9veIchACbUZ+kNpT+OTQBUtuGRxhJTHSchuiTckalzioXcDYCcd0VcYBsEfRaoPAz8AjLa1WVQI
gdxe7SBeFWFZ5xt4n10AkzPlVsjbcLIy6/LtkwZqiE9DVQLX5CC9Lt3XH9bNBF0Pm9sclZpmuFKz
cM3rAp7heLcf18gsy4iBZhg/SDrX2X8UHzixRgBLP7mm+NDddUKIs1Jr92DSOz39CEcPpv+qb+x6
VpJpz52SAdux6/aKbq0o1mox+AnJF04P46sgLh6/HLyLKUYG0c5joVAsFgEzA6KCFX0grFQ818Kz
I4uZc89mMlfLVmBG0W2EJrmNVmAYM+HwIGhyUVRUAbH7CLmzC/a+K38SdacAiOFwhK6VFIFnkYWE
EoqrdOd0Exp0ipvy7/gaDD22fX9oNLGkJhl/rbNezh+U5c4ywqvtJktFeEopfzlrHsvsv3lmFyzU
yPkectHJfVK8D5kHaQLWvTaMxLXAL56KMHWuvRxn6pkfgxmPHIN8+W27EAkVhgnka1fd5N00I8Q1
5+/XCNKYhNUAg9sZCVHBsj3FM2tS6t1l2SAOEBMokviNHgvfnxZGe/TR6Jdialk9xTZTwwUFlVzf
vMKYz25M0aZ+agAHZXvS+782JpyaVuywggD9r7vWvViCgBw7a00hzGVf7HdggR1AZhZ8pUAtC61d
VMBdXVnna2qpK10grIQPzRyh+4IskuayrgbinJHr5GNLWrcponPOZ0Sb25XQkCZY8mZljpQRbgp2
+sY/4tPaEy3Mj7K8KqKIJ2Eoa3wdY8vyxcR/Ho6PDodVNktdt20SAXQEs36hUyH01G0bdrkZOhyC
+QW/1SHD3EWctwGoSIpKn/q4H1ZkTScthSi4TR9wCccuBjU8/Vp77IIUg2qnqvB/ApW+JSX9Jnzl
zE+FOjRW4ivzqTxy0KAiEGMFPE23z3ZVyH+mLQucSyXFaVxVepiQTBvABDNHB7caGr+TbEm9WYVa
Xu/1rQF3SsBpIbYMb6HUd+cTaaJFhqkchP18c0DB1SzvW4leeyOwDvbUeBeih8KONP/hCcAsWu0O
AK2K4WmUbCZ2ajtTRwdS56Up12mizOI7t51T4LneOlK5ukI16iHXmlUNzLr/VjYb8YIFyeykwQ+I
tIRidq0kVEh7Q8sby5yN30hmVWfK+otNIy/XNI8UqZ5WN8kkqaQnNGj9oR9GTWDyqIua63cDw13Q
bwfLQ7X8PrfmNJJX4ak11MFnnwGUMtGZQp91lfWxQgs3Ms49jn0UItpXiN4/QhvhylEwM3HVtPOI
DJHM2uoArcwA87bX66DBr5BX6RqKDRlHqqbTHm87STAry47JZdBZ/xWXqruRWxQ8hc5BBCNo1gBg
OREQc8gF/S6gwOheuZT60xiR40qx+GyE8cFsF3pO6SdJgBKtrj/M/HZXAtBT+Yzl+tFNWuZ2sV1N
NVbf7lG7Fcgb206JgeNTosxShgQZw6HT/ptGbDpBlpEMgb1x4s3PU/ZFWy1Nt7eRsNi07vEJxkrT
JxhJUwtLb4/McA8Y7pFiHzOQJkA2FU6RsKDW02rawc2Z/Qf1dKmo9OaNL3EiEmw3og/hNagWSOkk
s48Oybn8TreqaCv1Gvbt7XeDx/ly9l+3nnJZejt3maeWS/+o3FpUezeRLX24MBMfk/OXSmLZNbfC
h5b4AbhkfIZL1E0MK+LV9aeYnqlgLy012PRT7cekE3yWrZX+p55cjMnbDJ9Dqe3JhKORk+npTXLs
W6ZeVjpX8El553xyNIIKoyU1+0tltYzj0r3z1GSVS8usUY7Yfn2LMtAjVc/Yw8lyrLAaCKZiWDGd
K9kh5CBJbDUKHL4osNOLppVqW3bIE862WOe7uY6mK8+lQFSYKG93YfZmBkmodOFbD7um3pNpZM1o
jjCRqTOp8FJ25AeY3Y8xCY8Jfa7WH8e/8gmXJmDhcRfNb4A5WeHWh7yCzHhy7IRGFzrnTlV3+i5v
LNhBTOSrSmXV7IOhrPMYTiAsKNQQtVYRIbFL2Z269Q9j7blPv2YEe0Dhib4z3z6AXPDWcp75PYsr
E2DPATVA1r/ylpc2wYRbRhFDCRzTFC82yeOEhawTNwCr1jCJGYDemKvs/mnSmTpzutSr4mpH80j2
fRz0pZ2BLVE5DJNam2A7EolHTtwrjJYIsI2u8BbRSjLcrRykxZiD5aBcN+IcFqoNv2okGA4gTMQg
DsU5UYAaS0ArkiVtxLoJscj7s0RSUJDMpy0aatvzVlYy29k9gNjsSiP+DjHPPQXMY1A2UHVi20fH
PLZNgCOeOsrQ/7kXTNmnUxYvOpjqUJBchwb/yCcISvB6qU5KKx+wJxJIzWeZdDZAiCDnKsW4mZot
34pHCOsvotPVc15FWu2im60vWN4RKsssqrQVXDOT66V02EHPzrkIL5mrIKdZT58MEdBIZGUoiNEJ
tahRLGoQ1wohqDxpk8p+DKBM/jUMfvKiETKESNMU/6g7dnjPIbtCdEsYCUBKROSi12AoiEcyrbig
MYEFremvWTDcV6IhWEUiNqKgArsw8e67uoAc25PkuBSskUc4oabhA/cF+tFzu0KOOKaoMy9dhDix
cJPhxRrLd3g+iUtJw1QTQuWbcbtfW53JNTepeyvu/C56rcXHFrcSsEHchKHGlgLORZXu8iAjhQ7l
zW7eRSk3Ad6hD6Obu2ftv0SC8CeGn4SQzbwjoZrUC7I7bS5aotgojHtnqIS2LVqSm25p2g7xs4ld
/AbUzo160hzY7u6g1o/mY2mcGWh4EQA1x1K4OYuko1IIAhVfZ9SA+pYE+4ALqO9GNY/XKeeCAR96
S/Gl9QGjy6ByodJHhCvYB4IceovB9WlviFSyOr2VbvTAZ0DWHZIHHvFQLRu4Srhb5huTwQBY01H+
W8g2SktNYTEpLAggrOdVzHEi5ULNPkZaDdqsSBi6aVY22i8evxVBFF1SIc/6lP5uGJa7cT/s4Zee
hsM2OAVnXicuOAEtichlUJFXf1WGHu2DggKHnqjSnkRgS9T+v50HVopohHKKb5/rA1QcETruD9MJ
w46Tk4vkSrfG/BG4HzSbWN3hfhacEwaTBWNs+bgU1CKA/4Tx1CooSuXfru+OfxGfXoaa9N4HJ0h3
llX8haESF9UDJ0vMhfwHytCkDXK6n/QCDCxODEK68ahZ04/i5M/5Nv0IlhwWJjLju68IsKIVc651
Ro3gH0QFEmUjvg7j+8JlUvdyql+mdHL3uJE6Kkw/lMKLdQY9HlTb6KVi/JPt0YO4gBm23abpX1zV
nouPB9OhaczrvfjZbDkp6DB8UODJgS/dug+shWLlT6TGvcIfdPZ+OBhX8kKWunPg1eXa0QiM+iAr
/gfsuAHIO/4tr+prbAmvptPW6WeaDTb5OL2oYS8tddlQ0WqUoF+Z1GhUYdPXqGd24Yhz4rIZHme1
9MF42l9pabCWTW9TqxuE/SAiREOlc4Pzg/4aZrZ2Jzf8hueLznIsi8n4EYTqlfdR8ehfOGBOeS5o
biGU1x13fFmr79iC9xkrF69SlL3AGksvGQm23IWgWi7S9G/VAIHbqWqLwKxxicwb4Vc/+SMuT07l
Tand33LZvTWFD02ADByaPFF5v+p6YJz8Us7xIy47pLxZdBmVNKpkCbjRcewv08NH6FT/XM9VLAFR
8/3wpbJzFMe9cnxQ1HbYnJMydrjzcrejRanbHflnvwZnxSgj991lpt9voXXxHFP1yBlSUzSiZ7bi
daUyiINaGnDjR/rz2cXxgug32H3DkIEZzDt+I+sUApzDiH5MTeKGckPyvTbMHZYJzpWnMXSNTzV9
g+5j+4YmKXQlD7j/YyURfAFrqfJT/ZHCGpX8qtuQ0nwWTO06MJaScTFk8suWxo3kCuMWAE5zJWyM
ICrtPdEzxmmGuUXHMVf6TB/MJwIOpX0INBvluugDDMzgfCfpCCs8NtHgC7sz7OR7aCd52s6imuNm
tIzLAUg8U1dZQzCQSgn6T1X3dkza+YVXDi0O61Pwzk3rRiTX5ILQKC+b6RxXlC3ogcFh+hhEAx3o
umk/vs4oPUHJ5xhNcBHPDS4pFiAh3hlQhY6SnlGqNVDNyXXmHWZCUXw3i6ldTfB+oG0KaoRQnhd1
iHvew557wUPkCq+lFlfqocSTCxj+vfBZEi529VX+8LNDBnRrsyu9B1aTWrWd3fgjsOCV0tedsmVm
INGCwEB440p7KFfp5305brrMorxS7Fct1VlsUrMfab6V/FDRJDJrRqziqe5KIj0fgYspJdeKbvkh
JNeNp0REG4s+8q7n8wbmEjPs46TuMAcwPvxKaZM15tk6JKs1Jx+0jhnmDuW+Y64btmYPkytIbCYa
ztIHRgoKxFylm1Ytk6VG1fQDPU064ip9UevXADnMzqal6xoUOpG5IPIp/LvBM4iZqtfgUb9xaTmc
nesJivxrG8N1ZCZ89u3Ycp3RrkOym3HFn77/nWrmuONvazVEYxWm9E5lnErQ4bFmZ2LDgJUx6qQ4
p4uK+DC7xHTnmPOFk6sKmQFDWi8eaOsA7j2xgkncs8uA/KmFgMF516OA7hF7zcPtaR43uYT/2dm/
lyFdgDJuVh3MVQMfXQ97OWbMnA/mANt3+RH1BVsDI+5EWgYy+uGKE7vyDmTqDevn7SYBPkwy5FUz
p6VeT/Vet3W89q22uZifuB/eEhP9KDl1XcFoYmJ37Ntd/mijnTyKzaaC5cbQTg87J1HyByc6LslQ
dkjUx46JuwOoJaw02BNoyRg46vfOPlwkEcDdy9IVfk8RMxz7YjbyjiAD8OKO/TsxU+pTGLRQP7Fw
DX/t+8Pp3gRlFqO4E9UqNtTomz3T5cuDqWSfpvmfQEF7l2f0YbY9yHmgu0KAsUeWOsdtOTnFeibI
pXWSSxDgSynflagroqa9l0habybUGOaafUABIYD/9ZPTu9oVnMwrgXIDaiuSvPZ1PQUsfrWGLvOg
ahy+vuvOb75aKiHDOqJHQ9ZsxYhBeZi7S5ef4Ie/xIzNiVzVMoFcfCjUYRKVf+VlqBVnjhMiBHdu
q6ANt4hogTaSrLXYyHrGBrxyIR9eyTPVdYJoWNFEJTSM/Z2lOg0SFX59FFLGtaaIUatZtc/eqX+F
NSGug4LH0s0bzT26AoLsWc/57lupuyYND9rAQ/kqyk+GFSXRmz1BwrVg6Ml/f8//lq5Q9wIKOMYC
Vm14vXetWLcmuVKsGkgD7PiSFVTxWoh621Vb9eD6LUcKOeMbQlJOWzLgb1HSQA0hvaq5FBJMeQ5h
vC71tcwHKivzI0VVC1ge5XJ5SNv5LDe+4K2tnTJmwYKsZwW4gBwVzIYQPwfut3HwD6309jshatyX
t1CBkPqaxjNDRJKcY0R2VN3vSXX4K6cBR5zcQDW57Wh/p2r+3HNRp2pIg6vr70u0DqB8Mue81VlQ
Uv/VDzgPpOk9sEyFjqYsHgX5GUEFMhLKgrvpGmz14ZapOcsbeDCwHfm5FYoNNHokr3efMlDK0O9w
6HMhR98w8N76GV5A7eh3X1Ncpw5Fa4H9JM7MIs6k/aON+5hnVmhtoSaa9tfrQLxJIZnCnwKvcVf7
AQwJqKF4iCy0LpN4LH7n+yrSSx1CNmmgbALxELlu2WS38GPItOFrZfO2P0MTYzxq3OfFF8DXVwB3
KaP4W4E4My2sJKoOA1qiUQxULvIv+UMBAavuoSq/S3vAWUuWvqFC7qwMtl/odw48kW8JbcfaMw9Q
fa+k7q4Hrj/HoDWO8wmyAn9S+HvSCAom7q8AfJx9Zywq8XGeKjuyrDRr2AnvhQruZuFs8JMzFqtf
jrrWTmhMbOJQu87OBpbHifi3xUNQMK+zEKh3VD2gfLuAXT73B6xE2NBG67mcMYDD8psSSzURYipx
UUDYW2r4fZdDyngXlcJLo0bRFrNVZVJm4mxnDqGyLvhoKo+ILGf08rkjyCfCYvgpdY8xVPRecGuw
Mb0NHDK8pfdmw84fiQ03WvvnsGPkZn0wPhqt7VHfyHMwySmH8fVIHI9uUqEoLXpFM2/lEFo38o7f
GqqQDiT/XTQ+qztNKbeL7vcNODAW0ZSvC1DgD9+LvwTAgiGwJqOWxMjY4AbGfaIX8/X/msSq1CUx
27foA/AwunhL1WBdbk4O3uqRxqlfTlGfyjZ/QM3cJ/OYQKYcG+qQfbV+UAn7UZ5nj2zeF+ndN+jC
fw4zcGhEfXhl80wgc+IqcpyRromzvTsYjOSLIi1h54GFP6vpRvchEoXppcz1UxhBakLbd1pKmd7Q
V4xqmWHaiIXgvMigv/AAbHIzUYpGa0J/+nRtsqOnUI9LxPuLfNJR2S5FnQqTojGvPXaM8TBVXNwz
wc4ISuAek135Q+obtyfYm3Et5pcFvgpvvTEeA1v5naGj4wRG1QJ1aR0hzZik+g0pGjNxneksgDoV
unzhnkKbficSqZfoql8seD/6rElCGrqeIbSa4IRADD74t+7VJEm/u2bMegk+UL05Km439xceB+3j
5MsSnAuMLeuizMB1lyy7noOFyjIQDJyzE3KeLxONhYznU8jFbrPW+jTbhUdrTgt6fewTb9pIWjuF
J1SeJw7XCaLc33r3i5RNVv8ete8s7JdVxIzDszBgSpAzukPs8UmFyo8Peu/hr7T9nRXPSNc0fgwn
QCygy0yP6mSTM96qm6DeC8eLS8eRHIvqa7mSt57A9XPs+xA8cp33ytAQLf/W1WskunAlQDFAJYMg
1rNm1OuzF8BMlLlT7d2mhv5Y3ToZdsOeb4MfQuBEjP3sSSIcA02+R0ECVfo6E2XnmORlJO/REXzg
YkTM8F0yhWAwcsOoH9xAydXSfXIe9r+8C6T3wbDJWB3cDEzwpysmsH1V6L4c9VJ2JKaHVB6jy/ja
tDNsU0MBNnCkK27o4Yv9smX8A+DNLVewMlZmdDoiZcGHnR2ZIzqkGBLiNDi1Dz+Ni81p9YgQ1Zzd
cqTmLHCP/kl13ioNKPoCtup6/Jaccco2dPw8Khlsl/XfZrHf099icsfhAfknhbHCf5ZlzQIEodcP
TheBhCMJEr/eaAXJKpss+4PsqoFgSJMYvmtD88CdssL61Zfx3JQe1SeWe3TMXmxbd9XIUeKFn5K2
l8uQ/PBc1tyemy4oTp3ka3yz5ucZiBmAkhZJO+6q7tRdleMJyvtBK0ZaSJjGFmr4iwrJc0oxH1EJ
KnmNlNa0CQDy707HpCMj7/9azruYxJ2CAgQV4cL5oGYaUHJLq1kZPFkZguAQ79BeayNvRaEFtTbj
/gjrL1UqbSjt0KnrGnJfEGJR3zM7zUC2WJ1mD/y2nhHEN9nLlIAXFuvw0QmSN6lYxWS6bBdADOXC
DWQ8MotxI/Ez8aillR7mwsK9VvkBN4zE/HTxnJBgjoMMgiQo50B9bvn+4lUKg8Yg+RNXsMVzjSJV
+UVQksV6qeK22zhDbIiMGSJs66hccEaKI26PDGqHNKGX9IRAHLWKmdru7R4enUtVxsd6a2HrDGwv
BwQaSsoJau0ycjwYQ6ANisYHUOcwbiRhSexZkwuV3NHON8mh38/xDfsVe3eB/9N2S6JVr7EO7U5h
+esbivUBPhwk1lq3sqVykXBndXtbUq8MXh+wW6kFYKIiN3p3q5MxxEFZBtPGu2Q45FZgfjdbG4ff
i1UBOKZzrrmaaz4MpMMK0nrPsFge8mtaVWgbtBDNlJS2uCDbJvoW2VYEHSn/gUOu/xAI/6WZ++nN
J646miVwvahl6DAIRzeBFXlNFfwZOqHBzXTGZa+7LVap+iyoX8t4FNz6JfFrdYRmmGyRXZ3h8uhX
S7UYuBFKV2ChjDss9UlumFXpvcR1/eP0y9/a4sUAA1YUijfBW97jbVuJu5SO31fzkxVNhXrFzuBu
4ky8xULQMubIRggnFn83wOYR85+yfPLtNElTXvMq4PsLbTYERI/xhHjBMC0wiqA0L/nQmZm2NWwc
13pvJ2vl1aQy/HQXb6KcRFHTCUVo0P2nCIk/hmocNkzyai44bnxdub2zlP2h2Q+xirZ48+aGk3So
yLcFOcylUs+omjDIKH6ZVBCiQ0DKpHg3ihTNQSxEbB4ORRu7q1GbjDt0f1wcCjJjeEjYP8zwRGtD
7KuFPt5pC91Z/Hp3fXgqJA7XyLjRzcTahPln8DkFk+r7ojoUUrw6n5jPeAkMbB63dBIIjVmLyHw1
rLwSrHKgeXAudzXIb2jia9wGI+W+K6gPZhU1blP5s2NIiDNFSK74ol89M2DhKiDo4Qc3oK5OXzW2
vYt34FOnXC+5te9jdLwiWKqlJN/8mDhmEhThuHI8b7k5yHnK1royKV9wXAHQfZQeQP3QlRE+CBoN
o/zfPkx1B1Dh0DDuNJrFTH7p7nFxtGp4axfb+wpT4I/K0oQNLZECzusywf1ojbkg+sl4aoXSfh9u
yP98KlDuA9mbGY1AWq8h51d/heYISzxfT1WFDKKA1/GpIHcj+qxtVxOMNpJOrurGiO4Bo4AB08nt
q/vGwgHefGHG3yU5B+Wzff3TsrqRQaHcQhAffeCeJ9DTigA8S1Uj5N8B54Cc3d5mfxhub1yxs2N4
NLfzQ/yu+jrc4w72/lR+5+IkjLbE1WXSlbEPJgqeQKH+XHwGTlM2ibcu1f5roVW3Crl5aVmAQ30I
TtUC+rb7c+2HLvijr6vN72TaufHSX8CD1SpBYnNo7BcFqgR9KKhC1rAJdnFfym6xypo/2HflNmmQ
H13mMQZYvok5nKUampCMfUzYJ4GOxyRmEvOgGC2Ev9v5UBqCSsAXLiqhuGxJTCeoF84vHsfv+2QY
hVDW3UXGhCvCKAZGA2FJnGqEX+6ntcLPwB6xOzrAmbzxNp1/hRro64WIMsYZiVuy+1BNz7qHyiDY
F+442b6I8WHyX5ocyB3o567yLq71b2sGsJgZBCRTcuqmQWEA0KIDM0N+cuEV0r4ek/gZr9LQHXuQ
EjHcTONwYLL2z69ZL+rqdPnwZDJ9EmXDvxRqbXhrjarsQPirQMAxMVhMzzscNNMeO5RbrJ0kP4VW
/IxC+eRBDkinz+mie4+bdM9xab2Igd28JNa5hQh27rmftKfUaS/HftQs8icfwN0bJoLK2a0eUXwP
Fm+tkSEd+oFw1XTIPx3zDI1qkT/0PVly9tN09QA4py7Yu10bTk5yvAMvyzOoJ3dowk4m8eoFilaq
cX8hz/js/bI1fy7QmkoML910GD7uUSdDUfwtiAVt8qcfK10mTfWwD0+pUj6RawW8UJwlB6+38Qom
flCT5vKhK4O1Fbj50azYU7Le8aU0+1n8+0a0awKH4+17oVsrFtnzkeSaj5zFZE5p7UX4xnkOrezv
g89DjOZesdh33dSATL1puIG4joBD2OGKTSu5KbE4zLUEAeycu518W/fnNoiH5xWw4994LTdWwz+Q
xyu3M2czlIky/jBl4Cvo1PNLzpWtaEf5om/OS8N852gz4YEgbyzp6RDXe8CK37eflzF3qKpptW0o
m3CEKQpLlPCLY5XL9nGef3OmVTwUUvcV7wkRZVyK8oTduRQyTgtyo4ixjQWkxHfUgNaw6zY6LiP1
Pcx1cn9k/I5aIHBPCRtMGWawgX0ZZMrCvrHa/E5EKzS35XSQgIAZfbtFhk7bgeNqx39jmJWhil4e
2t/lnmIbBp2NoDi5fkDNvBzPBTmGqFTHZyg/WNs7C+O2seWY8CwOkIYpyixREK3eOsp8pVSTb7qs
fmZjOqezLZZAtEOTBvib1KJZnuJ/aVFAmjr1FUWWf9Yidag2ZRkKL5JJCJRSQABB6DL+bUq/4SBG
lahWCnveETvkwtTEUdwvZwfNguqhRW92nILuBQENw4Y4/lskW8aueda18ncuQQVZbstSYHJsAPPG
XUoZB8QvkuFPZsxRxx2kPqeWdDyH7kZ1xIUZaOnhoqG9WjccBdNOLRc2cSWbDa+mVymuoBvdPqLS
VY5xL7QRKS2vT++RTEj7hxq9zZoCDe9SrteaLzHSmaccyJdpSxAX8Bvv4dXDtgAgA21wuBq0PRAL
zZWs6kMz4TpBPqPZspwmp51PdEvYDzf6swvXUS0PLCsB1BkJEBdp+5KgLL/f5YF2QIt6dnBLHRLa
rL8hNmbGps9SJrwQItZ3jzqX8GwVBX5hV38jOFBgnX0KHLe3oJ6FX4Z0yksqZYg6/bwoEcwkr/ET
lvGtIuELJfVpbq4hdLWRcXKRQs4+uYwuyihZNEa85fnstr4up2yvkmECDPeihdPWha84wQF5MVEv
auOV5fq8wfXrOZeASrvN6s1y9WxjzDbwtj4k2ZUTYKKF25c5KWsR0k7lC8ou8X1btt3A0yRv2L2s
YDjPDWZmf8gFALRjqarwHw8jHbHljYnvwK9K3vugKehgoIPh7lFodlNFELEDR0DWRN27Gi/sLR87
N+QxwAG5S4zAdFJvA0CRdjuaxYJYSfI1Ly9PSjuFBLIOCcIu6Yf/26YDv5OAUzMmGvrb+j0qC9FB
Y7YBOCUoAkGYC4rovGgA2qER28KsLkFLgufRgeiaCJQhCd7ul+MhDL0Ej0qL084KPylwWR6321lL
FRo7hs5BGlDXUvVFXEFJu/8mOMyRKdB/KzvgOT6BAtviysQn4qHKOmLRpvMMmGYbiNcP6O2ybRSl
QhUlkVm68CkFd4udOOylmztKW7kv09IsSYlNE/udrUcmqcLl4KlZb55JoqmLW/UmTzZQmmpG8E1z
COVi11C1w2A4P8Bb7BCQ8v+a6s8U6wGxppC0nJjik7UlWqKhLkVcPCMxoiNLWddmKDibouXiW6py
K81qVhWRSEpX3FK8hhw5uB3vBJ/9gnwtpGqEgoL1mAIFsDHObdpw7UaxmTLaLUez9tOQaqNPvouH
y/I0GwH6rC9M8K9H0TUYlymUrb5/CJFgh7l9HqrbnXc3Mew6OaicvsZ0p7H2qlMdjKW2OBPVbg49
myPbdBFdwtBzL+vVQPHuqtFPibEKuvgL3mIJM0YWI9phhVKeoKFVmNWdmHsoRKRGQf1T12IZywR7
cLG5JZGqiUuKEay/fEHFS9RYUfkonOyF9ZeAhp3GvnNKf9gYmK8K1Il8w5i1E0gUmQHwPhx6isiO
fH3JW+hNOu873SHjpBhzHi6m/5OV/Hv9vL0Pru5Ofq36n6E/GIXZyqmgYoEi5OrJwlBF34Iuu68c
AZklx6OzWcOk5NrGBlTFrG9XLVt90/BoHS3z5JbmhjQCnUrp2ugcC55+bq5iOsdmDQC4fMh6KNfD
tvi4VHoxa0qhsYiJgzqXOpgt/OB6fHDwfA7wgU3ID0q8uYKnB580uslu7+VErSxQRVVUAikMDN+1
RG24Xb/HX4IxO0okOrnoIjMnxVSONJUBSwQMSJ7/3akqC3ozqGEwYLFSH1KbF6yVWdG9i8QNo29v
myqozjCyhsLEODK7vtcuYHF8Hd06XnR/f7E7RqPuA1tlG4yChEowTZDM5VfNT6OVGzPl26OZvzHe
NedCyfWP1YfaG27B7xFN1cG8LYvgtZiHE77XyZrGv866qZAGD04HLoDL44EAk4xezyKCFkHPkKH9
0/4ypHwYjmBf3tAT0DoTgRErj7/Ka/1zKv22CkGNyjGj7pnagXmZBz62J+0PMcV7n3mZSeoFiZte
d4BJZpDA6zFujgdkhG0JRIaK6JgXlswON6Dw24tLjVnkiKb2qZQ1U7dH6qtOZiogXrRcCneERJpn
jki1sMn9/YD2HiwjWvFdeFCgAgFZuWlLp9FeH3N8U36Ed4FguC7CIDHCGG3zJOnHZ1A5yJL4v2Ua
WZ3rFyz26+g5itIFzWjytwH5QG3ev3pi0ts2L/BiHnadb1J41LhzKmAl7oH+4b6l8y2f/FVQA1SF
AS4P6BhNisHK9O9eOgkCMeWOZx7mDP4sbBchKjD9D+N8KK1WfPPYIkuM6trOK1bzxeiE9e2DxG12
HMhaklm3W7tHs/9ahCIUm1Eq3PJFWJj786cc2cGqUx2Ci5e6wFQnpzLgn+PPIn3Het3L2SzKf/nN
iDi7VmntFRg7xkR10DFu58B0sKBhVlvxcvlNSNHXEuNXLzdsmMetB+GGpalMYqWG1vzrfUu6D4o7
G6rMTmeSkykwGXksvmueP+JGIlZ67Hg61jR9bCIwrbx9GIqao/8rZw/SWcHtlg5uQm2oPDyRgZ6e
8YJAmwkqqZVgpeTB67SBdV8mESuujGkvfMIrASUCCICs03BPWDBkifqiGarzhwUvcsHbj5t/Nk7f
Umo2J3gOOnVWZ3HmW4M8rUmOg5gQzUzokuH/Jm4B6M0/9KjMIPJapaPLPhtA0cLKiQxffE3/3Poo
ukPFVCnpLarkQQZyaROAHnEtP5IA/wVLOQ/eCb3OSVNtSROEM2qJPpG5V0o6bwDFEJR/Vkw6fA7+
ly4FZx/g2McAkH560MpnSAOItuxj2gKbhpeJvutBg32rLTWx5sCzfm2b9CXUcjTWQOWiYWayLnsl
qKhSm3ftGOb1Gwzibk8GCHMFYXoHxvlRkJIZJ2ju1/50A6/qszHdLBlVcSeian9cteQnvjrP/qXx
XlVYQ+wGCx95xg3fEChnXpRek3PFCnvkAprB1Y6exSHe8AAhH/HrgEj08D3rWGXLpEcLT41gSaES
hAN5lNJB3sZm+M7TbYGL+KplpxmUpjmuSGCvARwL5Ld3s6M2luYd1yrJSALnU+GOucpORFXeyO8V
VYZsR//wlIPS85QHs3oFH01FPvA3MC+cxdkZuCFIJVckmWBOTVMgzRNMcc40jfU101YYr5dkYBaL
Lnlra9752J7AkuoA+sXAynHF36u/2Nds7UgzRiEXZtxfdHxrop+ARBUEhY8caw3hK5dStOqVVHMb
WMOpTAmNvXFd4ns9tOErxkZAg5eQppEkKWt0bcE14nEOGa+gifacBk6Ypx9EIcaIzEFlf3H3dbOz
AIwz035BnkAJvyGj/NSUFcMryEO/98MOnggqwrzlv1C/VXxABgLOzwlkz/lnmtHmcvOoBD9dsv8g
ZnQnDdkBMxmakSdcPdd64SHxUttfetD48bXyi2JSAD97hdU5q/Em/jXBKmFtdDyTkTT4vL65rvEy
cH5NjDjZZr9vsuClyCzkABjYjhStg+T+JXBGW9SywGiR3r8bXP/uVuEw+Gxs0UKvJmQRE333YE0S
BFkVzoCrRbhCUKqlpnUNyWR+XhpA8oFZfeoJS6ecQi5GxEWU+nZidJ6WVmwiBWc8lTr4B5CNtclH
62OSwQFVJntypGQ0F1oaJLayC1OpvFHxQ30uA7gpNDwSWjs7AMBGk5gWCCOMyiLBsFduWDnM83DK
aqeXflYqR3UzzfwwZqRdLZSZQN5CNfhDEy+O+8UUDO19h20NfaGrPNQW+HKEaEOx9yGfKa7jUj3I
jX9iBOCMPwRA2X17XPGNdZwDlndVXPkUC0OZzsrPPRi+t6VepEzAGcVuxpZVQpBawFcRv2r4jhCR
Rl2QlSSDI9SbRGBjvZ/t+W6hjQYjzBOp3OhldNgA82qlccKvWqlh54qFKpoXPg6L2fDIQMtWuo5V
JNS7vIW6u5BnMw0H1KRdmss4DgbnCLo/yVCadvi0tl6CpsUKdkUr7GwTzK6EPzLKlnahg+gpnjIs
RnQC6EASyTqCCBPz1Eq78e3j69c91ApVLCdhnk4u4fJ5QXi2mRllCjqugK1ExxBWox/g4kowUfST
sE5GocVkTEFKAeGQ65KqnZt8tHTiNNr2bCe3SpaV01WX/CuN22k2J1prLWACghiIBw4eidfGZgYs
8NO4HPwYZg8LTo1E0BOCOCFchC7e+0Ao0k8s4qcFDwN4mxIbOFz5W98jDbu0T3UOg8jqPnn7gTa/
5UR9j0puZJJ9Gw79jzaRCWYZ6xDoUu8O3YLmaMKZxbbSNKGP96K6la2yHGlnPu8wghvdTqmWmRf8
vrOpHnQovMN8CgTUHsvpAoBootyg4eXr8ur00g0ZEgcAffgQVsn+w7mPw5T1ib8YQ6cXx1uxWNp3
6jLp2oaogFlqOorRzC0w4EKQdTm3cW0TD3OJl2dfQGkhBVFvl63lu23f3LazxQX9LXK4h0F3z+jm
fHZUm2bZyAjf+rkIYEW9GeGK8m1B48ZGHTBvh5T2CZjagrIyXzJ36xcYyKpHynzrqaEjSRp9h/fx
40qhW4pGnCLTZTftzIROVWufIPVK5wa9AL5u4PolljiVcjIt8nkwGbkXjhv41RJ14DHTZHsNJfTA
dIZXVBFoPgx26Xhasq5vyYwZo46aHsViSC7A/nl4T2jOhzAvMDxHS7eUs9vIGrBcTQbZO5+x6prs
JbRGTr+5SV6Hb0lWreipZU3yQZ+B0yR2BexQzpCV+4uJ2bn1yIZnyy7IgQwjWJJ5O3MmhZW6n8G6
pxua9pielM0TmUVrkXMmifsc0U+d84p5u+4WZhkAyQmcjX67QQ5jcKMX/SocNdPE8pPczS55F9J3
MqkK6wQ3WJ7F7xemMpdrSIXFiqMNn7Z5PkhizzE/JwRmCqxsTBcL1JlnntosUDjpbo6hefpOW3EA
6SfXqOSsSzxHbYoSbKLSKNBXYYWXrtlnzXN3dnMLSAXUKOTbZ2V36Iwt4mRRBvS6wckd8AX+wHsR
UzS0/OKjd4VVAYyibc+3kyUP5IeTR7i56sYA7kLrY06vIQ6No5BYDheDuCSCrWd5Y19zGJcc4SfF
4qFIMsQPLzbNT1nISNINj/nl1qQ5HPLbTNGZHPGyo02EBIypCmmYx07QT2PPt5o6+MbCSVUwCrpQ
jkZnpUiiUFvx9zcdK5+DZ/NMciievywoyKjeAKa+O79PoVArjxaRryAzUqY9WLucQvdrxCHGHvS3
xopSGsA1FCqWRk6yWzYffODWqYt5n3Vhdj1ynl6B/uJxQWWaCwJKzZhjPpyfAseCvFDPNETcrSSw
agU569MSJtAijQxHw1S2/2vRF7og2ZHkeJwl3ISw3z3TmC/WA4x17XhOpblvoCn3gONm8wiTkwed
LkpJgegvkVtZAbB2eNg0q5wn2kbWvd4wd4Ks77BJ2lXb/F6Og8Y0rszIiL8F1jZNygkBEFDHuvGE
SSqIL0Gwizhb+RgzSyaG9vWga87T5yiAMAZ+LG0N2FRUJAWU24Ur1228gsy5DIiR8JaS7W4VM0wd
lujCnW09EINNWLWWQUK+Sf34LcpjDZqkAk2RM1V+ng0SPfU8zlF/ceV7MnVtwzIHswYXSiv3+9x7
Nr6TqCuUmQqYo/ERH/Yh5oYeiIdYTTQi8ck3JmTyNi/uYUqD1XQj0dlEDINvdIXzZsbfxTGWjENE
OjdgQMQAG4SvZurB/3+voxQStq5b4HajLaI0nNCmda+h38tk6oUYcEr6ro7u0FG+rcB0lyVysUCX
jsEHSaTxAqDl9ROPmO4RvQ2MXXu8sdRN77ODCqlxOsSUpAIt4mQc4CP8ghvj1ng2E+X9UGAXgYsd
EvU9ItK4ujmTT6kvVxx4pRVDNtAaXeHuDFMTnX1lF8ttrhzir50/kXVmgRLNY3vCbCT2SEuujAmX
5m+PXH1kB/9JYLrg6nMpLk71dR3XUbuK+6bX43xz359JxKWcJ+yxY9s/Er/Q7+0/7SUgfD/E3eb4
Dk/f/piXTgqrgE9CW54GwWUJNNg1Epn1vP6Fa/mH0DT+W60e3MVSgpL2JU03J/0YIcm76cx98MVw
2DF/+b0R3nfnsCoYXM1/AL+KJc73qfbC2ibdXQKXjmuvYhUULF5FTPPAmcPi/rTUio1R6xoKU0RH
6QGF2nkkRmCCmCTJ/Byo86W4kZBxtohhopwPF+Ts7hE8rZ67C7FPCulDFZp4RsX3RTzFADgrvE8x
8FOqIZyrH5IezcK7wXosu56ya0Yw6A0PagzTZWX5tA6Vs9k08uUIYh4tbS1C65i9w+5TSm1UAveG
aaviNfTGNNRjzGYTwWIT7JIFLabb710HqOE8zzYI3FLyM0eNwRXjohMEKYNEkTGaz0cLSKdAcQpm
+EhWXWDQJujvvjJfeiBqT5PheKPeAXY19tS5Iz+hB+AYB2wpa2ZUwCgAvlAjtfZIQajIGDv0wJoO
DEkwuLaMN63OE1RmEK5AoCAhxh4rayaL/UCKQLWpUYo3sGJZURlrtl9M+SJ6t/J2F4TKvdfxhICd
JMxcQ5UYDWOZpObXtzH84r96x24AcepkA3rpvV0rbCSgkLyrQqCAVCVvDq+5jyi8mYpnu9X1MYys
rx6gu4EOhEi2k/No5VW9f2mbjyCiolB+Fgh2du/k+9iHyPfS+9TzCbkYV9ICxdmOH+3BOxxoipdV
t2CcvJUp4l6W1phrdCVJsX6EpKlAe3jbF/19qH4aEG0nT7FOK9HWgV9LDReQqayxLcE5XQDASA+s
EAZ7e2X/MyVhB4f3Ib4EUkU1L6q9LG2jsR000OrDry8JN0aEttE/EQw6udtjlc0AJiTi7FySqTwb
DFUEVnauOgK7JdmXRoO6H5jaUWOvtDvheCNzudAqjUNt/8tVpyPirwmDjxhpNeZvj0CHF2CUD5SE
QTsCjE11Gd61MzTsuVZ+SFmGvjsxVC7Uzh4bj5CJqkhIkVVTUsEpHb9DWsmPIIMr6Q9wqqBICf/g
giSkUJmm7ZKgL13+uwtMnJcIu8gS4e2ZKK4unvfhdugwdnuTESXkV7HQe3xX/PSfXp8bGxy7JRNb
+809YqGFmK8Vzmnb99k2Mlo4e4INrP7v4nLLUQv6lyfHmmvnW7x2XLUrKcZc/+9SxoAC2P1H9EHD
DF3md1pR2+FMrFXpr70BZOgUNUHigWf8HiqYJ4xYwUdf4vF0ag0jGdNVpa8m8fG/LyUD8LsrXjjL
awA2TxMQXO7DRPSN/HjrKeFa2T6KrYqb5ial2x2k+f1dAnF8hJUH4jzzpZjL0SBqVLAcoKahLJws
LoewjB8R4vqN3H6TRslhJzglcM1W6rvzoL4okZR8yW2c5PGLnMy0NSEtVSvjVAIwlhNEME6UuKxE
lTDf6Sp8iuvQYJ6tszPCut4xhDMJuLKMN9pgVGi3CJv4IIsinSPCw4jbVAmqxxUNGMAS+cEpdWRR
qU/hHsy3IF9I0U9hdikK3kSJGVFG6PIALU4HkzqnfNn/mbXDAM8K8eHSpq46nFNz0FnWusOxlvzA
NWo66vc0GOKok8poIam8bunnfJ3kUOP7n/4CgZNueD2N0DFzHRY6QKcxvZCx4jTFmyE78aEVYLBu
1vJj9j3yQjaiEuQBK1G9LZeZRP3PgrwmRehnkHVZvC7QdulUjM0myIBHPHLZYE4NaCcdbU2tEa+m
dfYzQAedRtRHX/RBRWBfkyi1ZU7nDuwR/Nhg9COpqchh1zgdeqMG/D+xmrXpLHw/RU+IHTkDXNTX
4ffYzPRhitcYWHAAA0/27aUv/YwJTO8pIJ4yGPDX103EbEq6ELWcRUFcoUVvSoEN/NpQZRxhFG/K
Owv8azZgTfnD/+lj4ntVYCbBe4TxBHYh80LiVkBPTp44LlQxTaiqyDwOKNjhHjdJ4IAozZTdUR4W
fHM1dseUERKNOW8bbsPQSyi0kc7Nr0hWRRO8i2qD8HtvbB2VyfeVdC6EcWi8A7VYGyKmPaGNIUTD
sB8IxwF6GYlQpJUnkhSEZZlGM0xJSmLEo/eo1l+3CyqPgeqfL6hdyMYOE1NWyxWPYg5G4zEgXvhb
he4DgwqQLTz3e+8NVy1NXe+hx8lK4zpa6BrdUmQAeVs0PcMLF2aulQdJIzY5yqiBW0VGhPEEFvTr
PeAfBUZt51WgfLkOEmDkptCNfbdfXc5eEcO9Da/K6SBDEfol1cZVL63eVRIi6Fx6Ux6k4PYD2VcV
uMMMIIwvbZy/Atkx4vEgA/f+bBy03Z0KvAXsLreG1VGZ/dlZtt05t00w3doY5aWTn2Jj+2XWdhfU
kW4+Yv5vheqoc8AW8Xq0vMU8XVWNPGwqskxZvmfzGFec6ow8TIeXKCxm3kLcgRPY9DaQtaALE2ns
gssWsQdJyykCBKEcLXGm/L6eZVxmr13faaD26c1ATw5IK5DPZPasqO3UMZrEiB8N9k7R4/dMJnGf
kBdGm814qPS4pKOjzIJh26qsrF3Xz5kd4sEOCTYP3jh2hrEF72mdLexP4T4tIEsjU80bSh+r/DCX
2j9EXJNnTdE0rpOGxscLgPQHpo1e5CO+sZVETY17NeTpoWg1GZMOzuCk6bfwU0xqKXffvpHQ4/2n
vXy7yMH1jELREsBuYxgK0yEXpeza0nK+HgmYEMVKNfk+6cJAKlV0c0Ifv5VVhmKqpn8wyKV99kvJ
IgjQsRUBcCaAQS3YsER1G3tupGU4RJA5AHGVmNnvjJpHLSKGOXj8+sjP+YcsYJmFyNJI3OYo499l
kgYWjnQ9XVJVB7/GQ+q/+RZrfMgAJtkrU2aklRTTPA/4Um3upu0qE5bFCrjHJ1QdTxL2xipoGcke
F23qg7qDPYw3YL3fO8MJ/H0xGNcB98Mmdh1Zl3IlrbiXHxX+HwYPtLYgD3tGm4FB+FHC1cJ0MiTy
/s2DNaz7+IdO27scTE3SeHm3xJNm6nn0ySs/fstdHvFXej7rpujAEbHSe7TxGww6ylD/1v103My1
HsP4n99FAC2+EpWYDaJ7Wv4aDbO2tBx059aTjhfFdHI6gxWPsv+R+hqNwI7u2BPY0dqCUA91kJq2
S4YRD2MTejVXFHWWLc0cNFqORC2bMvRFWxbXTaXCDbqJ9BG1MCQKgVOSv/zrELMNPMHvmVBQG36F
ae6qs4zs8udEaHrfD0NK/iFFAmlWWqU9j8s0Dr1yAEzgXGGX09ZygNKZxLv6K4syfVYXE8bPKyl2
1w05/lPeJSgodMnG+d/PyL7RQw5AoCZI2fVeGBtz2kpj5Me/QESrHRbZ6FAhkx76nSbk2NcJ//nw
tG81JmdzoU9IxbNZtaXrj2lYZ6n7k4Ob8uyC2Nf1TdVJdGcP/MKOROG/uBlmQ4A4I0BkeaWpEhOf
+eaoU6eG8C7UCHlex+kTZAgHrAhFecgs3zKa4lfaxlDFAxelwCuAdRem+cNVlH32/ml5iPazTU0M
PBhklTAXeK2dvWfHBES27GNYfZiEXg5bMJg4JykBsFR9FcAT/m7bxSR4WHwmvNj5Evi9yRXHytp+
AdKxeRlffhJeNZ3zhN2ye5Z6xywLqz+cyjkl+P+xlFVZ9XsmW5VP7vi9O+BGcjQBJSxgEVBVSfnG
0UPCYs2owCDhy+bydsCo3GHcPQR6PqqmbZZD8Op4Blz2HPUvCfbuW5FfinISj6qQSJKv8U3m0cHr
gZprSNoR0MZsRlDvkXezuVhcPLEwUQL7u1lGsn+VRcC9Wr+s+sQL2mO4DEB4KjRmhD+JR/ahiMbG
xYIpj1EMZuxMrkFaqIyEpY8wB8dQ6mnmFygvUl3rK5Pn3jBLagKy+NGbhqUtclcLBk49nDH9Racf
5Blbxc5bPyDsxoN4/yFjNRFycU/9o8DKVKmQYhqWYHe6vL4lTADD9InMUIlBgYZ5ooLROdwdjjkt
jJiljWmFDCHE8Bq0kqsdPT+iKAZ5it04F5eocIFhGxj+UpwRrrqF4c4pBEN3GvT0t9IDWIZozcTP
rASP0JYnQ4BxWpEJ4B5oLV2UJuabNR5jzDlo43zmZ67xjrb46tMQG6XCxfP9XY3GLDOxYmr1ZC2S
04zfCv52B2312qk/mLxq0TE0y9DoytqA9xCDV8UIxGrXqREfiNScuO0+NCunfwstwKrdBzFQBkc1
mUY5+cpWngh+OQn5+v3OhMEYITb4RJkQKsWzLeaUQ6xwOtDZVIWOTrUx84XmB1PRLjvLRTXkF56k
hNeYXWnZXaI7kNDERnLT7f83Fly4I9EGx6eH2s8ON1yUjDlta/T+HgKUOf9W5EjS2Nvtg2bOHhg1
Hlve8x1stmdZypLi/PodloEvJXupy94c4RuqAhL+kaOHl2JyWwj7KA62r3/6l20ayFV3wNoA1Mv4
WcmTCfIzjYrbI1JHhzlYTI89tqJoIoyWrXkZpuTlXgK+qyz3Aj7G5x/sSxNDRzuPci4m2YB/4kLi
qEm5EYW4K+xKzh9KxVqhzGTC7G/jYFhM3q9VrT4Kbt7L1j3xUPNy1+vDzhrIiHG+O3LWyyqobAxf
zcA2eJ5g4O500fgBiITLXoAzb0mcgHzzz1y8NJwlFWgxyOY27uEZjhLwgv0ScnLMR46y7tDwN4Ob
HbJ9fUrX3iDEypZl2/L4BO73jpCaq0IFVXtlcF1pZ8W6u7S+VXPkFp9qIJk/rQfoqgR4KPP5bBUq
kHrXm+HqPBnPPiIDizz/7+UrssnTFa1UVduc9XwODbFbUnM2fGiaWxdcZ6KnC3cXSejIMR1AuaFa
ZbJMQ05NGDNoKJcFNPctvdS7tcJl+aX/sXtQkq3eFjSLe4GWpI1X51bLPsvhhFgK1Clb5MNvfcpS
eVPEGgiQYFQL1FG+xj16SB3TXNLYAbVFJcvxrrM4oyyK93hDgg+/NXfP+GyCQ+1XvGwXbU7lNuuc
6PRWHRttpcxrmyvJxRai1ajYwa2oE2UOz28tj4fRtQD2w+8AsScY+YgP+R3y19wtFPBmjUClXhXA
hjkV5Tc3xVHNfQSzIoIpogKRXi5nE2NgVQ5mABFlgITfR6M1P3+Qe87BgxPVxzQDVNDXuAcVOjj7
wuZQ3BZfx0kpCCN4MxrAxtzWtfmJIqxF2DlYBZ5/BdFHU5URNOhA38XrV3gPuC68ycsgwwJdBTvO
z9sFMPM0s3+yiBVis/JMLMkYJEhvPHMaYTXXhbhq8BT8F2jnnv54EPIiGObIeHiCZpLdkTqtyC1Q
Pj8Ed0GnX1jhLYYWajdFkKzwBipcbo/EUfeRtF32A59F9/O/FPp1NjDyWq/hpGSAaduh5EemLjEA
ruCSaUE3OpVm6vfH7WvMmTOG0nDhD+SKjJh2mR16L16MCSWoNuhw60t0JzH3MRSHwkpfeQ3Oj14Q
ycKy30E4b8gK9QgB6iQyqlD/aay1plITEH+OPRIf7tUowR3yJ5ElmWb3bBHOZTq2nIKgotETlVFC
c0VE+BIpQetULsaRkTwR5IbVZ8aLN2kySyQFKB/TF9a2wzt39+gXrmMsjl2Cdke3D8PaL6f0RusQ
EGLMpWjsExcWSGxY0wJGTJdWDrN9zaSlpZnRSTG1e6woEarrVzRalnuxTrNEqkkc49fIyK7GH1Qk
0FWtfR/90ieIdlVc9G1gUepuJrwSdubeVPdqKlDdzWQaccNfe2r5VWrGRz/KBFx+9PiQ3Q7phHxJ
/xYzmZF9MOwrZwyvK6seyF+HOs13ig6ZMC4Myrb/bFoTV2KBp/OoUnGJtSYIIIpg80Fg4aU3/V+7
H1pYOQVAs3vGMmwNUdOBMCHNJv78hRCCLKAzGYvW3YLnoSlxQs2WMxcm68PelFXcX3F/+aaCT/AI
Xpo0JG9DZ7ygDbgVw158dtvKnxWmAaBmLdOaPOHqgBeCvn1OlfOxk/bbhn0mYZ+4QmwYKrbo/XvO
a6+R/OpcJ/FDMtoCUBKh48/VNilfU7Dv83tgzC1EBiaZVCxZUwNqgYXJCu1FO0qqrbphEhQRsW3C
fvLDuYwwep0b2SaKovOzziR6FeZJKSYT9tABnPXPLUI3Mq7hiV7VPUr6rZ113AvGPQDdBRKoYGGn
zR/FzTMulleraNdbNJ8aZ5KYlk4efqNMVMSK5BQzeZTAjLuI0KX6587GgfNNt5F1Sa5dvTTnEwpP
aCXOUj0vFie8iys37vks5M1JTMiRf/+HdqNOL5GHixKd3JVICjvFUjUqfGZGr2dBs6Xufd5z4Hfb
Bij/avVabJRLgg8xndui0udyviJAFgkj5YeWgYb4My54rjrpNIsAM3gubwPdNgUj1EufFBcBg2WQ
/WrphHeyWE5ID07CxpAmhKKs2TxOy7mZGvU4yfyFcnH5D1gOWRgptbItTARV/nu54MRbFV/N0GMS
bTTO3nL3eaeEQK93WrCIitEYjA9PJ41ZSt1GyUuV0+SZWKJsLotPRO6ZJPagsFxpfG4afgDVMqJ4
oywHf2krd+HP6LylMiqWQL9oe5IZ508HxP1m72cQvVRGZZ8pBbnM4UwXhcHAVuHh/r0p2zjQBnm4
pykqDNSFZs9yvF32P8XKyeJjsYsug4CCuy1I+UXYSv5cXQkS7wNtxdHO94Ye6GC8zg6d1TG7A5Xp
IYG30TF2nN0Rg3ggNBJg5VRuHamiZzO3HEUasziBfRdcBmYfKl+XZEulO1dX2C+BUuEkL0v0OVO8
dydUNhAffu7h25WI+GlSnNypRKTnWjqWLvMgcbhpFid2EAJkpMpQqTW6Gj18BptAnv2b3BLhvnM/
m22y498nHTPM/eesmJ2rNL7E0gDSmuCndubsx+pi0iCcbm/e/3wZY3qByLa5bTGacduIcPrivznz
ar2qcTHg1m7Rgi1nNDjT5AKqP+haHHohE0kYxRyfK4DGBKQgAfyex43TpsbN3xyFYb6W0bNl1OCr
pphuX/TR6il1yse61g0zfF/Z4tctmwAKXRhe1wgoUTBpnXDiB5t9HX3L+Scf2O4/9RNBr4Q7SiI/
K9pmNi48XGZgzmYPtceNWvPedUFt44XWkT1v2t7XGOdk3kTi9Ath4HHXzXpMH7XbkEVA/Cwm1ohJ
lI06MRDjBdWIfrEdgfOCYtH8d2v26UGET0x5TIfMAo59MrxLUJfSyEdrxt17382OQ+f6PgYNynzZ
aTff2SlFVKaeXs5PqrKy/ujHjFWNCAvRddT9l7I0wf6pLW/f2ttMoSq0YYykQE4haxcsBXVYmm4I
m5d5KElh1N716EqLcFiQPrQDMR7AyuZLTAHQgcGXADaMuVMUglZeAZz+gQJRB3516ngs3LVmDm9u
uNatujAZ1lX8BcqlpqWjBH2kSp6sXmFwK09Zd2ZrMyTPcZVdJOHwAWatLzwSRJ/0gGh5AroJ5u1h
iS0usoA+ik6Lk87jt8hhHuUaQBN37j4bzlL1D7zl1jUHp5fWe0s8sOROQ8jO4tXWgEvhlLgw4xmZ
gi3qrJkm2YwZFxid180iwX6l9LONQOHvgM3KjztsT4QldSuGb7yNB/VoYholqqWXE9ILm0s4zJ0u
lN7UeDg0krFhmPZ7/WOEilZCYlxUw4mkiqvYre709GRtifihpKVHzXVzLFucRAvUbO7FAra5JWNB
wjctsNKrtZPGIU/5yRNTKqdWDFRLvgzSo6zwxD0BjUt2Lio73ERqqj8fxfJ+Vj/CLiNkqGVABopp
WBu0dSBYmcqa62ITXWuPQw0E08ocvWAosM4Pmcl0ne1imbKPM7jAS+qg8mCQ7HN0MZdwJmf0dxxR
YmVYAYZs/LQMjlbsZl4YD0kywc5+abTQRH7jBrpe1YejaLl2TGrwZPZOiCY1IemPeYp47atk8TII
5r4yhBOAPQLdAIj6MF8ZjYwTBBa+1I3Sr+p2ROP9K6Hmr9aYhbm0/8hAa74yTiPFX6eDmWH/yXC7
LgOLz5pvduZV1ZHC6QW3kBaKoYek0MNlrxRj7mvx7PzzeMEzF3RDhPED+VqiBCksadyXnfT+B49y
9C6bii/qrBvd/jNYqmsHsZ1iwOC8vTOOX5uWRthdcLJUU7HIF0cTAx49zrcKHpK0HnMo+JHda5s2
+KQaXlsd0V5CWjR9gOqZaunXybH5dfnmBanXdf/FVFddWKcX+vIt37nsFHSllmQFiwo5kxJmHeFY
gqY+S1uaNY9H42jAu4VUoLDaZcJJVXswn6mvQ2DbOH1fl62M4cmrzt1Qd8EU5rhGiCYKI0U6BrLt
ia/WTSxEmDnv8C9po5ryQRHrYJPOSIlvYHBY1baqEBWNxUSGVm9vJEVTXvef+PBcGsqCa4YD8Wm8
J/p7FZy1fEXdaGCKWhr/h3IEPTdEgg8IRfPhSYE9upA59hfKoyi/3KSZmUaUuJ+lQVzTU1Y8dE6K
Vsbg3dOdQeL7CV3JXmimVnbYvjt6wAgyQyNF+3dGRVZuZYbWOAjNPlSJDay8U7Fijj1jUb+RLGVT
gnG3b3tYgYm8yfEl+D32awrEO8sH077HprXQrs1dAW+8mdttPtcXoMNJ8z5sHECBp2FbKQvs8Pbd
N1yjN9eju9tF8kUFAIdUVcKl5cKxUtZZIjQuZ1BAUk5SyqU0FeLMh2uBUWStFXY8iOtzTPExSjAb
nFDFjCrcApFIQJBWczatE2m0KGQnMPkBgzTnc3aW+MoYfEVeRE/QrJ/2eUIiuxaKHArbDoleP4dC
dyjOeSH8M8q7T1r4u3dAbctEA9yutAx7frcDLod1ujgWU5Wb5fd8K4I9cwwXhHH9+8Pg/EAMOb2R
F2Ofy7CCy0oVUsc7yBkvD1Au7+9E/93LXoGLX15MMUVtxKy/binTp7+8e+MQMA8f3tKo8DvtEk9c
SIOs0P1aZcnuJGV5f4o37xwkw19kJgzXI7O0tmYQkR3cpFr5DrPK5gNuzsW2MFY8LpWdWdGCq91d
QALqPPLx/ZNB7IRrrjFepYY7zgf717B0+PFN40Dvmyg8NrqS2kCUJczDT9r887glRJY4IM28Ggbz
cfqR7hKT77SOyNgEeIDgexYmOkrxTGGycu1RZdjhd4AngtRsijXKhXn2OSmD/+iHoLzCeZyu2Cq1
d3dhbaYc1MN3D+vXVA+WaVZm6UR3YIxp5Gul4gWEG+7MWrTtol3B6T5JTsPzceGFH6gTUQXL/pv8
TKfm4L9XNKbhAQtoQFcotTjNawKCMaC4iMYdg15vl8g7H8Ky/y+a1U8R9OqHYMTrvumq081gNNNR
qoIGfgki8ZHdeRkW2fTWq/HiBwFTgwrQ0MuGNoW0WbSLZZgbhgC8G/4d+iF3kS19x2CunIgMvRLA
Af2ZkFNRDYQ+BK7aWW5VCUvQQVZ5JDDOY/DgiFrwak0sVOTW5Z6PZpZLeHchAfJhPEExJRT8G3M5
P1sIBmkM90MLM1wSux8hw7TJ7lr1tc9rR7BDxNt6eEXFu08KdZXwJfPdXd2ZG8NDDhJccHFTr3z8
/Gy+rtRn3GpuGxX2JrR0chAnOiL2iCu9sNUCWO4wawnz4Eb8YrBs6qgVII0qwhVuX3BO/1FsJToa
LoVJS/qaaSEnbvnZHratkdiSd+FxfjN0ddc0N9RE0Z2JJ+jpGjIe5dNVC/ylfo55NobQIM/sc3Mk
7L9zSFGGJaoLW4YpIDP+0D+Ev/57BlKNfoOjuiulFKSp35J+0EIgArusnphZ0bQJefZKSs1WtFsz
XlL7bbvjBN7GBshhWGpqPIMz6U4+yN9FLtv3fvtuuHJ4FC2Nqg2DoJjA3dw8ijtGf8xZkGXz9dVy
/0derhZTd8gi2rjsNRiHURw8lScPw6a2VdKz8oz/8rM8z/LFE3RA1bY8xd4RFqWJYpEwQhkmU8H9
YyjZgNg6bxYvx6eUvVG3LZ/ZTQLVfAMu8Y6VhY6vLszDzdcgR4/To10+GyR6vjxN7cbW8FvgfjzD
SDh6CJLug8w012GbtATqZhf3p92pJZ+PfV3b37xwmRZXgZdN5Xsmbf/GJV1/gMG3Zm9++kRvvKSi
DDMQlu89BDJTkYJnvJZyIUjuheCqPKuVVCJ48ZmptAr/HUp9643cO+2C57vvH04d9JGCV8DNLe1a
9E8ghUo3nrulw3XUtPPUUuq05RBp6PZoSzW/nkMd+41m67gz+xdQGAjbFHIA0lxJFRrr3iCj40Ws
jcj7qiCg6l7TYIjTrA19wZRjohhQe9hIXQE/DQ8vWtT41rGYLNkwSK3vcF/CU7dpDdWXgIZCLqE/
be+4fYo+PHtBkIWL9G/P6L4IAgA/5pk+R/fmYckrpQDOU0yydYA82lDGWoAUKElvV4TRWsKeVFZF
OD/DE/MMaNAoCpSGUj2UFR9ISq37y9AYW+2fWumTX8ihsKxuTCFSn9sN6xj1Cq4XBghIkx5rvDQW
lYEU+/pVugA0W6RV10sGdr95BSBCKtWySPUN8wdurNRz6/JrcwIw9voRlz3HXjL4KrYruyZykFEB
F8EZnjWyIGDRSm6GzJ/kVu92Yqr4WFr4CgMAHpDmyezxq5WFOmm6noS7YK8XTE3DurFzO1ZlnQ99
hYxTqodZQdPabv2D1R5KY0C1Zrb4JewlI5/cvlmrRdx30Vywq7zOywyv9ex9+tkSLYc5Gq+6/MXd
u5lR0upYayaQnj2bPpnPaZyX7UQzgbm8t61Rq0+kftZCUJchd+wYBV3qFCF+EdJPpHkxSStV8qo8
B6/EZAvnKej2zSixlm5qbLJpnk+H/kTR016GcOBAztnDttE0DzGemQdMPpOqmCvHz1cu5DfNDFL5
ankvZRn2Unvo5/hyGVcgoBN6yPWDSzSc3ji9Amg86TK3Z9it3RQM2+AykVi/W+r/7Op4POTKGq3O
vP0F7YXHHczBsGPMJXYZb7CFtADOXFp6fk8un5y4N2WVzx9snerAbqDcLjzVpqJ7CnVCE+2BOyu0
FNTc6yPPDJ7wGdoVpX0HKAjdnJnIGM96s5o9mIuMyzKVK18CJ3uYATUEpbdU83UrhDHBl6M6geTM
DIM280TWaDw0geXS36KdUUTMD48FkCJlZOfEmvHl6ury5EvDrqm9QJg7HhXrJ/IXRwF66iKCKYr5
G2qTGXYPXEnOy8sd598CYVSRPLlDyXEy57fxP9zrAWdjFqm8uWRYiafE5cXNa9unr1eRAB50CkGh
/eK2gORKDrIZaUj6eixgM6puKIQCkTDGG++ooU+1IuCNakLoFsBavlpAB9ITFuuCHck6rS/NQBGf
YscdYYVAfPaX7V7UCJnaSwLUHMcegfL5eZr1Nfm0BhyuRnK2yFLTFbSoHDU1fCiirkkIU0uPw0Xb
paE0TPSOINcTJ69ZeyB3mxCingqbkulCrs7pU7gdCOpV3e4ayzF+qeDa6IBlddoa7btUsGikVlxU
mpJET9BiAdGMOz98wX6wTiFy5TwyGXJW7FwKI+qm3XIshHtgZr1LjaTF4BV30oQoP3vqBSBUx/TT
oh33ILMY+Labcy8DmADCk0DW2RWS3/cdkBi+3Mfh3a1/WGThSWkQqxyuKnlFBfTyRGkl7kSNF5Kn
03x3+YSza+Q7uX9K75lzs/qn+fMgH37nsfq7qaF5Y/vScssYErgM+XjLqpi77wN3y0wgzl8HMNYd
ib9zkr1BpqquRENm3xgdyTVbseLVVm9Jxz0OHpU3gK0VLZWw2/oaQP/ZT9Gimuz6+r0xAkXytlyt
icqkRjk2w4SkiJhg2ybyYecfgjH6DoNiN/R9j6+/QqFpQzOMNUOMJJQaUimfEscm6CE64cJpxj4a
DPC1E8DbhXcTemZWE1uCwVWf693O1/TEu3CxfaJwcPP1mefJtujVSYI0HoLjK3j+m6/3i4H0FTvI
R6Pm3RjxIZvRP1ARLeocqvJitsgq0nlYig6+iIYKx9blVg8MLhNkLGAFokKWndKpZJI/V2oAwx4j
7LlIaRS8zYMi7S8yVDr6CZZU239fMXcsSyzng9sFDCLgW807lVs8xh39HWiE9aymXCO1OAuOb0Db
oslcdXbONk2BnE7YqbPh8BnaEoy6Ec0t93OK0GDJT1zbh3D0sL2rCsf7/stOLpvTb30WeJURRPI7
yH/DLzrJz730pSNdWyTcw2GSfJj9PaH9+vJSbJnWsG51FMAh8n45Jfs4eLkqPTqZ5jFTdNN7Ufra
wPmcnl1OGnB8t0rlfEoH9WITN4uStafQ0cWmwk3tWkl0JdcTEC8qtUncabrUUtQjAYZs/2FsbyJU
AVTamsuUibQmwA6nRFSWBZBxp6Viws75LFJId19Ix7QMuVXSFeDmHzkdCX5a6NNtv/Psn3+Ubt1d
8XxFvr4EE2loCEKZ0EF2qSoqIfnQWWGRzPXVRQsVs12GU+zAUm4adt/Xl7347HmkiqCufpCwaYaE
Zf3JgYTLuqKjK14PUwqLtvLIeYblpiyby3zP7KlXsLyiVj6IJJVgjrg/sx3/DdeMqJl5U+tYMOE7
e6EIVZkG4fIsl28BKYiy2fCafaljVrETUYsj/tGcRNA35VF6qVTG8Wt3+1byVHNA+59BlAFrqiBC
QnpgTpexE+9/vbZ5VenRMsij0cgvDAqiT/PrRT06ADcvD34w6lf48v5w2ksdIz89/t0doiMEjNQT
2WWn6vIyxeD06IBUVfnkv3ZqltidPUsoigcqWzwO7xFJk/mgmL8Huxqth6vCtt9MqiF8QY5kWGJj
VG8soXRQPLg0a6QHSSJg6bGNNo54w8cUN0yq0d6ZB8y2xK6ULCBuxgd6jnuAQwJkHtSDuR14hD2+
I6S0nduc4mrbPYetOCUY3bHy46c+rvmcQIpnak9wBiRmPsYbGw2JDcernMOx4jS9k1NH9GIcxRd0
WietihOjZ0ai3TTuh4qDDeyt2TqzWWLJy6f1dfdf/8m1mh8eOavNUPPNq7ktadoMtQaq+47BaAt0
8L/547FGNWadIJDpZ+M60MJeslYiq0sKpR/n+zuM8ErDoqJao1geRqawlCuZpqwMXEsobScGnW5t
rbTrWrNKXizP0JNe67GQyc0n4qqJLzKoTBaMkeZjDMGNpDhSoP3S1X+STPwxDqSqRO/qr3/nxb49
lL+JhNI7lFn5lx9v8fJTUdUAth0E4OsKMlOqhXJq7W2L+LbFqlJRBgxQhp6Du1uog7P7KC1xZauZ
fRVXnEtQU1VBbuPKuMkDmO0GBgtqHE74OBNWehWwu8P+KMDl5qwCAR6Wp2BSEM4Ei+Huj+sS+Mve
czymHMDDcS+yFRpLhIHmk/z3majeBogiERRcTxfU5F3hxlXlWGoTkHfF9MY8INTcQs9aKW554A9S
0c45/P2CjBjPiJow+NL9/+weLpnXLpV60k1vKn/K98wpBU8nXb26yvGGVVZ9eqyE/l2lTPUahVmX
DkVVGuhEQLvU/vaodpdeZo1tOpHnQJrrUFSFf7PjRfK4CWPHPvt4qX03PnhyS0wdY48nrPqshkr6
ztxKHp6D84/sT1ORek0XE34krJwn4wY4ot+6q+SRgmPidIDOUFXyACBZeDJBWm4kQNollJuHsxcx
L9tYWhUPG7c/5sNJKMPKg3jCTVoJCpKvQF3ojB/lQbuNGJDCXGbJKEE9v1xa6LwbvADxo7hZxdWi
FiMu0usAIrQrsmSYen1gWJ/dIbhYIe8JuJvvsWvtEEuoyRzM9USD51yeknMzZDvfxTrZ+Jx3LXu9
MMFd7OMm3lOfSYUJleOUF8hOwVrEWv7SA9UU2k4XdUPqtZ0V5oQ794SQ/j0dLar5o3EoTsrOIMSU
Bw8e7XG9dpEVtX1bRgHv/iKTs4tQg247vkap1YC9PN0r0Fg7dPsXguG4kDQX3iNNaPPeODpT1JbZ
NfvoW6A8mKqEaZJAXqvRyqscwZeWRbzLsnCvdbOpSt+8cbnZJLh4L5jEZwvG8v4iV1bEk7wHGznx
0dAsqrd6wSFljIUu9pWUhtwxCjVYSZGuvdi4cI6JAKui7ZYrdP6cascKwLOPfO/4n+PR7CbwfLFM
FhHw9t/IKoSH2HT/j/Wlgj4Fg6bJ4KCZhT6waNU2KSPIgNKvBNzWV5166mBWEZhVh45yeTI9LLTo
F6kRg6HDl/p/yzZ324LaoEXT/F6IDd5yc+YMsD/FZn9L+xeWmS9NrQFwwYT2MtW7Pv6DI4tCaJrZ
nS49qrk0bwRuaAizk6/9G9jB//5ncrgipClG0PRyAdIT9FPeO9UNAUgXNiP482rCIRtSnTiNvKsK
UV/coh4ChQ78fuhEu/TiEUx2Xf2V9ivn1cqNbW+Tr3v2XJQqaPKrn3ftQ+Fqy2DLbhxXruapTh7t
cXz+upQV4Gef3EMKWX8G3lj0lMV4STUXbiKq+dkAYS/lKLwDv/PFn/hB5Wp0IF1xlvtFZE+kvU6H
tiIZCJWKRRNr/4OXFgr5uk4qKWiB0Lp4DTczV7Jr8CdWT4d5Cu5Jnt5ynQGKEewvYjokSp4UMgy6
CDeYMD4UG8gUJxJU5YthKBvRwVX6I22ykLXZW7cHUCDr2HoqXoeVuLWt6klk0VmLsNGCmNmy28wB
CJF6VwIluztBA7EzZbKHOWVTAr6WAWd2pqQ70QqN9J2ZKNMZ1rME2mQ2Pw+iHkeCqou0vHJTGEaE
OL/rUXTgS56voUJ3gLcspR8cTiJn+9pCHj6nnVl5TyqDshK/ecxZTc66Apfic7U7uOGsiq7cLMBk
2oQyVvscgjkNaMmmuxgokCoUnOT6r4hiZWT7DE2aaneVYQnsMKvcHWH2HFctPlrYwFFdD3B5Fye7
KiwHWWJsVXlr9l/GvDB0pSk0+BbHFI7NMw/bXJ8POO2l/gAMLXR5i7P5hByS8uepzWuOqCqEXv8e
BTcf4IM0ATT/aKooCYdBsZj36cco13UHs+V3vKZ9wrn8SkC3mSad/2SAvssURitwejgYy/eHLlY0
ajxn4zsQ/shlHMLa7tz5I1jhKGBKMYE/XXQfRIc/Cz/CD0XJdd9RO+bNceKD+ql1U95HvYvuPcZg
s5/z/mTQE34NyQDJI8b4qUelbVOQAM5bltRn7VD7Sje4Z7HvXU5wlypsCy05zqbX+N0R35p4QptW
p9Hv1kMu9oYDJfvg6htpWW5KVJvaajg2IxzWIVPUn6p4kfZbiZS05gF3p/JwX+W2tmBRCnjbye11
puzABVFrgHwQHvsI/p0Grkbs8mncInRMVf6pxm6hzZogitZbeaVgECxawgG4g7BKHDcA1CnMzr5M
7PVuIuYkWr5vDVF112me1Ownu//rlsf1OZz9psYmm8nGDYh+YWOfmJotTjHnckpSh4zlA7zcMXB3
HsPHzD9sAvIXNgKxzt6YimKINuSM0dl7+dam1Xhgnrd2IixVRKYnhaxetAVVw24z21plIZnoeJSo
7pFDD97vK75u45Sg/ArDbIL7DzaBQZ4lcZs0UU2eVEQIpoBLMsTmHrqxARJKHSliU0tet3gsRq8Z
ZVK/9XUQk+hZTRPKiKbyTjEKCx7WlXMNjFGNjkIK0m0yPjFfk8mGRS40mA1o0DKfmtTbjrpLuvkb
3fs80qLY0tABnCmjjB9U1I5J6ALkDtYGi0gpWhtErQ/z36nW7ZHl/XFvgxqTUnyNf2KdeM7zqWk9
91mDnahwqj0v7GQM0xrgepBasuoJI0Jyvu3nQEIyiN2mzjseKKVKY1IiPaqOZr/6UAmNX7Dhn7gK
sq7gp09nrcYUgW0IexnsDwOioYgZckPVs1eRFE6a0vlDSegHjb0CIC++nRfS0JOduyMB6P9IQSbc
2qy31Z549Tiz/7t1M/JI9QSpDBJViIhuyAvTcLH1gaKx0p72zMX5Bl0M67U6SelPaD3cyZrMU1uV
ZEdO2A7Op1AYRiz7fqMF/iO+xLBnQVfY2iq7MXTaX+67hImFEnJGSy31WEYjLQp3LVUVGsB1ac7X
MoKmOP7gU5A4vJanXpsm8A6Fy+W7yD5iWLDOhe6wiiXH9DquTCLiLErc02ganjWfTZ5alXwkXj3C
amsqF5vU+5qTEJskQVKLQdyFFTHGlnbdbhy4dwEJOFYY6Joq/DFAyMqqh2PrS/DfgGCmWuRrKhWa
+jmEVsKM1ZCt7W/1p8dzKvrCrR9cOwMBEkR7FugtvKLAvKDQMFryKIpQ8lCQncpCy90vQYbcL1yF
U/tWxm0VjXVlB1fbvLRzxqMtQmhSi/u5JfOcE+3fOdGbzdCKhdO43GB7hVN7ml9Qjtp79dksg8C8
ZpsyLaD8Rojd+udW4F1lq1nqAji6l/FxyOm3TGj0cvRadJcA/5GNn3DEzyKmFg6HXjUE8uHZbznl
odsf4NBzjyPMO0f/B6M+yKzdpZpYx6mSr73H1zzrTqomedf/ouie1rsFysCAV6cgt4auPrcSpuf7
dIRON989Vs3GmrJnENZIGoiM7/O+YpJlokWNoIoA0suzlgVgPOCkSnPKrs8k9gfBi/94HEmhz1XV
wGoNPYCufVL93xGKmJNg+kLtkqx6R412QmT18qgt5965vrMMdcPQWki7epQyGewILnHwGIgz0IiU
slB+d5+q1TggvleUWkaEH1QL2jWh67BnQVol6qSaisKUEvXAeijucvPSY77Yb5ZlN+Uk9joW/9hn
hpHGTAXeXJgH0i882k6ZIQXKKxBBpP62e5HN+YxgtSFAWravs0aBY8NZjZn5wLUTvMKCPZBjlztU
6y/tgYEjoR8XOVnxTZB5zcKGgzj1jPPBomXHWEc06rZDylQgGw9K9Xr1BG3Y7t7FQ/Q8pmrgyaIB
cHKvf/PwvovrnRrLG03gUoM4L/YGpukndtTxcwbxN0kLga+J2eUfexQPcfHu4NiPBhRfn44OLNmO
HIEZCVCnLKtpFlffYZ/t1njGoXKDvYCWziGle2Tpg+IKV0z4t+TkhLh8h9EfPCQcNdGOT3qfA0Eb
xrlkvOZlQNHwiKpuB0JaWmfsiGAg+I1rNczYX6yZtTdUSMtFzd2Uq29K2VIpayOIpzMAOdxi63yW
plN8/wsR4cxhplSPSxSnUS7JbZYZgnRN5tG3Royusp77d0x65trqyAFRU0B/eUcN2T576Yssqzt1
+dVzG2o1cHegGh1Ym/bmFYwiY8kWXZojFtJJq+pH/j0wB3fFaqTJfU9gKr5LvJVJh7cO1cFA8+mz
pAh2qyzjJMlD6RVB/KWZ3K4+zrc5wS3nz2TbVXsMSoofFkzK7M/J0n/+VM4rfXVrca4GaAvDuREd
NV+7m0fmn88jvgdUcbQnzSanH9yspqmTZPeyhnDzYhsc4ThIgzVIeacnztPxvfMjIUnmkP1+SC3/
vq2euHn+trmbRT4dcelrcdlLF8zu8PxWdCET7J+BUbTzZnVwsy6oCPzDdTJkroZJj+stMQvbn40E
Nzo1ttbq6YS+QqGZ3HZOm6odSg/DQBEdAicrpI7wTIIx/oFGQFb6dXnGlQFwInLN0LzguNxhIiFE
I6shNDusL0aVbHzWW386fbJ2DdDiTOPkfIgb+UlxM69XqRbrNLDrhEXkM9vMrAAQ+xPuUSzO+/Bv
xczQJMWFbjvIeNt9xmg4l4/Dc7k+8ORu/X05cuzuibWf7vfrslySgbZL/0/k1hie9VoE/MkiHkCe
JNixeKZkOMxKRLru86yF3tbCARQdlTs7I2ainvgw1Dr2AkKSIgdFhfVr1qQIQ4e1mXQYY6Biczqg
7QXG4zY53YiBXfzzgWDL+1MB2lrw1vRATVVanLUqqBZwhE7QpVYTX5bWbxMPOrmtbKtmac+3eeAb
PgTiKYSuUExn19/C35SPVrt3mp0TNP05abTUQhigJZidjfWGJLlHjezT9jZWd1aya1V2FA9axFS8
XxlrSAEfBsiw7d4rOs0HVBBX6zXSgYYxELAQo5d5xEN0u+gJSxwML4b0IjLnq6p6pnqajgWxURv9
SsWpqA/7+OS7UT4rDRKRiboB9J0b1xEeapak7FvabWyipisIhAqZacgUOpFtrAHEKPE62U5kEwJd
/0HSTja4bfC4Y6O5ksDERCIdXqYea2OuDaOVgRb3CxTu+vjwAlH6u93Q/jj2Amch0wFalbqM8OzB
aVqlApFLW28WtH5UH99QhomVV3Ex15TIDbfP6fihzqlcB4I4gSvC4OE8hNa2vXSwnA3hae40s8P9
mqMtEO4MX79fnJgBYeKM/kLGezf3vvYSuU7yApCQbs4+wDEPqwToXttFTk7StDHCbavxiH49bRuP
6P7U4+IZxcbwX3pAfBvdreZM9b88/UzNlzb1sTBOmOgyCRrZLtNfEo7/aElnYsKxFh/n3dFw0TpB
BRqOcVQ8sFYiCOmBPZ1+tADCl7CAgP+QExPWoMkVR5rxsXjTc2XSowSHJYWdGBpUBS37aZXFVLor
YxOgcJh5qmdLmucsad3SLa/k/p2UKcNBy/HeU5XsvQoIClANR5fnSLyQcEEOoaGS9xtzE7qOnyFn
QDeK5r5Qkvs+S9hhq3geZNaIuko5dLHQC840tdDntmScUEni/lwrJvQ/FcIzc1TuH3Bjl7BLbnLQ
+UThIqg95K9mp9zIUwS42oGeqmqNX3px6+2wt8hp1semz3Bglx/lWoK+StFi+l8XXdJqHxPRpT6y
2O9+MtqlYlIug8c9xBTcCFZuFWf6Ukrk3tCl5iQjfaZ0k+wqwV2XMUGM1z/l1eFLwWRzPJHe5Mvj
txvVXLGqg6AIENyBtX8a8gDLCnuC1XEMnH776wNdlkS7FvThkhXYA1DVlkzbzSKhpNJyEnVLOyXm
2PDNMLcCQGib62VYjYuf7UQNrOf389fCXakMQ8jjlP+yfIeM8+d78bJ4YuY5SFaAJaOObZPUTZwo
4HeMXp8mYka2dY2QcRveasIKZGF0xw+V9oAYJZB5jVodSaWUQKxT/rZjmYujgrncr9fplZbiVR1+
g1+0pNmemN5da9ZsXbY0aKq7S+1hxt0w+YEbFvWqoT5SdE4VAFNTSeImu0oA2yW8OgnflL2MwnX0
dm8CE5GM+h0YJijptpanJcdnd2xGB2CnHMFgv4V/cef0mGlwcqKQEDHONhgnTMlZlYoDknTvy9S1
sPbUsUekT0RiiNNc2tibCBiibMZmtO8TVedSz2odNvwxv4gwdedgNAw0+2x7SmCqCArPX5nPw6xG
jzzeD/SM8dF40sOCEGt8eajm8gllKUh1rmjAAH6NEQCR8wNwOxRf6xKsplTlL7x36heq6AXq1xIy
O9j/uHX/rZ2Zu+jtD1M6bCByIMzUFbwoP9VkrN1LDmYWKr2/BpO67g+nILXXbYKgUSy2cobZ3Yrq
DYseWXSVBteFywkzBeg6ajyAtFpdxxZuanAxV8gbPjDmNwLeCiBYdLS1lEj5S4IO+09rLH88UuYu
jzIA5Cv8XGTJap9xY4BXkKbiMCWW2mT65sjxasvO4VG9DOVFtQljDknslBvD/p2gaAyId45ICaIj
oNWBB4tetKLWuGdr6p6LQbZbxZA6kmceL/oIyetYAsIiLD3GRG5SBp9hGC3D/O4VoSlUBdvOoy9q
eXmky7RjJIf38WueJjsQJ5qmYkyty96z9jvTAVRROK2QGZDUQbIJa8Inosx5NgnIKMP9Ent1/Uae
zKfiSm2ODlArmL7LFtfljH6/pQade3Lv7X7WCFjUgP2+Xon29AzKqWIuDwxCmK2U8NDz9vmCycUu
mfx/Pabr/OVEeEtDbxWnZTP53RP3cZzvf28rzmzQqZg3dGbAQiJwSqTUGBAW0zHabPz1y2FkHhm+
Yhpd28soDrrhS7LEVnKhhQeTbu688cIzKWNLqybxfhcaLLlbd8jpEDbyj1fshGnZzl66QL9loaSB
69IUnpq5rM5H5/4QyOfK4LJu441kVuuzyIr3Js3OGEallDtLv4oBGx0LB1vSfFOc9jXgIrecobMr
iS5uxnjMhGdZ0HWFfx8aRrD1+R6s8E+VhYAKR6j9oNp/ZzlM6JMumzklFB7mzh1FH8CEay9kndhu
iWg//stfvSJVk2m4LHBQ2znK0LFv8DnaWUZkkFybR6TC95siRGqQzVFw4frC4BymfyyBYRcEzJ/p
EpjN7XkwIkkoJyxo0hKLGoR/OjsT/WRJyNASS4ct0Hf5xuvhy9uFKYi/A2yxHPstSR0c13nmKuly
nRa/0hS/h81HwjiXWOQnKSXYWn7AZxHaXIy+D1GfDxkgEpMigDg4l5NLFzlQ4cHUJLHTGgKn9Vrh
aU+scRs6tLo2gn2/OV8OgxQR1aA8YiZJhLznGN09DMAtmr+reY0mShEusRHnhqs1W4zRFwPAs3Ag
55I/xuCBeq1a5/pxGeJYGlEgH84axp8ZLRl4m62TiEnaJI0SaDPziopi7Yn8VmfHdKE8Qy5502nb
4JywjA7ZZhfgI0jhtJZU14pOJn6TihzRRxVf5t1x3yn+RFNSL+3pvi82CktGcYx0U/zu6yPTAOZZ
GNI3nNsYfnr2SdHm+ubI9zk8GBhzOMoGmMFO9znIrrX/p28KTlHfDXry6TrK0AQRq/v99NYP7OV7
cUd8grCiqCchguPNwtWnYouY2+ddmTJtJTjEdBMn9IbPnigHc5lb6Ht5hOUh2rOwxN00Ul6wWfMI
SnSWxhOyr3CTRKbmR1u+Ji7y7vWjMmmBZPbt/EtDmkwMyZnFMsuqu5E0icIEbEHChccMh9MvG63g
fcSbB6X7Nc5noe3v17wtvCIssLP4k5jSgMB0zeB88cM5YVEHQdyUjLPTPXg6UsptnjDPn9CqB9lp
562gLstbG5jsOq/+zQ2+UX/X+42wGvJIsngzMnccTRNCK9J6FNVNHdNvnpQmfx3Jo2Rb9N8z7eYV
4535wfpd2Ar8vcK8HhTY99T+YBzsMZrydJsHmYGjvuhBUnsmQq2Vyc9C91vonSuDsxFzHVhZM3ZU
YK+n2rkHfisg6QFXRtmpfPzxspcRZP0kcM8CIlaEv9bXkn6IrsnjdQbfyfBcSPp8USUwXoQMm7kT
jsRfdhlBIa3E5YM6dcynUYy6+bdyKw2OLOS+ecKm+LmR/2FhTtedxSg6T/zmUb2jLBtPVXexHT3C
lSW+j72Ec26xoKZ4r4227kpgNGloMAuOw09+3NgBFsf1OXASgOH+m0DfqPgTnuWTWTKJ3hrlZXoW
myQQbqOv0ywHxuS2vbTQOO9t3ms4WyRE7UwSCDmrqEPYKy50KEKIfERfCJ7Dkwr5KIZLWwDKyvlq
TSaS47Otuvfdb3HxEnugPt7W5I8TGjWtkoGjz45biuJwFDq9eR5tBDzjNPIWUQdrq6j6GxIuGJOn
W4zyOL+9jz0lRqDBf/OC64yNg5EaauSbdRtvpUkndsaMbwrKSCq3hgpt4qZ53xoWDirljk7C3Sk8
3kGots3Z5CVZnww804T7PCc23TkZNoGR4QgIFwlf0GyoAUMHORjPuC5Wsx+IvjRHlE01aP1xpQyG
oKqPLhSyEEb2y2xh/nZzpZAA+6RftbO7t13DU7AtAB0S+1LMALeUARwvVQPU82AhtkBquTiatgdF
RH/HBRDcn9wsjwUup/dByDIJCKo8BWJIvVwaO4pBf7wcxm2aZok4V0LOiW2SynQcISZuFdvB2lhV
hTUNvUF3gs0sJjZmCrGjV5S3Uf1gnfvBvLM9zpkyTxew2SyNVbgGXfpG0PiayRNMjcTMUf+LfwIB
nvZTckCMTk5ZcISwGaYCzuyWfgX+GAwkq9wP3r3gqnW+3hF0AKoVGIJxX9PY01Po8wbgLVr8eGxF
rTSlBR9ngf+B7hgyfNH7UoBsxjebzLUzYaTpTMFLgOr3QN1l1FMF/tNJ/idU5nPQKGlLFpqqmHUJ
saU3eSH7eriGL5FK43BovhMw3I9P6QTaz5sRFGfrSXUaYXzInYuEyJN3jJDbupLL4HyrZCAssx8Y
3JEyi3iNJ2FuC8hkKY1e9Yprf07ho+S4VAImQz0YqVGl/k0IVKkpH69fqDFEfX0/VH+9XJqnbdW4
MKvhgQy0YGadKXmX7+R7ieqLudrFui73GJFmfYRVjwL/U8xyQN23g21NmE/b149RkwjJ/oG/1ggo
4a0fhwQqrRpbTdVP7F8PCCeQMAsVAx705n7UeFwUgLPsycpcQWYp7ppunFbltZC5xWzNYEg50zEr
uxltNHFdfqcH4OaBk6jc8w55JQjA8+hdILOYkOhU7pmpBzqufwUZyKF4oifz/hgXuIdcrgVrwvC/
6fvgCz3Jhb2lOTq9OO29uBq6Jx73UvsgO+PCRgZEh79j+Wfe5q/FYuHQGGSCoh45GUtzp8yWClSI
tR/5qigXNiksiewATy3zEcgkXOpp5z+1bAcz7XSvYbflGQZlsnYGPydvLcb643S3vJK6x2QR7Mmn
VK03TTy8e/WZzE2Wpjh4iUB5VrhqvPJpjv7ZTfXYpTcuAuOhKj4XNnf6dGlwl/5RBdP+gh42vX5e
2z/lg7JvHJ4xdrA3tcKmU+VOL/JULIOxt3uotXlN++7QLtQGdo3ldeHfcIq0r1z/93UpVO5PV6bE
HSx+a5VwxaeCaweR1EmJeilx8MO+3XEZEdKVEnvz2v3NHtiLjpkjSHL08s2DcDCRlM8tufYH2ht3
cYDrppw0+6bApokFNvcjQNgef6gp6OKy1+iQzdDJ+L3wEvcyWk3N9Rc1zUoRVLDdpa2tSTv4DZUY
ZZdXJFJX1j7+MQtythoAWnmLt6+MYjamttN7LbGyE1qLRhC7Y126n7fTUB1YOwrPa6UNx39GQGBe
1vbnLQmYd+IXOiDq7ejK6LcuqmvMCLo7JaUCcODDznpSeSouG7HZZFiJjDdAQE6WTyEWwRyI/bdU
v6s/tyM5dY6tK23OdM0PWcmPugO+f+XEhsZIuQCgyjfIHTK/cMkofWdql/WruTkm0f5A6P/owWTf
ENrge0T+gSQgqcW53Oay5fO94xSprFQ1z01y56+0RHi1Z3bM+XkT0xZb/BEILR70kRtegun0DbKf
tU6kSrSQ2j8J82RuK6brgVLVim5qYFoq4ocLgtkmC0Upn7eM/w56xmgin4EDO9QUE/+THiJmSsOt
pvicdO8he5KzHg2OMqsIOCe6bjgtZRumnubXOcC5voKlyTY+NFzdUd4BgR/0zdPUD57EObYpO+wj
tD5JRtnp2Vll6TmrycbacNtJMRgTppWrkDbQmcPS9JAMdGwbM5PAgc7rz2TQNztX0iY8oQNFG+ho
XHgkuvf+w9MHgaZOxZ8QWl0KoGoDgGyroETKA9oVtf17khNmW9RIko+CLoq0f+XuzRl+EBhQyU4m
qMtIKXNPVgGgNNyvk1hXNouTndJ23kq9FClDterC5oJjHncRbYxBT25muCWBF7s9Hbt/rLtzQE/I
xYLsfZKf2mFS8Wnh9DkYAYHTzMuRbPZAJvqigS39Q5ItLnvbrGYNRvHqr+CQPSbSf0UCNdx+e8RY
QMclSNEu6BBjkBCV7/4dbsOuXNxxverZcsx3+JULMOaJpD9adxg6zDXbn0F8IAAa0lF5CYoXKn4l
zw2jZrTg3LMYf85as1iY2NSIDVAmv1ABiXOQ+BhIN8ACHI0qqGyCO/NdcPFFKZW/m4CvrIynjPOD
E4F/yI+Zg1EuzlaDBN926c3Wzzfqib8VzZ4hgkRucPA+7rHLS0hAIxWuFlvm5MqNSk6zW61GkSv7
pi5UFlB8otRjvrZEgOlcIxAI6+8KKtGMpkrXUGrABufDeiaSGzNLXSFBGsoyUdYBZ3Ai0o7NAjcM
pptrIA+8UYdZtcqhLzP+bekC6MFkJRppZWZUrwZgOfLegiOc3QPhvixPUn/x7ShFeDysKDdPuXuv
mwg57wPxI2HdpfI3FMZy3/2k/nR3ei0RwFGOlyqf6AIjsP9Pi2mf5QOsWTNsdCRSKFgfk81a3c+o
eiRCazsRpRMr9uG807adw/Vf4IQ8MrsAYns3KJgHsW0b8dv20r8uc8ekAcqjMXGdoC/cKTKqqApe
DubZgkWmMC64HyyT/ogyGdRG9UURvKBlvO71WsKIcmGXW4FDsBeqA/8bF/Ev+N4UT+a4aFG3Ch9J
hFNgCooiLiOQqnl2YLlVEt2YNDd8R2g0ZjqmITfmKSug8bvi4S7L09Mf4pibACqZD9dQX9towoQu
AVd1KAIQD9xn/qIKq72g7s4jGTffh8C6/wkrjQR/yINxfpMsb6xUkYEE1fa17FncKXnxHb/KOlez
pdLNtMnDjdXxrg1ruTooxeTFT+w8p6AHbuHZdP9yrcE6nt2MpBEeHMmvLABmjBsJHZggDLTXyd9v
dv371JieQg+qntxDbuBlOVWMKCXBfWTbCSfGdxd+L7A2YbMdsXQr8EiLb0nH5WeK4EN+ajROZ+id
Y5qCxrczCOCr1lUDAE5kGjktWROfwcOksF4EXIHm9mQgW6TuGrwsEnMBUEoWU0GCaBLxvEiP2xLn
KBXF0ZsFxCZYyAXwb4TFeU828fOmBYTBHKMLP3781lcUSgisiE2BMVMYpx1QlfLjzg9gd/7yZGFQ
he3+dAyJHQWhNaYgonFJvncoUNINJND+pLemuLJrjUcRhpvCr4UWGzQk2OKZF73AtX/rmYQPnRPX
lx0ybTMVAgPI0U1PcE+H61qod8eW7upbQdebbC38yUJz3jzGhAodIOtw+bPPAuWvmMA1aVOglf4m
9Uy1QbOPqH/LBomXk4gOr3cis89yHO/25YS+ZUNlP4+qnOTjhPqUV7R5YFYEZKb02x8t4LVwhfx8
KLDYNgjVcF/EL/qsg6nKKQmUsxv5FwHNCQx7lftbWJWabgHCS9mXEIG2DX43aTZhavCS13keBLC2
h7NDdsXxSUd1zXfbWbrm7MW7cOcK6RNnQNdAZZmV5RSazQK8HwWmN4cpBKAwETCLs6COoKfYjIsQ
qO56qR6JjV8hhYDNSrUxBwRq54+eIShFEIsTMpHh/C+MQK7eokuUW7JInXqB0euZsD0xAvSeUnVI
Tcg/dibxoWf449+Be5TePPttXJYhS7Og4Mboehc1HIqsFntdBl7mRsp/eFeZa+wcWGhIj6QsFqYD
Oke5OS9p2KRowpV7gvEflee/oAlZp3j92LaesebUqUT5r5cBPIO9dYzByJ6ZQmDwrGwMHrt69u2J
kYbNnJ579rDX7BoiEG+NQMyDgcouIJjCUkQJ+8zgR7MkZ3RbMJrtF4jxAo/5d+0ZWrDF2NqnEvM9
FyKSJ26n9JV3vfkNTZBdysAKq7/05TBV+U+s25K8AWtZ5LfoVEcTWAN2dAhh4pAQkUAqUBMD/8v6
19S1DPlMh9RY7yjBxfe6lyYUThCB/UExbvPQxdZCpz2byukwk6tlJTcMQlJmTfwbzyR621psFrDM
iPVQhkpI/y2QQr9H6yCJPHB8B6RZx5pmGeJVs7VZkrVyltsKbJXKytY3q3xV9upxvwBrfL3oEDnl
ECIikm5nLE9NzC1oKiowBuUWImKBG2Q45rkUvmGgc9Nt3CT49f55UmyH7YjK50Wxk7FRcWZip0Sa
Mtcyzt12aW0KpE5DY8Nf/xokhhnpK5BV43aOWnNbU/t+G/p9xIuoKAh5eOmnpACtaoVrAzQOPstd
Ebmy1hkWMwRyfN4UvawMGizfmwtHZDXtPZBydOsogxHuZugcSe8Xmikdr8Y+kDBtL0HKxIe1NvfB
LCy+rcPdk7vgXFWkJ0AF4B4NYf9Ze7UvBjXGKeMu2htgy4MYT/d7mNdcXcos7353ByaWQ+Ip7zG6
VW1dOJYV7tBQ5j+295UT9+Hz3jXZA+V3RxWmU88mhrCO6cVlH5z8tYoZV0rJEQH6fgxC7xs2BQHo
9RJziM/sQNdZHP8LgnPlfLou2ncHiCEKV5MAtQ76ckDfObarPokXgdffvPDJteGWsz6ijY72cuGV
G9MdvANvK1CZ+kxPs67nPPTjm6L0zl1JSGyL14lNP95D80AxYOYVUqJdW3CPArOgJluMZCdmj8gX
6v0wGSxmBoDMfmOxLDBA4Kn/TC1xLJKyR0m7QUW/12bdTmhiWlRVxScGqmSrufVSq9xHBOvgiBhX
B/q0oDlkW4em5jnrG2oZtsw33iOhtx/xZAjjRinur3IN+KoWYV9s+QHLerAKWjtyVCB89d2/NN7m
93zwz6Fp/h8SRyZlON8YuhBGnvdba45IZZQM5JRhhzqUC2lgsiw922JMpH/id26WH+4B3ppPpfwA
5I+UoDpKDy3pR8WQmi2Gf8/8d0soGy0YcW+1KZ36McSNCWowDdJ/CHbz0mYlfvlYSxqpCj6oSve8
DYMQ50oNMYj4W37GBjHbpBuPs035WU41+O4wJCz7XeZCsEpaBRfkFQ3i9ZsrT5y1P5WWotM+y6kZ
xobMiH+Xg909/xH3YIunmjsqb2k5/i2rBrf6uVPKjS8PZrASs6nJ0lztB2+1Ivcw+BR3WM5jngTs
Kxh1P93YA2ax+5OMx73S5gtTrYT8zAVBr6TF94c0vXHjKhMXaZmGsrtUGV64mePA3/2J2zLzW98p
TR5+9AQovowEJcZON11SgHn6jYKe7FwKwAr9oBtLb0vU6lLtKpsuzGMZ6Lu9BYCbWT1h+ZjYnpSd
7VoGFghrez1ylfakDXqYMBfk9HL1c1NJlHcy2//TL55iyxVYKhqC8gfv4msuSERM0ygsI5hwFHjy
u0pVL6ofaKB3G/93vkNtA7HpsIAGs+rrWoYq6dWFm8PajUNjfoECaVXUPNoAae06XHkBWldmQsvr
R2EDkIJXuNe3S7WnGhBgW0vziAegnWqU8Off0cPuCHXrpTFVupYbQ2lbsAi083hkEun3rIMs6lwa
UM9mnDJVNpSTQzj3qfvctHU0z4pRSLTiLLukZyQ16o2h/OCQ2T2Zy+r+3ZDuh2uM0FYvCjEJnTL0
ORKIRRH9G5GSw8oJQlp7bSMXC8EdbK0eF8Dlhf5ry9+rDntyc/XPhc+5jylHbcUZt2ajPDzT0VgH
I/WbOI/a5lvdLeQK7RghJCqdfhUMYXmIIR1YY2VzHHT+ZwAjKQAzkE11/99xO6Ehh6Txs6DGyKEM
EMdd9sS1DxMl4z/71nL7XZuPVnUCu/fAUvJSs+7E1HphiIZGKDeYWXmDT2M7vwVlSPF6ZXuy96zg
1sguNjcMViLSQKkNNdBUlBTq07CgD5gPoLbaNhZzyIsAo74Gr9xPs5C1BfU1P0sBRKk66wFPXdFL
bJ2pfzmSWIAfEXTEw2YsHI7Jkw1eJZmWh4SWAIMjvAGX4vvrBn0e81Da2M/K+8Ox3AjYKCIS+rA9
xoDgjMgBZo33HX9lH0i3DfnhK1UClPDzrBiaiI7pa/33kMXOQjDSFCLt9vBWDn3G3Q/HXJhSezz8
9yp33GAjMi2l9La9fCVofpHf6jnv4y4/3Hbxxz7+C4Bv6GRcwo+M+Z+vyQzGiYaYsWYKAIp26Tto
uCgw09oKIHsmi2NK2kItp6I1oYo0rJu7/XP0v85hDXfnpFe+pVIaRedDdV+fnRLT+wZOwdPO2SeP
9LHTKAXx0VTQxUrXBki1fTLz0A2NWuIflMGvIV13xTeomGfBq51zfMLyf1fqDqnQVk+aAACneXli
Fo7gtAOVA+KD4rXcOaNCTDAH1vVcLlbsWen2ciWeAMCJYwvtlJWIj9NkzKgKriLcOQrSdz6HF4U8
9qYeDO4vOcUvPL3hucqhI5tG7cyyIE2+YMuydzL7GZzlMy+596q7mQW3h+8VTfWU1FXRahyuAa41
UoHajX5aTK2aRt1KhPjOhEUIxrdXe7YS7HRao6Q9kZ1o1/XfZLBdYu9Y3ratgt7A0MxLFc9TV5XG
E2ZeieABco/QQv5VvNt6YCEjMZoGYCtmPvLDqC9GN38lSGm8JWeJIPA6+PmglxL79h99g6rrHu0y
rfQeBAT44jvnLfUlvingreMKNV3OccshfkK5Rpxks8TB+R7YbM4DY6oAcQ7W5Q8QzX5KczQCbkmF
107Ay7zwyWS3u1Bo13zP+DzUxgSiI1uOln3NXl/WlP8feRQ8uweRaoYllv431yvsMAb/yZhMOBk8
pbjWYAn6jGfAtSUDkTKDWDEjp7fOK+vkhziKeUmlBHDRy2tqQz1XBxqnD2olNmt6z+5jVLh5cKvE
++whJOA0jgd0xiTj2G+jCXl4KAhSGLiEc4xjHSnpJOKrYYduPIyISU6Dk39mH4h2q1O9bFYuSpEm
W8GZ4XJC4ZzoWuoM899Ew90F9UOoaRv4OCKRDKicPX10bhqceX+BeNxg+gDbkpHrZAYFJwFJ+TmL
ZBWuH7CIHo1upl+KA/BZ1SUXl4zY7cq4R2Vj0JVG/ANG8K6z/xJb/5T3XeNHMrm/BwUVisXtcM7z
2MiZspFvAQhoMNFHR+cqNgBeATZTnBIH5vP696CcBnH2pjCjSOoKnY1S7+6znKaKmtuWt+2iWvR6
1kp8LbRDv/JsfgUrf/TXwv7O9+L4qjfVM1m4El5Oxc5DsT8SteJcM+FcpaOntudQpmTNGhVqshzU
WtM0iGgOQ68YmckMMbgd2lgwJ5JksIFj30fts7/PjOSjJl19/ATkEDXj/NQ/HVbhcd9wh/r+4GEc
nssfKaOLVol77cts4asYq1ok0gQjTyu2UgD09fGkqzcIkoBFibLPbUn1CoAqJhTjVPBNf9c7kmqi
+wIozmOyappSEfBiu844gRhNlmiqIgY8h+jcY74t+j1S6wXGxZObd3s2UXauAaqMt3s6kmnQykso
GfKwJ0PttsJV0o1MorA5Q65EOsUmSSjsDHZZlYg5sNWyo77hC87nBpPKDJ9mat4GtSYfooWwgD9Q
40XIZneIcVeGCuW7OWK2PbQKtG+96s4LPmpe/QIenDsowlM4+Rh8hOr3GZfwZMEyssVoaSdUq9pl
DCvZE2CYSjmM+V+OUxjWyJ/49vHPkatVz8CD8zd8ZsQo1eKLud1GMWsZRUYdnedsCD+Ummu/doKs
+/1n7oTGhKdhA9tYaop4LYUsZDFwTeb9KMIvZ5e6ZtCTPEqGSrFb9xVcMKeH95FM6Fl9ELqCOtR3
Se+VKg6KOkofkceIRUNca2kkfIi5ato2LbBef83zygGfCWSwe9IAqszllRROqBOlb32iNaram/6j
ba/c1InIUBJb1sZgDnEYt7ztKYfuUm7OpYffjRGu4VxjGNSaDfCIvaNa0HusF3h6P/FJiMevbzIQ
9hgcsDBFqbfd37kpTTpi9AB84fVkYNxeTAV3CHCnws8LkULuzcMMSUQNxQvhyEUjLwZ5GOjdXvPM
UyKynXTlAm0nUH0opz0c+/o3xwnG8GeJ64YBDk8F3/rfexNB4/Jp2JRuxGDOsaQdF6uCbOHiW4Qn
pIJPDNGFUJMJyYukWLl1hbN4BGfDt6r70ogjbjXmtTeGLK9VlU+gw1sIGXhfeB0nPfioRq93+I+C
zuJOwnnYjCZwMQqhPSPgrQvOgfOrh9+UejUsx9h9iAMk3Qwq7tyP7ZEd/pJoEFa7dP/kKFK+szEO
8IWPy7VnC58RWKpu6L7CE0+wTl53+8oQ17uRxAdAuW5ccwyMkLYOLumIkanhoJirodcIb0yT8Oaf
X9YrfET/qqy3eU1MR4hs9MsQi8Zs8/Lkp9wCP1XAn0xkuug3wRRctGIrWoUjYXMzs/21P5isWp4S
tOVntwyan5LRJemN3N1i9wH4Lz57yRgXBA1VvHGzL4SjGoSEC95JfP0bt7wHFgWvHY+BfdbKUKYt
z/MK77ulQOwSNXEI9hMSb4rDSf3JWKHWAcJvjRaLplrY7AgD+/4Kw9yJ8lCM1tu46g6S+RRYiuFH
CSNJp+u58ZhdiF4r04CG1ltjuCzNgczhH5yK1PbZluK2/svGvmREy5Ip+fMqPNMVitOm3P0xgahX
t2maVBBAWYu3+lcmtbT8RozkT1ePcf9uVwy0r5XpBpILZyoXbmDrRB00b5kDNgYu/KFBzlRqtC8G
NgHOvq0DJCTWUVVy3XqRvbB9MKH4szVR6hsFmCqR27xGSuNfAr/MnNdUZh676pBfz5hfsMqHRrBa
vHbDfQdkINC15U2xKMR1a9Nkcv+MZciGen1M44LKrsQbCOGxaCDnySOX4QRCOhKyl7HPsBAsw80o
kRm/VDrwSbqD4OvQFI4fi0W1+tXJfvk4WGOwz/ytojuEgoPzCTqP0iUWVT1c//PjvJaUhxuGulQ/
4UqyO9t40BE0rrgD8ViUb0DFNuWiimTwUsnm5oWUt57mvg3mVeLUhuotQ6bSH/Dqty3/1JlCphtj
vfvp1gvJfPn2X7oOISIJSt6nO7a4Ryc0jdBIxds48UrhVbCXzMWQpyWkIsCgFVG9lP+WulGqgf/d
S2/kUoZUec1UVCZK8FXF6jR3OQDfLnqtSFholU7ntkhLHp7IAvGqA2u2Csh3LAJ4Yjsik3m0RkRA
1tAuRaczegS9gIC2Koqsy0zVLeC5zoVysSeBFXKsq3NaZfa+3cgFrkiaUXpKnMdzIbBly1cbYeXM
OFqB00T+M1qSA2kl1kY/85AZ6pjFKuP2auRC0YGpRhTvPhtE7IlAPONQVQbnUHBrEaw2+8mE0yaM
qKbePCJp8UvqlZuONyxlqqLa1nZ7f3TXFMlHnBF8vg+N5sGzU2wbbgXIUM9VluoEQ3KJNapJHV9l
b59xnfJbhfpZV4BheOPSqHuAq0ryGf5JYNBQlJFyFtgTTUArytNi86GzNZRk5as8IOi1VDJIM1Mk
DCcOaBXgpygVnYyfRra8rS3rWobioMd1U9LcovFbNEbEcG9GG57YBvbtiHGAg2VyJtnVufh7Nrt4
Uy0fIzswFPf8ybMO3icm0lYtGJyQWZTH/cEujkeTK3jscwE1lbcWo7kmJlDKkZ+M4XvUpChKgkGa
AiJBVa4AQhux82lWCwnI0TGyqt/LapVip9RTJJVbE4HxPUCSrEqDCbmYrQdfEZleSgOHZCT2gc5S
eUobE1uq7poxsKJbAhsiCwfSOj+Rj0NbdtGsRoEswqLWBk9fwH5yWv9LAi7kRvY5h+iRNTb68zH7
rK6wfzbMRgNYa6UfkoInV7uiT6UHKERgnPHqa4/+yoP+pQUXMpIJTJhf+iyI5EFMFp/5ACW+5zc9
KJf5n4UeRPu1+8uBhL2kaEHq2mRkCNxHRhoLjtBje8Rm+SOiAu/ZVWakeTFYX5OJQLqQAa8o9gZk
EYpAfS5E7UEmcv+DKB2jnThn8ncqxkUbSqMthq9zqYl/aVCE6lMrP//KTl/boiQ1x6TugotsC/LO
5eQK48uclANYv+J+Ox07el9RxxXQXVj5X7uoeMsXtcKIDPXAGanXoeYPR0a7cMJiCsHU1B1y30qB
YEffZepuszf/av3iVfKDrahlbxIcv/IdL5Nm3WuR5k6bVrSFcrGpjnLuJYyZJdLN13eJWGaYTf3r
a9zybLWRzMSvcGsLUjPmdBPwJchQwHaSbuV4oeaEjx9CFthr+RXLtqVJ46CEoomSYpdTp3GvfEB+
gTHNLIrGK6ijEMaG4A33hTOW/c9tphDw8tCtwEc9VEwREB05gJPfDCQzBcpcLQQ86jVX9FnTjVeo
zbvzkj+N6wUiKKE4q0xLwAnGJcmstkqmd4aLV6wyrXMYKPs9j6NJWGHHY0Zjy6e2iHJNLWayQceP
wZkTImrIhL/c7klDBqs+zxVEKOk0A2OQNP6oUmzz5P9itfRddxn+PjaEjJ1Ak7EoX7LvoHzgdZtQ
VwCLEikgfZnS3jmD94H25WlzgMaImb/080ah442VWs2ZW32hCXkubnIVHc5IHKp3b/YahaDsifcV
cuLw+RsajP4bhRo0u78OaFnlA+mOu6n18RdiBS1MyGqS0eOa44fLr7vLRnLT0EBNimx2Y/Ow0JmD
M18PuTYSZmuE8M32mtCjeROEQoT9XxU/BH4eT/okyOcT2inHpn6HNeNmankBVuuDqbAccOoi9MTt
2UaAoHYfYpQKQIKEDfX+J/FwK6THP51X21jfJ/vr7x0JOX+0TNX+lr75AEwCS1uMSKiSdPNMIFDS
EFrsNDhZjB10DXrH/WLJDDaeerunTXBEy4LxeZUUdA8DJb2F57imVa3O+EJY8hc6xgEd95pty0Cf
x37uG5GoBtOgk1QB9dYp4nsiWkJ3AIdsCjNR8VCMFknBHzqxwdQcA3TRzQdofiXeCym3zkRQX+Ya
Epr/TGvJ61snTEBFhqZ09wRqpAyiG88zktBa9LyrPf4toqMAfnJUtPO44r8xHdy4VQB3L2/86dhw
qi6FhD992E0BaETVLwwnL8MGd8/MB0TfjAnzPJDQBsV8wshZr/PR4dpViOM0aH2wDL/jnslHujft
N6Rv4n/lxT7NtbHAoCMxZ1jOhTKGMRa9YE3YG6DWocznZZ3OzcQfpafu4koBx48VUpwQQ8G3RHhF
TOqPdVp1ltocKeBbRNeWQAtt5vNimfG/76UHXHmPhL3EM5mP1WAV8jfr4ok56AjHabrHbcRK/iXt
jUYDZh4eYAxP7kPBFaAzF4tS2LZzXV0EZCxgGpTsuUH1KXT0+2bADXlbp2306TfJMWfIbbI8fuCz
qgYFt8mF1eJzDn+izy25sGRjHdmE1sgh2ns9nyanJSeRM17ueYPIzRNElvFsy95S6x4LjcAuSDHs
x8KjPzP9hX0zjF4LxuNa08sLv41fkbO7OOZYVBGyeSnIjQXiNms62HEfOicLeyNAIX86f1/jS66G
HVnRi/PfQcUdfRWNurX5ftIR3B8xUYF88n2aX9SbswVVSmPMq2pci1t61Fs1t4LY7TgH59HvNzcr
073OrZvnmTHZacpEE+pGs326sBeLqV6SG5bAe8svLwPcnlEMZx6nu9EqmtOdiDbb9TZJnNS9p7cn
JeHPgcUIahHm3jP5N6EleKxV1Hife3LcNKflJ0tKLOlxqUWa5fgSFnPAFLtVvRz6Q7NIXwRt7t8B
atn7k2cgZOxmbPBuxdBJniUnQUOA5+3YR7jpebkin0v5eFe4G2T/mJ5s2TtH/mnVphE2oO0qS29/
BmJVNxjHIB8qiKyiiQJOtDj8YtrY75grBI/1QAUiLhw7Qtj4SHw5nDhmntLLX3IIMeHnDgE3+l9B
fV8+pqxp2ipXx9pXMHqklMzNZHG1sSTEyiZ/VJtT+vrU/5WlFkBJOHMZaH5gbEJ1sDex9uqng/ld
Zf5e+iUR4CPY3dnmw9HmwWtah0QaXhr4fg8gYjPfBsDzOEu+zmiVp9p80AVY514kTTq5X+edPd8l
a3koz/HfLPdeRa9GpozSmGlxzrHtB50DShHl6Cn8D9E9g0qMLWzyRDb3ylT0QvR2fvFqhA4pba6g
fG6Tzoj+1e+kBxrHM/JRb20kJqCATrKUQu1Ml4GZrAgbUjKjBhsHYoUYglS4RR5rQ8nWSvbxhwua
+9THGU/L1YgQnmmGlb3gfnHZ6h0OnCE5C4ZPcn3CJduB/G3U2/SvG0zdZXOAUB3KsTOnj403JI0l
YOz4Tis8r4nSX6/op0oaOlqy2MHbsF5Q952atsBrnyJx4Mn+eHMdC8Ots4PQAPthq43Fl57nVnlg
FY700vB9z2ovR4r5LsRIJYHwy/cWE01sNZwLDCZS7omuOLoMMIaHaRQNo3pf2mgGmMxHpGZpGCpr
afdmBI266tmwDYXV5aFRnQt3AqstwMCjBkc6Akoc+Ok4Knm4pFsjzNJG4S5B+Nx8bDVEGY1IUIpj
GMHFEdRaJ5haA9iCnxUI2+PwqsuztoN9BMOYgQpvRvVc/siHzEtUPQlBuluTk3GgbHJtV4ej+Ujp
1YovHCTQ8NV/ZaqLsx150LFVQBHkLj3XdbTFwsH0ppkjYPyTwK1AIUDEKSkInEjjfDr5QXQaTk1v
Oys9XpyIipYQVR4Inu1StHaMlJJdXt6lWCwZzulnpOJCl3cAesyoIN3T8TMYu8Zomcdn0zm8NWpG
TsguCgWrUGVe9JD80ys+oPA62P/9Y/9X0L12C6HUqeCNdgt5IhbL8duaLyeG2SkYL4Es4REYavFK
TNUpAxpJf+4FpgLaLmZUn2XmtkUD7akgyWYFlznrWKQ687Ws5lXUcVE4gTns+JfYRBBFNSYvWnGc
7sSiQyTFsCOKh+V++m30DruNq60abdS0KWoK3M8GA+leeKs68/kL99ZbIWGUGHPCo+dXg3Fonu9b
263dEIu2HnQThElNXUCksUyHBM74C1iOPvuHNV+SJKhJ16ZQkx06Oij1dcp55u4j4HUKh18e/NF6
lPS/D2s+kGIyvJSHRHX/9pPY9w3+RRQvUNxfUsf50xkuyAd2iQrIeNt9FzsTDVMqMq9Qk6ULQ5YX
O+iklL/HtyXoUHir7SVbOKXIw0D7WZIiwbxz88+uiXYA5KcKlhCRYNuSvnxsbQ4SsewRrIb4o6BW
G3JcI4vx26H6HZiL9Z2SHBVF8gN3AmvARZifWj1GuEHcZKsSdduHQpe69you75Hc7SH+piS4CpyI
R0oLXGa/gMwFkMjhFSlc0BSzz/s2OT8S7xX+U17FRiSuhzrLAvo9H2dNAFuoUDo/rtWjLi0zcjL5
27k2QT0BpOa8yD0eOhXkj95Psl4J0jQNAixPN1Ti+b+0jzN+snYRtSkm5yZElYhS+xzyDUC/wb37
+R0DYc+XVBtJ8tY1L/dpLbaheJzYa3XflH5JmVC4doGgcyn/wBxABf1z9oKkUx3s2IXzD9hPReY9
lZWgDyrObfmRpOnQlA+8QRsswlTCJgwbAo4iq2fKQ9dQQcVhlE1XgfxBOvYShb7orZJfTcAh/JZt
10baxC390hCDOA1ADGlFWdHQgUo91wLx44tO4d3bN3aeJaOP3M9IyLLjKbxECAhEpuzyNMQfLTZT
4V7LDjwNJUL17SNmyoSimcfwC4nat9zUvFH7ttzynblnSFrFveMR1rs2KMkK2g5KQDBqTFdIGaMt
fOqeqo/SHbtYCthKNWsEGr33kyQ3JQ3ijVtdzQfZcHtPqPqvcQvpkFxcgfu6zftKQ/N+XK4XUuj+
AFMUYL3fz0FJFWTT972uYw4uLS/nGZx+L1HLWzh2+MnyyWvG6+SUkkFxssbzg4HbQo5+Egc112SX
7NsJKhJucihXzp0gJJww4tz7pFgwpwNLCUoBxGFDTVZh3oJx8X6ewQ90npydlBZHAPqTQwM9OhAP
8wMkVBD9HxVQYky5v2jZVPYt3WkxbT6Wkpg6+bsknM9Ca7O4MRBbZzRWDy8je2mCfVULAL6uYLRl
HEPVm6e38EG7Hg1+RUmePA3tRoEa8zN56n2NzG4h3S209QVjukaUoKFsX+pNItThezEXH8oPKpxc
ha60dJAbmV1r2xuLvhw1Zo0gce0ynumVJ0YM57z72eqHoQTnaGpQ5aBHxOTIkWYvppisJ8sKoepk
F98RxI21CE4qulHgA7wS2XLtLihQ+uQA5aJII26LIYTML+ODu8CdcJAgGFh9xidO+/UG1S/IyfVz
+9vMxZkVOz9uV5qtAXcybFtovIhbdYL+gl8AsMMQtQeEn38Or4ZwgqneMykLW3a+VVFoHCRcGbgv
tKAIEgiBwVXjhMnB+hofqcUdJAaF6xwite93eTQBDXwezvuGPeOxGujYCh0ZMyvNqSNUQvMTN7Me
o4D1CEPzovJvYsKrSWJmrGthS0VmoV7Jgr4CHymsHZux5CQTH07vbUyAL2xESBGQga3/1emxiJS3
br5CWbzx6w3RgMKwwupuV077kScjfjZlIkxreHTm6d0izlDt/Um1kJ1cPp5MWY/OPoUxdhZfQsAN
JrYFMckaRBrxC9CVn33PV8lgfDvaQuApdKFtfaOzncFnnM4xLIsm982vzCjwGjOH12+jzEB7tHbj
3M9WCFZU92VZ1ZrFoMAbtDlbExKSMH8ds5VFXcHUXGXu47RsbdiIJc1+iQzK6RozerwC3tx3y5CN
KzAmXkFLXXQ8gS9z4qAJ/QcIgti4PyhosZLgZCA1kK19vYkTBSUr6aSboJmYgDrE7qt+GDNe5cxg
rC1W3xSZ4HmC3BCzZhn5RmoZHFHuJErsO9G/npGL5h1LcznWQkLh+Axzf78yI9GQznopvE+FNZQv
+TB9QafqGJajhNHetWoucL5WAVmI3FtvJGdQGo8hx9cWYO2lNeyOEXa+0ykl2QPfV5LeSyckDxHk
oOPeLnv/w8BJnaXYdVRVDhODN84Is2NnuXKsXgzSi1psjYDajvefHLN3wWM7GM9XzxYkj88PgVrY
KA/005N2wp1JI0eQMQAQ66j88cP1XBnH1eDWfgzG3N4lP9hZhyixfBlUjEzWpwm2cwX7SWzTedd2
Dw9pWTLVmRJRzmumw6ua72B83ddxkuPfbA5istVBjzx4iNFRydRk+9mKPAn0Y5Rf2N5jaZzOl6n1
BbsXHmt5E+wYUl8z7UZ1Y1J6xp6z6fmldpe/rU17DOq3eyapLljVWQNuq4TzRE10eIQO8MNDilIJ
AXh9tWRLOV57jLNRbNUzJmJDtNaV9DzZWXzqUzVFpd0EVSwNM4XRO2mYUNe5jgX7LAaZzQeVAbCv
fU9rYxv7nVBn6/+lJj/MvFvgIYLlDzHzBhN/EP7VqQET8Gz8my3Kb3ivPcU9QnvS88sgFyaKiGsC
zFEblWIx4YIM0giRyHwVs2wI5fZVs6dyCdU/RGUidWQQMFJ5tv66djNn/FzE1fm0T0udqDMTFaxC
dVS+UmZbZ5vqdT9eTjvNvgco2MwyBsg05IvrHzlnOWxeP0reJHOkNOsgRnFvb027P7YeyWeEkpR4
sty8BGhB9GLD9x8YZp4p904SEOgTNTEIQIplYTo6qeNwA9C/aKLVi4pH0H5As35xWMtJD5JPpsgt
iS18H9UOJuGkUvgSEkUEQ9hOfvEBhnTAGKj2EzelAODfIPbXrkK3IUUgZZeTRXcLXJ4ZVRnkOyQ5
PKSGb7RqK/r2sRsvu9hO729Y9qayBYF8btkACgJdhDs2yK13QXnfX0Jg5wTu31aiOOz0safJZbO6
U7y5p1spcqSfBEODof2DYFiGIhmJ2wgHkxYJbYoZF3LQIqpclGpDabFWgh0tOEoJas+NpM4qA5kn
F70ReLR0empyGw6SZREQEBnSWnQsXqFhgs+tGbOKdSguI7VeroxVgjdTeX2H33Kq3s2cl7nE8akS
ltr7ysfcXQD0LMpZKZvPB+nGBiyd/PBuyEV3b1VPk0F4fw+OFgxEtDae4c8zM3NKeibLYHRxY4a8
zJlKMvS0DEH40Y5mkbs625M8sgs4+wjlsSCo9IUnzUbOw10QoEOd2h0UxewvWxQOm/Hn1IOXpQKZ
JCFkBzUVPJS+LSxMHIDabdJ/N/Zqxmf/JX+EnUraxhtagI43dFBhmNYoDBvDr7GheC9PJHmYgpOj
DgfSkJaxCZyTiXO/W6IDgeV4E7cOnVR0RTkNwESuM7MZiOaZp//CtL/tQlaaSS4FcckG1lvufeHW
Sj4iFUcsHf63THrgboZRhAqFJ1g0sOhP5PC61U7kjpuOUMMxwNUS/6YWcJLSpRUNHbxa4SFAH9iO
Qvoxh6yXVJ+Utaey5/yhiXItfpYb8jTjfTK9BGv5nSWYSeQ3zGYWLyjkH4R8ZhRMnYpz+dSC8Zzd
qJGV6Rigc7JxgvMF/B1m472/tsPXMG8g78K2a5/tI3UzBVqS0s3HaVfaQr5bq8bsfkT6z6Xo3S6i
UfHzrGlyt8zhb66aPDnOFiMQHJncoDjmGBDatkCtevwhO5h3CdgTiGnl4i93HzffJep7roNDlb5/
h9tcg0to0eRinu/8ry6n/RmpYjbQMZ2n6j9Hc0Y9MPnCTwn/e+Ihl5cjPkiIU4gflR5F/Pt1swCH
TlbdW1DrWI4b/6XOrtYE9210wOa+c3ZnFKyafXnNHKhNEO/ne1UxTSAgMfEeA6xqqAOCt/HGCd9g
D3quME0L1BZ2U92F0+PQSWhYXsjG+YEFGQ2b4yOzzjAh6xqboV3sVjlPy7l6f8V1tGJWJbXaK5/y
pjRxsXEl41SVC9OrrU945UtsIFnTEL//Yr/JyTa3qy9ECAz017AF7tPV9Jt/o1rUROcuvwftRp19
baMfyo1eIBEbpVaIqo5/qlDjqgaqjq8FZ3s9m36VLWnZ+IjfNPZyEpW3gSrPiu+wMeMNkDdSTW4J
5x5QsGlXPJLXKAXTiO/XHtP5NRGDfx5vSyBpD3EbAPlRlpsk02ZhOliY8ZQY8pZIOt6a0LxgUQgJ
vYhJXPVhQLg+I7NWs1Ff+Rg3Id4YcHTMtCeSsC7/bHqp53SRomWUA1UlX9QkNS9dLvCtKLxrR45X
CFLXfj5XbAG78KuN4mVYQefwh1tx0Ty/iZ7K6c81eeHPRq+d43pEWYGFCFScjUwdkHTRmiUoQ7MR
YV0jDy7dnUPe3HY2sxDjxre24WoAW3DUH0AxOIihLIEKNdRKFx+7NEnJkClSre2WB866DpF2KPc9
aNOn+8Ka2cnTUAKRAtKEmK6Xz3Ki0lCEsaaylR8a9OOWi1lkK2GNYaLoJs8icpNLb0prQ1KR5uJ5
md909BiKyjy/mEAKKWT9P7uo52Hw8wWBsMGLVdhaw1VXKp7mD90egv6NroTjxhowyxKLbaxXZsau
2Ab96fiW+i0Fz01tl1C6IbRuyKH54NA22W5RLeQKf8Qvm3g5fzNed37h+G1eNuGAp7g7Whc5mUZ0
HdEOFOcuPHDq8tQPfbVH3UDGC2avQZ2EzzkYVpi7rGsOWQL5N3R49kn2xnvk//dHPNFu3jzkbLYF
9o6GXUKghmXsaSOlajCDmfR5SewZ5jaZne27DvdJ6FJw6nO2Xt/qcgBZTDJfpu533XjsojE6KlCb
1jpTok2ajvmiRRfZ8ey04cuylDgkecCQwXCGQZfyzG1vg1EVg4UbAvFr/VM/uZvCkXx1qRPQi5Ln
SbvLhXL8wVV/5ZZhQHOFJcLM+HA4DUCekuVPKkJkZ/J9jZCBtFqwgTGJTHtUF7Sms/Egu6DOhrvf
S116RdBNRVtQIXjmCGKOKgsom5sVObRSMmL+YAb0f6lkpZDCTvKpP/pYmrgJQ+cCxlDoS48Mamiu
8EL1oTCn3UeFVUZXpE8T/i/zSi3OKhLHEZSRpnDYetYWeUKvD+8Rkv4GPT5ymlkBpeRKcZiaw9kX
/Dcqk+GBwtTejaLGtD83USY3pzvcwja6gnwTcCi+qxgpmkgN6M8MF0Pjp6JkIPpnsmD0Ksd0U9ln
62BgJKBKcK9u0/PT+pf23hA/5pq2kjhmbnhNOdIM4U+jHnABg0zYqTVHiZ/cCGEYiMdAsfR7YTe4
Bm5+6+M+uhm3VUyFHujLaFrVE1zCIHfeVu1OFIkj4XsvWViAE68CPm9p8nCvxXVYI3pq7bnu3wX1
vYh/LphniYtHTG8KntPBHHCHk3ese2Bee92H7fopufL/zr5NgDDFQ8gnxUtY62EXnC71izpz0NU6
3vrEYEyZ0eVLCCKqy+6rZ+E78Dh+HZgfXkXlDcacyRVvXsMFXYly3xE5eVH1AmQHGRPFTySjiPUN
fUKuvo8sVurq0QzQYYu7c3lcwCAYIyVG8X2UT+SYNagesElQxUYeDfjlPr4z5PJiOG14Ry1wISBU
gzEVU8zj7nKTEGxIhHEY5Ads+uvEOqHcmjfujX+t1o2FWkuaa3diFuGOWevfWr4jtoWWu0Fa0klO
11n3mZqGw3OW5ydgglM0EuyxjX7SfDKudbuXKgkZP8qaDgWbpVBnIyQ54UwZR1CUGWORyiri7Axq
kaZp7oQlle0seZ/pqoP3lCqnTqHR3TO6tgT0mqRp6cPNJTCsPuHo9Phh6Wr9HW8aWxUa+YgfF4n1
/rHwnZPPRP0V3pBT4ETVh6vDVhqLZAX4EZQkdTCF3JVyyMLtfZ8NxSZ/JhWom2sGysoUUL+8oY5N
sgMuFERi01FccLagDWYSEbv/t21tAgkDzMzu2ZEGEJjKU9P3Wo+NLN9baqW77kjupQyfQBvoRSfP
F2Vg8JfFj6675DXRW+WP53CZgCE0q43pcUBaK1efS59AENo6XKGwRpoxKWqwGo4I09TZhUHgSrPl
+WCle8ZEET4DoRyEDpFJV6bh0WYiRhSejHZ2jUaR6RxUdALA5SbpJlD+WG4/C1fe+oDEmQGj46Px
CotRlz4MMf8WNB6xNraJvH/2GxqYYv9/0Nj8glp5j2esXhhEVAs8NaVu+7fS9oQ1MLw+eT6IG/QO
ISJhGlzk9fNaPi7h1/wnyY9+lSOOkdJuvMUkulFjgLAHhT3530u4OLcJ+FBSfwP6LABWcwnieu0n
dUxo8R+7vcIfnfYioqUyYTDDVuTpCFtKqJGhkYR6WTNTPRVQ6XHcORi4yzMEhVBYFZMFOWDlsW9L
0ETKThSL9g+QjA64YTTO1TSTusFz1/RDwplYK8oJ3MapWkHWY4EGmdtrSAfsJ2AilQ0rjkwsbLIf
RMSjdZLSFzAHAOtaY5EBCHY+MDH4G6fHNJBCxd7s9icbxrKowfrIeSGPgNz1LXlPgifAQ4VpGM1H
irbapbglEJwYu+cMHzWxVhIU5zEjcbTULzZyAnUoQvGENirC2KWzGGAf7f3jEvuEzVMvF7JqTRNU
lCdt8lvf5U1Wdm2lSk6+uA9kIsMqR+/dUFQnqOPGj79WX8PfwkBdgJl72p2rbulSf1R8eyWznjxi
Qza6KmXGDZBWxMi+gWUluUKszCcYmtiMJ6kkQr+FnJr+1wPR2RW21/YKd5Bb5xpCX4J85N7k3EsC
/xB9BriA/1rQBcj7VgVJM2+VPNYBJvk/y0PFXSRaojeph0GEYjtr8ylnIPUBKUK3NoeSGwDqFdpR
6/PsYAXcAG42r999qB9L9VM7xRPH08uAWgaim2pXMrTt2jJAsmc1KRIQr/Em4Il9R0BCqcorVDB1
2QNHWjRIcg7cFPABsUFjHYD0JVSz94OkHc2m1gZZKR+eSpxPBfUQhCyxrt67pN+vmMGoo9DlMA51
XYciLi+3qEbGqaGzkqe/KvPYP1R1Aa0YmpBXfnue0K8QhGWFKGiztFabXu9+CWyIxFm3UkP2BwSw
ZNv9SRRhPvgNiJDgJ5huK9EmQ5vR+yphrH/jUW31Xzazlp/yC79NZ4spsQwQgLe/uCyrSg1XPLIf
QgPzr6dMQk/mWmCoGGdj/jUn/dirAjmrovNpZdsDNfeqggEzjAvOw/nh2CN03AkGh68LeWiw79uR
ZfHLSe6HdC+Gqc2sAHAPPrt5KNahnPvDCXpRs1OL9HYuWfm+kD6xtkruJj0nhIh85oQx+Zd5FJoH
jIpUpz3hY4OKKenLqaSaI8KIgyQKwhRFSunBtomJKEUFiClhRdw+tfQ8pn/XmWp553BDVNjzA4eT
3aTzbXel7aToGluc/Frk9IVuX2jUkKM7MH2TzOFc/bH21dJLV3eRqZDywwPDWHThS9MMAIV/rUOl
gmxSLiRzlLjdCT2NFsP8+m9It+5vu0uCJQm0TDwc1V74o+WhkjRT0sazg9etOrC1U4wKM3qwusfn
XuyNpIOcZFUloEh5DMGFAty/r2rTOZnHaRvoMus3xV0z6XSHV8XJW2Oy17eBWgwVv/12Hk5xoDIm
eHV36pGLRvIAY7rHpiRNUCZE2baSWzKPNOtJFDi7f2XHZsPX2lGRfv1/PlU7rpQyrtAUQLN1xdH0
UB0kzvOUE/TKe612Ce/SwWxeTj/WxWbZOWx1d8b0hnhhhqcGrGbBsbL2NkeKSuliN7lwG/qIGLmg
frZrXMnvop/FNhlmgNT8QD3skDeZXWPAOE9dHsFhAnWzEKGMcU+zHY0vme7Ei46x5jRPYrljB+Tp
xUY6WuNlgYJEug36K3oIRo0InHShGHmv6N8vNk3bQ+V7BQLcXUmDfeKNfbs1sfp226TTlD/DKIz0
9aCfhmUcLDlHawaajGn3LK0hvG2l1IB8J4RUn0c7BzcsuDX5dMRpa4hDi1nJ4GUQ3wG/K4RUSir9
hm5N4bZVN5iyBOT6oy16M24XiQ36BlTcygKyCn3UF6P8/GlsM5pkaotjoJhC3gmM7kKVMIUAov1G
SRZu34Kaz99gV1JbJm5vvAFiKvj6Dx65d78RTOIeAaXLcgjNI8U3fpB6t0s+iVpMSnEHZjmoYxKw
1JCZ8VDx5FHAGepjSSg1ywoRoEwFw9PDdzk9lwMpDQREoJs5q+sIb42CKpGGOfevmaVKDBHmsJjj
BzZb0anmzmpHmltFu8DC72dma6FrpZg4hgvswP37wu2/YCc9BAQ0qnWTQs15rypB9hAWUMMh+brH
9b/riOrSemahGl1kEQE6gNXwTIhe3z+crtW4zFdBZ6Ue7n/Fwo5WiE54KxtigJjEcrclk/RQ0edQ
fynYobXfLWGNuKKw04TA6EXmSS4iiTmCC8+Rkuwc3x/fyTjnvO6St1Jv8NIzcKlZElZvCIaJws3Q
Mg4MUKM7cXMZ54WMOe+VEZ+X4t7XSJnnDdliHhDbpAX6Kbc+ec/YQiUR5ZahySAbLWw73Wh1BwQd
+75WQ53PgkmyzMBwhWtLm0h69k0VPrbYKJfmhpcDWZ/SWTL9QG248P1Hs2Xj0y55u9l1OROcyp4j
xpgXyBeerOku6ppkaWHEu2I2BCWLyxHzEMplSE08asDSDjKG9t+yEZkgfNfjnzljeZrUmNW5QxnS
kNQjH6BORGU7/MAqw4avl05aO4ignb0ZP/Ig1YopGdXkAP8UctUiKlFNNEqx27UrF/xd6/5T+lwT
Iw0FWeQQ6znP7mKiADyOteqD6Cwxd27gcKoV36Rz6stEWg4n2bYtqnU+nQX+SHqz30kmSa8YXB7E
et1f1BjkG6w9FrAm/KTQt0zuS2/aC60jhuAFiuXFjwQXTmGOYF3X0ZB4MrbJcypVrBoTPMyeexaH
Ll8J5ie8V/aXiuX9UkEKA0uv8JZ2qlGn9zkZXErq+JMOoDsUuzaUTySICyYK3eA5y2geFkgJf+qU
Wg8gj7i2+ebBCFf1WVXkIKn55G7Bh9eATK4pcPml7ts2fiI1Ts6UW86gRtE2iLJd3foe6kaNG78G
lUicXusVbR3xwHTK4/i0Z+mq0fe8uFk9TIbzxp+Yl9E2t9Z694F0VGveY7WudElJR3Am1me19XY3
w8wAYt/xuvtfq1LWMUIRNaR1a6lNk0jutTm4lT/ZuUv8e1QYB9pzqxlhrnpvxo346W1h1TsmvlVc
VCaYfyXz+dZkoQ4s/veP4iRWQE1VJPzRtBtLj8u97tlUtZ+GNS/VYVFUZ5Rx37wYaq6f4eTGLURS
dLtOVGh5EETa1MWNC3/WkYium5ngru47AVd6U+jRiw5d6kocni+H3h6s3mESOqOay49+1tN0jbio
GCnENnb2EWiqqBin1kY2y8PfTODYET1SL4mFqB9Krgw+01FRbUFxUZ/0c/XmTzMm21M1uuj81wDf
lp0RTDwS3oeBTVag0LPQBWbOCrfWmd0Rxul/FptVL0i+hmaZCsYsLgEd19A/RkkVQ4q501O3B78V
XvZFe04tpLbj1s6ZTH4CAWACeMji1VA3dgX2LMzn4Uc5m4ruW2lpOTpOC29HMwmze/T2HpNrdAOF
APee4R5/A5AkcI3lVNrFmyLBC+PF9JOkOaDx1sQOfSojHmWmKeWfnfyTiXCh4zI4CRdO+7ifkMYR
sH4RsEZXgY1oni5OCSL6gw+M/carlRoM+XCvkg+Iq1FFqd59AtBjs5sCGRDULGoM3AiHztf5iitP
G4KksFh6p9vQMXHJccQF2GVHziFkI8BpaM+8Rkzm1uFQeyx2lpRMSu3DSQDbC5IjuuHnff+MZbOf
q5EAzIN2rFlx1wg5MpmLZW34Dsy2eWckUG1T5uzt61m6MIHFROPxXNrXgAtbrSotpiWjRxEBn+Ur
lBtj4iVEUOlnTEmS5rhp1lXs42S5GW56pj/NlZTQ/xm9csvmFUYY536ufq2XwYq40mndB5oOnM+E
vmLMUyUXlQlTWLP9YTS3YDBB/JHIjcFPDy7fnzUnP7Zl6rI8eWP09i3oaO/MMGfaIp4o4MgU6/gA
IwZRzuSxY3KmM6yOd4w7tYFyhjX5yU21TpOVKq1Lt/T3/D1KxLSnrpKvOy2c/0a62MM3mfb1tHy0
OsJlijg7DcCutmjvJb4Ff/BBRA1tGSD6oaI55giuGBptRY25UYqsRWt7Vomne2hxXV0gAF3v+gM+
pek2wK0hZ3UZKzA3h8VHqaLpKLe6cLNoca1XQhW9doTSOEzTFlWue1sRrysq6+AZjWtZ2mqii6jd
S1koC4Zc2WYyxSrw7ScS/3JP3reQw/th6ZDJpbJDvZVjKbK6r/TrzsPE6sqAPOKte+gPShkxWs3B
DBb16PJC/2yeKo8VKMPh92uwHPo5N1q9L3yBUV0Z/ohmSR8cI1oYShLbGp+sHb+4kPcvUdM93/C3
77itkVkfl7AXK3DbH9Y3JZZL4FJyZwrxo2C5F1yM2uzs9xnOu1pjZSHK20d0oN57Dl/52GFz+x4l
xQfg0bYFf63QhBKZNsdLHO28SqtESpJszu1rzNkOp7mVMPkW2lsbdE+czalWY7oI4Ki/sSwUYrDh
ygpEBaoN8d1hGGv98fKbaSDQLoCl3atKwAtdpH713yib9ZALduzl/tjs2LCRzjgRlN1Yok4Ph5ky
t+g8O6j/ZejQo2BVt9kw2E0mw+/orNw/Z/W/VQ+QcFBfgedEznCM/hqqg4FGUXmOl9uY5yDmllFi
KaajS30qtk6pFXVuPjkybWhQ5C8lSLRYx4kFU1hq0DrB+xGDvGAfNUV1wqr6GE5RabziXr94kVa9
0PlqV/9nZrSJfi+tacpMvTtuS8BV3u4Alata0DpSklh5Opv01KfDeIWdLGGo7SarhxihbAMjg2xY
geOdV7YDRmIRTZrytIkrCsln70XrhpTjA/B2ZrJBDqyuhK5yBTZmAsYaKyFiFNCBrFC9HExQO+U8
UxUQpQG99z/5oUQcG+Xfhpvwumn5EjyCuh7iEagnCFq7CAPTVAm0HeZptQa9cSZUs1GuqqGMD/cu
h+GLvG+CO8GdQpbpPWdKft+2U+yc6+nuqweT6nyN5aHFISY/lZ255pg0tcgwjnGEtY2/NoKYRKCU
QB8sOzlWaLlVKfZA5Pmu1SVn8PmDTK7MgPVEE3syvXrWdFc86mBPtuZ0ip/11YZ+YZLepjhDFMGk
uovY9z4Oj+AwgesHzw1G9U37PWpTXUhH3uzWDepMddAD7yNVWmiB0i1pWskYEhxKWGAOgXguHyip
lLF9h2SNhW1eLbG2kuL2w9uwmWcDkRgLdDg/aOJrbe2zg2DYRfHl9rvNMBHdqZwjyQLDqwjEeOb8
jyuIZRRn1MNW2p/+d7x3K023N0eXaVbxaNkZ3r1DtzuGofepTbHNTZiKDBk8cjBknMNtqGFynAan
huvtevgSWxtQUYBX9rQnhrTlf8cxCqtYXflpBJDbqCVHXSxzrcu+A9o/Ja8L87KJsGuszK48NHC+
YGDAPxnxI8/LM+hVUcwZFo/JvppQ7NTJwEK6eQ5Adfo4TMxx+OYAWm2SuUHTShDKd4WbejSsQWML
CHoNPPFR8pfrkJY3n0MiC1AGNcIA9ZWwhVR+RCyXibAeIq16nU4LXrCS9fI6xXXV98UASMxm4abb
hYiwFBPN4pSBh4Sb/ZQZA+OGhCU+8nv1ysHGhs/z8eTVaP1nMjUdUNAr2BzU6StXRlwXF/2xS4uf
1KZ8hLk1JAa0MKVfd12DWN9InNDMf/rnJ/Tce1Lf/IY11fV6oEYq96uwCSVv6EX4RON8agxge3Ib
2jS0ZIgtebwqkw+1ZpWs4Lp1YaqCm+0aoGRp1jZuv+5jmqTzmnPOXjtE6TCw91sldglde4qyk9yu
jo5SchCpCDwCutGZMNUqeD6urzgZREXhNKiVDU67c4e595eEE8dX0OQ+HoLK3Q+IiMtUUfB6ed3W
DpgPOhqR/se6PwU6Rc7UlITyfO0ZE4x0kFtOJsNTybB6e1XY9JtUg7GRubosuKH/J5hcxDz7+Da6
Ie2D21Ql4ZHyjM5LWDJjrpvj/qXWObOJ7w9M+/rL439BoBYIxleksGMeLUqNHlS2FGNu9RRQZB2b
J7JrV05z5mn1dAApn1mf+DZ1bomShJ+EstPHOEblM5Kp18k8oSW5YUfHtBgOjIbpkyHAzP4KGOja
m/TgEeCjbaWK7CV/TYaHS7MkLa8TmT9r+5cGSJrO+Rr6aMgri+K2MkmhDESwp+OTC559JnOkn4un
wSXtmT6KWmyOsVNeph5VyKKWF2uWzuer9qO2dQeXn3RnwhVlN+IwOtO3zG/rGXiu+izq+ZVKu259
894iWxYUjFaE2NfmXfRI1+K7Tl4xuDBQIoRe1ahs0GL3UYbZWmOW2p2sHJjTdt+vKp2gOD57l56u
tDdC3r/HkTn8zBPiwpbSYGsNGvq5+sXeoVBDj8dodgdvBWW1vPb8n53HUubBqnNhiEwNXRjtzsnz
TJSdD5e/HNzOIq1Jh1H7IiacnbL38yEdWrf7UtxxlCyL5etWjP6lH7kYjrNzcwjndzK7dC3fWgRn
2eV8l+QdO6w9YEY6HluuM7GQCSL2jHx5My39hGwXCJ62I7lq/ofF0pMNgA3AJnvDH+YnYIXJbyQz
OZQ9XUEC9r4atWK/3DtnaaRkErK2kz2HuXLasthILXzPRnqwIJa873W6DWcZkIn/ckIFsoUKa+d+
6HVRnjrvueWkKqh1jX3MKeKf65prQDXoaT42keJl7yoyXGchrWCn8cSe2iwc8UnT644cvzVA8iVz
hwJfHyZD1F0r4hXWBpJTaIam0ib+VAZC3BjmQU6dV8YMas9UEKSaIFkXFwC3v7uCBShHFoulvQbp
eGO9HyK3oADUN707Cx5fZD7osw35muU87sjNuzCSr8YbES5ihkO+AaFFGeawHjTFPaI9KDRAEPsr
FRWhq5L32NpfNEd0x+1gn6vS2u1cpFHP6CA8M57FOW7mof9PKRiNYI7hqkwJk08feRQ3g9qkau/8
LWBc4Hz0VL7GF66xyN3Y30ocYXfv6aJfFOjbS+So0GhdTT8/xjwQM6/EUp3tC+kcdw3hzUziaU/0
wo4KGSKjHLKfxYXmFzmpEPo96jT3iQ2+nB3QjNfk8WjR8Um9hIDFsBG3DaBTR/UPnZk25vvhggzO
QsPu8Mw0mZ9LDDS4nGD59Qx+sCVuL08qo1Q7rQNUMhxONk04KS7Rak5KebQlSdo0d3KXPFQaIeAt
W6Fzqxtq2qaLGDn14zSJLbYaD4gWS5ssB53+1zb0yWwG+PSEGbtpim4A3pauOgUFWpMKZM/EwNNA
FZ1kV2YoDIGJxBT+pjqIcGAWT1Il+rKEccFU123sfmiBmoXLyYzu/Cz5ueU1iUGYWCzXiYbU4aQg
Lf7Xm5Omeve9kkqReQDo30NQc0KAiSJ/zDf0oaa37Af+dOxDyYu7BVAtIAuwyVaYLstBtz909Ck1
YEvetewR0hZBB7rC+CVwpAjkM9Q76wzlJJEXC9AOCJUF/PvB7XYwUY5zkXzoqVz1zKqQefWvfMW4
Y56tPRus5BW1/QqAyvDjEWXjAXUbTbYbVz64tOF6ib3s4y5Z9Z5mP6WvhWcoC4VK+mh3VeZyp9Cw
9wkKGu0oICUylL8HM+MYGnFfE7ZkGi3XrEEF4mcpjIBYoS+BdXXDOQ+c9rQgkehp+fT7xbQU9rC/
AaR1J++OvxiAnkYV2mPOc05OQrppEjWlYjFvNKPYBNsEz9+GUJmT/LmFZ7xNEeCTbDq8OJXVCxOv
o8T1Vje3oWbYRP+ew3KZLvrU/htocCowfvByL/hQCA74CCnR4LlY8fCiHZ7c0yM32oTNZE09SEcF
y8qBEipEEMPMrNec9lI/zhHCp/a390aFGsvgq66ZYBrOe3UH/GQ4Ded9x4BWsb0+8q/xAFuSpzUL
2mrXzkONdkpaKU3tnd1Fm+pVQcf3/xAsX7J2S6GbiZzonkctKgxNyf5um57QXh8Ao+AvAB3ObrXT
+DEL4rHSa9fk5CmirMv+Kf/jAWwE7D8k9DJnzybLl6VGxy5/NAO8w1n5Kjxa9Ctw/xR1XFss76za
eRKDMbK5jOsKrVdVPYZrEFBsmb8sRqDgVPtG1Aca+2IryA4/EUlof7EZvycmzI8uwRHnVk7mReDg
nMra6ZAIhwYTR2tukInBdiElv8Bny0N2SnNu6/FH8m7lVIVE/3uC/iz/Cn88rTlcrXIIrUe1Nawm
q1BPo3ydmFE/t7feSSQzYF4O7h9/v4ZiZtJ95BoImE9rf1Jr8gxj3bOFxhHmfbHjCfims+DaKRZF
3y16n83baDlk367lH4Cjgi0Fp+U5UnbZJ790Hs9BEItDb/xGxu2iMk9vJx7dqK3+01SB6uMfZpr6
H80EZPNDVVvf2je4cGa/KVq5DtAUtwEVu6d2+tiD//sr2Cyep3sB7dN1JfylXGQob481AWmrTOxE
VuB12+5fQyGuIiCi0ajAC9OeqtU52cKDrwaFBKushZTlQiOoEdRnLF/CdGRg3TbRx37L16ItnkqA
HfxhAMQ8V9k0YGnHDGDCx3D5k0kbHe/5rRNOjHCrgczTXjGSvZ3jHjki3z13R66LF6bTr1fa9Ose
EhH4jOgz3H835PbpxT3HJI1kD/mW6ibTY34dpSXb3Z0XFep0ZqUGdUfyFSfjVN9ukXR7Xw9ql5gy
Wy0XNjGmnqljJeXRtpQCAMadFckJWqvBC+oMkFs0NElbAxAF1lX2vOJYPJJTSrfDUHznQajb4rkO
BTbIPR1DITsRERqYWzQNlJTn9RJQ4ZN6FDai436ZVH0FW9h4fzTjyLa2dN2N9oDBKrwgp/uvVm0S
xWV/82Dj852Kqpy/pCnxB5qbxb2GC/h29+oo8Il64gAlxfMho327IBngDHTqeiEFzjLZu4I2ytHh
b8k5iXbKc2Qa72vkNIU3JD21dyAH3/wFJKyjIAwD7wLy3zZrnLtLrjC0vKVAzLZ0ZpdHX7Lztp7F
AIYdX8aUBSDz+qN1Lkv4yjPCpPtYsmn/ii7wbmtCrkbbNB3woaMsRFshldX+xQqD6TelGgyImX1z
3gPNRLjexgVBdc7sIqToT0Ah+A/QL3SXAdZlnVqGnDrsOb8T6CZDyyBpjtxyTOuzhGxJ7/TnD72B
DC2B3ZYB89I/p/EMzg/cMxtcxSYcF7k+0aljUR5VzROD/vAG70IOkgum7JsBF42qaWxS734TJpdb
CAoOhHNLjSgVNjjDnsSU41qlJBXAKCWuOitBKYO/WbddiyH7Lu/Rfoprvlg8+Yt5Bv+vg/CR8p7A
c/in+Pe0pyJnF+DpdcpntZB7sUvspWc+h03ZduVqUbfIAZTrhsR6uXY7Dh/mPW2UEsZT30X69YGU
50IgkqsZ1S6fUbY2dpnOA5RmDnkKPzN+jwmzRtKY/P+KzFTKiMCQj7mNf3xDe7IPxx1GwOSWmphM
f2/uH1hDgmXn9zoM+XE4FqAp/RlFcBkMYEDnqs1V0P9zfij7G1Cc4RHTslOjZOVl8WhnPD8UP7k3
8jzTmU6JNzggcNfZsVCoipHg0UdNeFz18Ojk7RXOgid1gFMqr6fDZdj3ma3XxCzPB9zghl/Aj0cj
x4R9WBPoNkm32qBGpvF3mjWd7YY1HF6Iva5/sYZt5NwOaNTdeNIEb/1piJZxCjSru+iT+OHmZJD+
R7Y/m6kXIesHG6LNYXKamK/gPOPWiZYq8tqULFgxfRHlQxh1xxwXMRrBw/xA2bF8XE6doyeEteX/
Ma+DdCiviHfLvjn31noaSWAj46VDJRrnovy72veL0YV14rQGfligL7zhsm6DH1kGOzH4UgCmozmj
PON1OefD7K1G2rRJzlPKKLo3NLMvy+F2cDeD9I3VNM1Uor7lRodaW41p5uaTDacIQ/wEWOkIYLMC
ek0DLg5DNuyF+zIHL6C9kw0gLCJQm0glqmPabqkpoOEEg1+IhakLvgYuABZ3rf3YWA9cV+nLwhub
A3mNN2b/mmk7eGJ6EMwASI5hVsI/RQ0QapIsZnZfK1wzUydKO7VA49qBCX1fAmIRuzzWO0VthDhk
m2EdR/+PPcC+3Z6OItSZ8K5h02gLVK73ZV5i1b1TzIFFupnllz/L/WdHf55R8kObZmoPlGu14oQn
skN8LQFLvZakwf9GIjWqJAjvzHUWK+vF8ppsqQqAkLdCdk2uIK+J7e3Wl6mU3XJqmL4APRnNGF0o
HjmADyYdmn3GGhRK6kPcnw9InHo7cfZY2toYX0dzoYp5gmwpUKQPyhyU5KSrz+noP62RRTCFvpeG
0gqnzqeLt6Ympn8gZW5PZZZcivIb1FScKhhzB9d0aUFTiTXorvBvK8h2a/yKrEP8MJBdt+6pSkQ+
h4bcAPAnRT0PkjaSVvY8ueCbHD60IJOm+X0w8CqP9dyz5FckvM2IO3VD9h16hih5U7hwOKnVRUt6
jH5o8YmZO0P8YuRLTouE1fryFzCReQjiwJAeKt5FfsaRLqZ1h25Gwsd/lpCBWXebQju6ymAA3rPm
3dhOJONXNu64LAtwtJvxS8P+Qlnx30Qd3GBltghM2BVjrD34x4OmqNAhMkjrU9rse2oxk5qJ0z8l
Xk+QXnCLF43bbcC+OK8l9xkNVy7a3nwerTlI8IVgezBu4Zyqer209LnPtfFFBeIB7SFERxvaJOmG
E/2jCAKYdIqYZbsU7ugej8fClJqnB+rI6qsENUdSF/P50Y1IzgUPBXJm8IpjdlH82Eo50xw9A95V
AwdM31AAEseJJ9IGYxTQAaO31RvppiApGvxXgFjSSohibL12OKezRICdnOcbAcYPoksE3ZG6Rcy/
A8OC5FTxFPkW8frDEKObMv4h1Du3zikIpC+Sh/HnzqEA1hur+bbc4MVORTCaWg7ToMZlL1MWsnmO
LzCa4/hHu3jTH2Snx7bPMRhnTy0yndOjxfaZCZzv5JNOGwc12SRCozTh0eRJ/4AqwzWKSLaDNocm
4RlQ6GFEGeBBzSX6FgjSt/utA0mqilIjLRVaJCfKNiqrEZXYqnAyOdKUbYGoVSA1d2aees9E+NpP
wGBiRaD/rNCotNaX1+AWg0y60wmD5IAoRWtuvVjdw7CZZbIsiO5JjGWpUL9JXJ71VYd2ZMP+Vez0
RHYdK+XN8nZdE/o1c0plsecokW7Ks0FOklKYPPrkUcHPwtSGACkOlH/uNqVq6qiD8ryyAD0D7LbX
j494HvfQETfzgtJ1H9VJ6WHYpLnbmk4gTurLxXVB9G+uLMHoah6b20oGmR0OZjCC0Go8zR24Gl20
zjaA8U6Ev0pNffZD+4vLy/lrZfZJNjiWbGeyEHnZ1f0fJXyX61WT6wh+9Fj0J6gfdE7nst67c7gl
wN5K4XFvIxx4PCGd9v2b87IqZ6+HVj6lu1H7bv80r2pRXtVkhkJ/Ywf+SBbt/YB4+eIEqOEjrnoS
IF6dBjUKBaRjYzoDKNv/wZuLr8H03RcNotqEEtJo60mZvie7TK3z8AmHaJ0E+r37LJlBLHylj8Fi
+5FiQMNu8e0aAeY+I8rTDOHcPs6iFfVieq3GcecYVyplE7K+ac256J0GY1Cp+jGqEB3H0nl9MvHC
K8Umq4+lmXOf5Tm7Pe9SmLsRez6pcB40bWTuqrZkWeEUa9mhOLe0NRKxAaMqeHNci7PShel0y7vI
oFvPK120bzZrRMQs9YR/KMrzryDz2qbWJ6Adk3h+EtrNzgG3CocuUAnB4FCNYuX49UZO5b0jQaHq
xsObFq8PlgJsxsGKJOyfrriIxgZVBBND4+tp7yrbmQIkScPPGAnnKgIUa+Imk2p1HNjBPfhT6/0Y
M5gVetOjA+IznqdvLuff2hwkNlZXtWCOLkVxa7uPp7hXxJaq4NtvewBfV4pcJfh+u8+5lFIiyHaN
hkniOIYP0jHQzDBk9tT8RwmcqKQ9oAy5hMEKRIvhoaPH7khzqgIc+F1fFjAcYDkS5joKbkHL2TxA
EnaaDetLqrxWOPOmVx3ofUBKiOJkiHyv7IwBw3468M0XT6S3QkvsIAnXUNqZ37CwaID84aYk9Xme
6suF0uFB2/fPaVD5DP+yOwYFwpORb6XCyVVBC3I54i2HzuWUUicHdt0sAfG7K62i919U2HyNNp6Z
z4haP2yN1BsoMgKxZea4XK991Fo46QbVsISNUTnkYl1Y9Oyvct1fmgKNFCvcgCouTYoXdt1EaCES
8gtiHupeNDKwZfo/zgi1UliH0iiSZj6dOHcWwY+RHPIOG8ABgG/v6+wrW525cYeYAqAOWdOXQp2b
xtICpwC2447se69HWZS4XZZxP4J/Y75wdWe6nJsfyusjngiNQBgn8IwRvV/8/HFYEpP5JVCJP74/
YFlEhWH1Z5dS/sdUrUskekpp41+XDnZ8mGeGSdwdGG0O+BzBAOUcv7sxe9l6JcmGLqvnj+Qm3grS
YZaJ45dFy6OtnRtRExNUV4fcBqoo0MXcc/WtzbnO+or+2rrPn9gFrlnPbiLmSP+5Tg7G4LNuz6i0
pj/NHI+TdJ4jOEPR0VrWrDt9uEOs1xZazTePrjFh/H1p+LVsMeLZtPlq7+w5dqfKzsq0uvsuoH5Q
3VmkDj5P8IZlTIFkHsbqBc8cGXPIoehGNxObL5H9JFHdOxzQKvnd1O5Bpyjr1Ky+r84asgm7HVTz
oLCi7QVWPywUibzASjDE3k/fVItidk3gdEuaz3knEwegdntCtHUCzDldAWVRS0WGAbnJrvXStdPk
5lGvUosvvDnBN0N0/ghiiXd1Fqz/2j/8oEWi3d+SulAu4DibiQ/oix5nTUKV0LOg9Wpd/4rQHwz7
7jDPzqblgcI1pmyuRIgYPDrDakFop/W6cdIfKIyQb3ZWdpxkVjiV2YQzsEN6DMQTC4wAtOPMtFN4
3NpSYLEpDVAfcZlE25riBsMKQ7eg3VSmPWTrFEVv20oL864pteshb4SFuFT6r/MA62I23g50kgr7
cQFQ9k5Epgih2bfKzK4YR07A+2dwJ5Ydn8deTXTcI3GHiGh5zcW91F+dCHHdgdhhK0f1JSmCBH0T
gFLjVzg+fXanSetgXh/SwZiS+FlX+QPZM7vfzZ6kqQBLq30pzNSepV3dF9pdE5esxvPdNmIT+FfF
Ox+9336ZS10VAbsbtWcDbbqW1TcKFYHQuVdyo1eqgM5rSZ4mFJridVhn/euutbsFr3zCqMlV0X9u
3660+H762F5WDLnZORKk9b8hx/EmzYM1Ee10kqQcFzpeIs0O5othwnRlupts25O9dXAjf3c/ROtV
lH2UeMpEqt2puQFgcGznOhGw7zRRZB03MCAxuy6H1/muHXk1QNi42vhSoq8WNevGwnsmlPvJmDs7
Qk7R7Qls5aBr2J+IBdcWtFJ16P3+KyMCqYWJqrm2ah+IdSsTF24Pn0wWkTftEo9+wv4ae1qXIBPN
dxTeZY1DWbUVaJvLOBWSQpCpJTdzrvx3Hbkqi3HWw6EIxmf4ZadVdSEJLyjxy7EuVj50M0LoydAb
PRiASC9FlxXmQiuMDXPfYLjI9fY9yC13k4rxkt3aGpbhtzWxwkcxx4B57UbH6x93YNpOz0fdHftW
+YzuL/zonI00/ZiNb/RvkxhsqARWFcFMYUsDIzkCxoo0Y79rvNLly5kKj4hlzz41Hu3demgPKKrq
SzibOBgdB7H0yP++k4q0Y9pTmQoR6u5EjRmzoZ4/a16Yd0JB7c8NNHKpc15hiW2ePSTcsIEh7A6y
xaOpad+NkVjRUxbnbXDh33L4vEI/KGtvsG71Wr7hSEU3QeGBBCqAOPTq99uLNJ72DKXw4b9mYETh
gQyZg9Qq8xaocBnEybzDvCS86TtH4sGkuHQI/xru8gQhSUtDD2ofKN+5zwe9xDzK3IV2m3f+aPn6
Bca/492PPk3jqFFs72WFHNcN0VMfzzCrI7W0pyqTD7+HBrNzwvRlHbdR584b3Od/oOE7Ua56saa6
TAni9JcGM7dSG+76Pjwn3cJJOVVyiEPVl+ZlsdQf8NYD8khQPThoQxV2OhCQvMy9pAsHzOQZuSWZ
mn+boyDTgfJkEvQjCsxB5javpjbtEwBbZz7/KqUNe/iE9PtcX4l+Zm5Bk0g/C1lo0irtSYHAXMzZ
ZHX/ZDNF7EjYv4yWJnF73nV8KWyNekhgJR/vuPylcQWqo5+oZs/tE21oy5uw7hPbWdThirBuDUQk
1RmyTJ8zce7/Wbjidad/2GNRKe0SzwagzxYUabx6veRLIn6/fNuU40ezVILZXPViLJmkua8Fzw+/
/ZyF6unSCzx32JhmcZND3qc0ms9lv9ZSP7p3W7uA2Fg9VfnHY2Ed6sV4NhZ+KQw7n58pC6k3PZZx
JfYciqMPkIgsYm5sLfaVTvK61TBRRcXqVl/jM4uhgLSzutTRMNihh6lXNoLHiPKmoOEvLG5X4CjO
3roShsgNm5IugJjcHn9mlmbWIKNEHkLPJ5tD/dAkdtqDuxNDfn9m/btgHvPhFqEsfW4JB7PO+RcQ
nvFGF/GIYNoe97iakhi0jl4f47A/zqVwRUDKU8MGWAKjkSOF+mKs2YIMaXQ1hS1qq7cn/7DEiJ7k
0YRyW1ZYgXHS1z/CqeqVWZUk1bkuNgf+cq4xGb4cB8YOEs4oXmxTx0FMycoxp2uHbO8xgoxTf+Ua
18xMjcOnTfjKUUStf3i/WZFIYcw1DS7B0pXYaa0bhrqYiKSxKsj367vKuVgwOyWJyQp/8DI+hzWy
pM2kQIDSjfBZ2IEfn+VKtHCm4tp1NemBnBLWalcDuwmvMlVW8kwUVzMely1b1wNzl/jkD9e5haZf
pQL7Z68AqUfMMbxAAANxS6l7vIjyChsflT48mujAXfCOHhZ3ABz+aGjs0CYIH/RKhxtbcZQYpjzl
4xgSYxFoKeB/wEKRjOO46S3MVeku0/gSMiFTqc2ykT8WevtOIk+1+MFSTh2739MlxLmuHmRaQ05H
XKFcSiCoHOIC1G6lopil1izeXw9mMcf9+GCATiICBba2dwVTleYTcwRfZcZ2MabS8wXMwftJpZQK
B80pUpa3tldZjkv99tg1lYrRcrizAebqF7oa0tPfELaUih5BC9XkFVmuejNtSU4mHNrKRaJiid89
DefJlcno0drNhiysit/Codwl4eulaE/15bteeaRxpKqa6/4eMdPZ7h5YNernKQhUcRAf7gr/w5vA
AotcA4yLiADqABeG+NZsdQDdsCuGlGyYi3zS/68dMyoqO4ZLChMYzO9DG41VJFPioZkO2wPBdPDP
ENJYuoGEvTgVvyE2BbboLNlLhHBuxIg34lLMbjEglkpRmNtXPTDfqjwmnFPuTzZptOJDDOY0Ca7q
AMIqTO27E6BxpStWEpPGHCJYpVH0FhdjrlI6Lvptjgw1MEcYCpf/9m1eJAWBGjlhlbGQQSC/3tbw
DBOsl4MJ/9w23zlc9w9VSBJjEE3QPlWlq4S9K15exZBXPN38c8vVbRx0fLzUGYpZPjp4u+UbaVby
2VuUN1ft8BCq3KKQ7OQMcjWxT7g257tOu7Lz24U8kT0BJQAtmUwZ3R26RkmRDcwEdMzip2QOFGEF
AqLub7tjrUA7vNL+hDMpEXp5xhRLLfEw/RdW8XYB3Yfn2W7Sa0fwbWvrHy1eZlyEEMpDS8ZV7gsq
z8RTArymS48M9P7z6n6sZe5QmQQYAlDrcFAORV32tuCE7pgg6Dq0qL9IvuHO98zeDLns2QzPxVX4
h+HDCPguqbofYil0SXAVuduDNONjeaI0Popj9pgWut+sYJjTchpK1h5wvSCUssC3lWkgESZPxq81
IRWqBHAsuWNH9AY6/lEY0zSJJr1re8ImmqTjFMbFUKPpBMQAz8/bSyZeoY7T+7EeZPam7Zl2suKo
8i8Y5jG4dVgNjK2CJnHUJvj406kxNIvzr1qayoAEIiBpgVduNPvkU61jKXl5cUO0VDjAIJfu0XzR
k+40ITlmfgYYi+MB+TVYg78NU7zEjPui1DP3RirVQNeruK2FHupTVTmJVsTAGPWSn4/xqV5l/A4x
gKInxnfv0E6LSrSmDBkCQXk1CySG8ysLh1d2w1ZU1FjtmXny1XjfKE9Yy6oF0lGL9QzoHLOIodTP
QhD7JHN+nrlB/x3OSvUDp8tH0pDMtzElrRtqLTN2fJE9Ol42+wK1OxK7Hf/rQGOQjTFbXkhurWqW
rR0kofAroR5B/ha0i6OHqLzFBOGSBagncG/4l+QH9mPlxI+d32bt4iA/eHcqcfzyWcqjnh5w6Ltc
xdc6F4+IbeZC6ITeS1lDZ0nfcM3RnaPGuaO0mvsRLwS6JWHV1bJ1NI0H7zazKTdnL0ROqEZVIm/8
WaVj5zJhs+ziT9dD8NPLnXUKArRC4OrmJL3KL+44pk2obsWea/WRBAz59m1Vr3tajJWKnBYfgfch
XL+/ORx2noujstmFh8KbmgEjrAYkIyAUlLJnqCh8GAO3hrErdnU721jndcxDPjft/vESPw4JXWq1
KSK9EAKVMX9SAHTlKxvE9CeLSxY2aVxYdCK0h9cO4cPdCsbuTy7ztzQnQ0HVDSDhPZqwNc4oLBDI
81nT+wZXmICHyBLj25Eenl8U0KB5uMnYtAXUkZdcAB20hVXRPygDUnTad9kNqqF2izAzgsayYBAP
6xs+yovdlxvZe1noNxHR9je8QqbcFChp06LPQrT8f8mbZ+eBOyNsv66TcQ8fP4hJhZexqkzN1B3Z
krzTZ2kN2fLR3halXM3Nirw/bF+n64Ro0MicehQtuxMiJ9TJ7wM4cp7bggTSCUfZ2153gz8WTPQu
RPfu63VBTeREVN4B0/GoObSQ8kqpQPZWrOzewdOJhHw7UjXCj19QKICyuyZZKBD46hja78cr0Xl9
Wy8qf8cp4M6S9a1EgsLAFk4j0aubkpiVaEAq9LPPnDOt+7vQUFo+JOXx7cegibOUYJUF4q7/FMUZ
gMfVCWIkgYPacsbpO+X9RZiMkZ39m/h/FuBsn7tBlPBS6CYxiG2EnIryhN5mUT1odJQW6nexlcTY
x3rmJWgF8mKNJlwC/xjI4EBkxUDRCjNCb5sGxJymuakOorN6YfIozzALIe3sRpC073s9Olfek09N
pA4mMSNv9r1zRC/5VdWyzRbVn78aEC7gG5CY5Nq7pNiqAUsbI76JrNped1MG6n8E8Tfr4BKzDUAY
aCxkh1OlYzqY/eOuvlYknYo6EKD/i62qFsvgGozJzmCZ594VE3zrLEyJyfNLFJyaKc5+eJVi2u5x
13052x8NoLu1WfYXkcfyYRR8SFL/CxvoCp9ljHNV0h2nYCClJQJ55ySRyYPDpmCCGnMMMfKYmTvv
Se2ZdYz5pKPwkSwosx7ZqXRPCBAEi/XCYGeU/0kual6xl/SGGmQoJEdCkBzNajoXajGEGMGqlc14
1NjE5bYWFaLpFN45DudlC0mOK98frHwKalfbsmi/APFwRGD+Ks4DX8L1ZrBc/JU+qEO9tHpAOgFF
ll3MQHIdG0eL8kCA9ddhWeVeQUR4uHFk3wOyRSgBMpglxyo4/uYZ0M3mLrQTpGYOYphENz07xRTR
TikXYl/4A7WWu0csZDIDNOY9s+hUJfMp66joB20g+YuYMB5KLkKfra2oA06Jo08BnBYaHb51K/Ep
IG6qiMat6IpHA2VXrAWbtFCNcNfSmQFNiLkid0G8WHY7o6Wua9xgdBVUN7dt9rTgUThLfheQfaQg
/1kZPp4G+ZJmmviKiP96UcQ9jgA9wqnWENlmxXwwGGz7mbkus2vezMxIsROYjRaVqVA4IRHuTuYd
3HQ2z7cTmZPwFWnt4pW57cF8KbQ1FzXEJqBGMGAAXe+sPl+ar48JfNd8TDAySFnBVifEFbSGYTJM
08cnU9u0V9a5xclvFyBq3nIEmf9FSz64DKSt28nPtl13edebZEjfUmpOagGI+TptKOzfFNxHqvRZ
Jq9E/+i7BsF8vz4WkeLh+6IBmBrgPrPpADJF6AI4Yc8f3rC9mEep600Cwcgh9ZmTwd5m+jr+ASVG
1pWhcEHg6DxrfRUqJNMUMPcV49b6jMPQ7kD4U/9bbs2LeSXlxevh2XQeaVVuJbWKk+LvrT81h5rP
uFr+VWbuqg9vSLqLxS5wh7JQqs/OrZTQBKStm5botKpCmkKD80JaA9J1oRovAPrYXp5USq72VLQU
C/Sy8fs8EJe8DKSB4jk2UnRdAkoEpOY0lDKKmwpFoFt+rHCdTDXsxSOjNYOIz6m1GKetkzY82JlF
l8RuASL3MV9xVbK7C5o9cJLqEoPeNzFPXmhhqLVVFp1B9Meu9W+lWLUep65XnU/P+7x41IXIuTQ1
uDZlDEo3olf3TI7brV3Gr4fO8kYThvWL2rkH7sPqOHyLo1vIq7QKhOXU7+W0lPlFJEz6yRU4pTqF
21Lr73DOj/qejs+bmP1H0LNQ3CJG6SaaK4eBdK06rZ3XOpajaZLNACnVFR04Zuknzd+jUkFaaZx4
DB6ZnJzOWF1h1aBrzmSNLcYVv+28fF1wr4RZZ68M/vkP71VqH72yj7eDOTKgJ1n22nTpHB6YP8Gb
iCuHXiD/pYCHvFbLLW2Crbcs6jlIpoNWrPbqryH/BAOMYK+Uz3gEmEo9ZVgGUtTvV3kb8FEy3uj/
RBAjK9dJGNiqsLCEjFZ1uZj0VHRpMKf9CgcOg0537wtw9YI16h8etx1vO6DHZMAyKMvRkia/obqO
FNpk6caMyGbse318ITaEBJsHc4z3K9eFdnmdqWdrJ+rWMz1h7+KU4NkGtjem4JZmAcRMwNHZXnS+
6pjfDKXLMoYsK+MiICjVx0VSt2OzmqYYYq+K2V1DpGoJcuKKZrpGvS8LBj17/pRh/l4PIaT8qrr4
6WqOdrTAUkt1bbr6u6lJ9PUlJTYhuXQV9DPXcDGi9sdPeVuchb7kqXJfMgqhVP1cTMo/yyXGdj16
rAxnjnbZHDdbxhAGg89UeLqgmkO2F1xH+GSj1XRpCgYEZBGFSjZvyDwdUtt7SYFGHX6HS1idj3xT
QYgTrNKhwMyvoE27Fo92IcbZbJ/2k22yVr8iyaR+DPw0OQGao9qapjOje4tmdzBbKmWSIsuP8/nV
ZNZ9w5gJz48KZv0wi+AE+C23KxZ17rx8TBRaSXP3XSkFLPAbDOodPR3j/5SZ0gLtSRKW5PqoNJmb
9SnXezRkM3O7sKA6hluZBtfY0QMhfgi77zUKtj9VAhWi9ktVgkMZDJEUCkr5d2o677aU1FbVg1Eh
ng4IErC1Uo1alBss9Vq4ZQDXpfhcxOUy8OPVBUA0O/FIKzTAEI16WPfxnf9rn2Z+VC4KkImjBEVs
GXwMcT9UPAnWxIjTGcK1INNxmTE7FEZZH37+TIn/FKUbHwUqmGGli+FFZvGhN7IQwOVkDnNqyCkj
2ExLZDNdWg/OKjf4x+2bwmCpIN/+Yu4pAJNV0SW3sBuY4c3HWhgAcMPj77jALu8ad8trj42JJ+qP
XcmnBRYpj+tszZ7e85JvIPOb931WKKXo0DeflHJ9E2L7N8tV7imNNfR6Ap5+syyegalqEaNODI3f
isyfUgZyqYh26M73TnCJNYvkNQg1l60A35guUs+NvWTUS1Gl0GhGwGSrGzG+5OM/zn2QmbIex8Tv
kD3IzGS4x/Qj9cqW8BMKvRzQ824NFwZYFe0OYwm65xABJjjBP7AvKSWirxZJj+0YDV/C9cS0u0wj
Io8ggU6RD0sOVmycDv02xVovKB1dPi+ky3bzzjbbwwx7Hm4Dn8Xo+CXctR3NRrwHDQgaQGVB8Ug5
8/LrhXBK1t+cZWcMJTPqq8CK2ey6osH1m49fcmqBLDZJnjL004HnY3vvYIdITTPKVSorfRrWkDi6
YHIw43SqK9ietBNbLYGjQ/Yh92erZZ7d90Uv3dAahlYtr5CC0XU8caOyzWLuadojnPwWYlRie21H
cfNqVMoBjLkzE62V66XJGVHvIPTEczvdBremXa7zL/sVZK2k5WTyS5FoLdt26vMbPpHQvTvq7XR9
0Ki+pKFwIud8Z5youfJuXQofrQa1Kqx9orwx91GLNxTV21Kb3e644R5dYKXxerK+wZYICmB+7hVV
XDztW4CsrHi5UYdQw+qZMq/9EYYIGVZ63tpkS+WEEYVDzs0VILnlSSAJ+iJjwU0f98acaOPsomYT
BFjTzauSb/kZxx8C3Eh/PtNsdOnA5WYV2NfJR15cIy4zCj+PVSSBqIBjpmvztPu5KmduFdlcJ7IT
l8VxraZa3En9pFsfCkOADNaN1isYtZ/Kj+oKsqAbV5gATEYfNHT3MXOP5hnBuIWeIGE5HsQ1nPSk
zkK9mpe+rsl9N1JLMq+JJ+e4ozGGsruccJjvXeFXR9DeeCKGw9OWwiua80dXZJCfi/5GxcVkJq0S
EXQuotpPIURJFvBM7HyICnWGwgOUu+SQh1rrfa7s0N0x4IfIYSfSdPE/3OvqXd0NGuNk8Iw5H4t0
m6HWQ7NrIEWPRSX4k1JPfjvQ+fU/ORnaZLlRnsFItc4qm11z9vuq5GuvWgodo+k62f0mweRovref
lvVaa7RJzFMFxmeGOOICIVnekNfJYDPPg10ozflCnrFZ8xOL4jYlj5s4H5IHAl/AYo6qQUROdTtq
mv5rWKZDfALMfG/g72dXD0sMpFZcAJvRnqBnlnupxUYqNeOCIOaRKnESBE7K0jjCFqIkA30S+wco
adYw3K7tnvyLZ1mEnA/fL5MJKTADneiRHlUSU2tBo8adc9qij3em6btTUuNh1OWpUTrSQQRPnu9G
MZzObAr4SyTv88X0irMtaYFs2kCbw2GYFTXIt9yQdlme0SFULHE97Mj1tSHyubapFFhsUSPSmPo+
EAXYXACXn8MUUaZTVkGBqZWX/Ah6SWXRfNQTJ55DiH0vMtvKAPJM36CO1ZeCqJs1CPi1o8CKZnoO
8nyP3y6YBs4asQHtKpoIAPSCs223Zf1qzZyZ75D1MuxkTXX4Pu96hR1L64w3pVZkZp2mn709D3Wm
uxTaFsGcFY2i/PaosdQ3x3QIu0RjUsKakKYIxna5R29Om5g/ZvUiWFj5Dph/tSx/n0ep2q1o1QAz
Gmp7aTROAE7SyQ9s9qHSa375o4ElVxxUYqM9iz0hwMM+RSZp6kAPfn7OiPUnxVKmfXsg9L2ZlLvf
U1vFJQ0zlMtLt3VzzUHe5bT8qmvHi74jtzss11bxQisoKDeWgZUhhr0+MOluNpn5zEc26hKoYxTa
NkByrBC+yaqNgwk52jydVlsSUSGMimX4X/iksdk5nXPrr0/Kb8MyrQqN/X00+NmzcJJ7nMl1l5iV
VMCyvn0dOcsVNCG/1NktDc+M8JuAoqYskw3YN11vgkFnJNEJdK4z8+PAd54OakPFt2bDks02JvRB
eFlijpB2k7sPaxNxGy78h0na3P+RHTAVst/w1AD2AqkORSXUfxdNxgNWYgffI/4fSwpMejhBqr+R
jofzcp9Pc0RhCUBqThIT0/ON87Uc6AxAdMuthkKOeb2/y9tA9FAtN9IvuGCC49W6nhH0n6IFvC0+
C+PgzjQc8lu1Vk3GtPy9qX614PbXakJApefvrdOswLSFxaqKvPwALSdZ9BQ0fPUGzJljcAOst6zQ
4dAtJz4rMy0d3o/uQ95uR7WH4OAo1DzOotsZJDcF3xCt2iQBNJo/Kq07ypL4fXFtaImBrZAY7up2
EFoYTwbohidoOYXvL9o5zhz+A4BVbfm8jTB2fNx1sDDSC8i/McquJHu/Aj4lfkJEhYMd/qYClXvf
T6JRkSf2vAZDpfWPq734Q9qlqEyTgv9xB1jZEBFhFvYPVLhlmnGfNaF9UTp4e4wzPVFynZMzdRyl
QDPCUpEE0EDj7ikCuqLEQc1Pkh8WlE41dUdg0PjIgspARE7liuRidIYWJOWdvPr6w9wvfyJFfyMR
Jao1WR8E2rVwB4AROnjZJ9xrvS+kN6nC4LvhsY4800bZAXpYRYEl9pUl63xkAGEaiyndJQ5mySkq
yy/QMn/HVvCB4DaFUIteeah4l+QdjpYy5HdcM9kGIeCQfLPFtHgUNgl5qBXZhpHDEtII6wGsGkZh
jDt/jKPdjJBmSTuR+FKWCBE4XrLVj5HpQKFw3pCLTJV0ta5p1JmmL0GwmsU/CLDLYXFmqRJTHmUP
dKXhIfF9INmfRBYL/lHzB9aFPelZ78qIY2Ss7U+eRVr6ViaRY2huLVmCYvkYs64pF7yWgzi4x6VH
PZRoDtN2ApFDn+B1ha4rpeV0I2YWoTfqx5abrGhotrlVCPpj4rycdp5zar1ml8HJvJOe3+PW1+wl
TXlStYAocCI1y1vr1SVqcunEm0rnDmnc77WQqP3yr/e/fnhRiXiVya81n1/LgmDcy1vXKDei8HVK
Eoh51Zzr3qhVi2bXZhuOICWmcw0BiBrQStHUK7BNQf+B6MPlCtlg1pFfGtIFU3lGUQw8nef0tz9M
NNCdpz5kzzlj3KaOR7Ip8WzleBgfHoj0WIsX6XE/OUCsAz7qyAaC4tz14hvoB5JPgkBKs9vuzgAO
UXfTN9FDiZJhChlRqUEwNAW3zpzsUZChynjtZlVOUWdYPn7/EmwvOfWdfhmGL/IwK3JnlioZwnG8
suUKjlSEXV6LudFqbJjgKYHZzSfQMS2BFIIc460KlpDRetMi7Ir82QIWwHQAuSqs5S6x2Z2dEoEX
oEE+3KLITSTiqYvswPuMcGOtbkJGywyssZroQ/+r7qlDHZxyrL+XT+SHynzRDlM+O/0c+NyIq8bB
lLj8ifpkRArUQS47cXIAg5T4voMdkB+eq4E2tMkPm6EdlIHDF+/hExVMpUsa1S5+5lysIBRG8sH6
zvjmN4jjgANNEz9poXtJiEZUrkWFqvJ5/UuHyDkWwtGhZ2rndeo+rOSqUm5HUtwPXSi52cuOSUr2
n540OSeM4ULWTCXgJyopqUlc6pilce8GlU4q3lDz5+F1aFmPpZYWRXryjofGwV4EeH+QTUAeENVf
NEUeCHoYxWNThBCpGWmrNa9eOnPt/bPSNRBjb4VNInAvBXp5o/+BUb3T7f5PO8O4TdGGmMxkeT+w
+hheZw7GyAnbVA+sYkPBLm+w3YziXWqNQq9fC8shBD4BfyF8apC/ysoOlNY0C1eYibl8ll+paM76
qRlg4Veu6cKiI0AA4YXUgjgDmEEPDIYgPvYI0Cz4EEZz4m3tU0NPeOWizd1BUUu0bCwKZdJYc07/
DjfXJ2TtLAjV4E3EeWYYxzWZvZSypHZffT+eJZsOEPcjwaXkmdjy5dXDf8kSRUxd7RJvVVidqSvl
8aB0qx/jjVgWXoVu+rcs5t4qXh34MCnPtGOLFksjoTTF/bPGnLJo2V5Nr09JW4N/YAF/X7GIULvh
TdmD2t1sB6ZNKXj3/AbH0VdU/Hw0Ehpf5rsEFoikwpC7ObnsTLeDV0Kb4WXzrKeXDdxM21VIzdla
BwsD20my3k5hKoIYuJyBX3SmMzf2TGsegFClKcs2CY34sOy5utbXEAXxKIuy1OXbk3oLFW7I0xAv
D59JEXu4yPPk3Yd562h0I/BoBbo1DioTX6hxlB2OUO8lWuf2Scp0GonyEKnc1R47dPBzalb/McgZ
DyJNmzy2KEsvgEuFd+lvQjZkwiU7cmIR4BtLbjXmkBj3ERL2hCYTMJRhOmDeWnlDw4ChIZYLEMtC
PhH0MF/IGEAmcAxxW+soC0IdgZ5MfXRZp0NwFDiO3O4iGFHfOzliHSz/qLsB4sPRXyk5ptrqVzVY
cv1dGyd9Iv07uR6oel9pOlX4UTGkrQ30iOt4hY62Rc+1p+YmqDzRlnJ4+W4Qq1exmcjgF/77ril+
odGcwlEkQvT7xIL1n/SvCOjGlwTq3aVl+4zlGtQJ1i49aEC5FUJnfudYcMzU828S0gD1cECP5MFi
Y781envZehgazvQlj0s81OOdnKqdX1veDc+RwGJHccWSMWjp6IXxHxqzqYcrJirVtfEM5WF+tX3o
7G26MIlSJtcXwUCssWjE8jDdxy0wEnn9jdJnBCYFkarOP6DNq8EehW7aiRBMiuy1uoK7IG3tH78b
lZvHEcnD1tz1WP0TjcxHvfas/wyxARqJbuEvunGQ/Q2wOQqiDRH/k8vtVlWGIRP+XIFKm7lAFolY
Z83Mucc75QPVJIW+Ii3hS2gB7xm3/2OdbVxXN8qYERh9c93z1KG7M7bj9Sw9d0Bkb2tQIc/pdGdC
KSg/yJL7ICvHMr9Hg7oGm+5STeIRTjWCV0lIbpU3ooF/Ie2aLcXgaTkxN+HOLujdw9eXq1p0BRY7
OFQLol1WjFy4mYzsyvCBC/JE0P3iDKxejJBcnuhm26GIcne7mAHjZzeqIjTElcZ5mU2dftZyXGgO
0hYf/vQivOoGvzji2ml+LPbCk6MPVjqJfxG4VaPlxc+ga4O3EODDWHqcUVoF7dfVH/2bCnC8gCOZ
qpYK9ZLGKI6UNtwfSNKVML5D5VfBcHszp+ijZpxvV6y05uxKITRb1ACK81RIfnMcT1DFE8HY7qBm
8gYzeDwXDhgvIEh5WSW1GTIZ4uePEinDVSNlU3Ag/196tHZR8P4H7/IB3CokTqPpigR6d5X04Zsf
5pxmsrUpCWofiriSNes5WMgVZ8Nc4bVRfXQYz4b+OVuIrcQKiWRdHPzgcNJNk47xcUaSpPxBHnyQ
9nOBSFi91ihgnMiL+WFC++VOGXlKiTc7kKyCepDCOcmXxsT2fY4nYpkzGP4OqAJh9uE++U0mdLFh
94oxp20207WNACLm1qxOKpfuiwx5GUe6WKoQzRoKh24Mnge5F+z8wGv0Hz3lX8RZeRpM5OKysFYL
BgJAww2HrTVNqbzsgty+8nIBU2AZ4WpvmcHVmQXEaQHzKqWe09SFuuOcmumbLOIhBk/8A5VyEXe9
R7q9ScMMRsrrzMJbTpUJfyp2PEadbNUIn6oY82Qqk82Show8mN9Iy40fDPVLCGdy4znNq3kC/eKM
Oy4tBDXXTR1KJHNh5XxtXQGWeDqbNPN06oRo0eP1DieX0g67HiXxopJXrErTj3S9emnioiHdcvuv
Xyz6H0NJcwLb5/rqtblzy75RMWUwgLltGlD2hstQt50tiau7UIATgMoJ7o27je0xW4P+I28YD2gG
Z+20xYT97cfZ7lvWbIQwmDYck8YCsVfmZh0YO77jh+jeSwbiSKWDgfoejmlt40Feu+C1daMSnH82
b3tDTLiAZU6+1Bu7PkGSBo0WagNV6oDsvSnEUpU3wJFUOC0P2alclbasXKVQoEWIg7Fwh8eeS2By
Wxk/z4ZEzuKpzjZ/rMus91UOz0maGTXuVYmVxQe1z8fDX0hIKAO0+I7kijoRj41YxkeEmH9CpYwu
IHFOGDYtbnKq95XpWWYip8LEy8gNqNtNgia5XprfrL5sNdcaIiyZiXwZ9f4X4U6oyjcfU8Q/hHy5
hB6W0MuQ79E9WKQ1hF5jsCEDD07HPWhrAHDxwvDvJr8g28Vq+n7Jxb5DalcSmQFiYwswZLGpye3J
Dtr/aVBE0i8lW14RYgQxJ8ZWgDsRdPgGIVGHPLYcd4m1P/Hb0QQVu9qHCzaOhrARWzewp+3aFHp7
4JlWCNn0Lakt2gj+ixBqwlEKpJYtE8D781fJKdmz2PHyO4ZOEMqBW6c81YKvCUK2eK5bLx330BXe
gS5mIp37nSqDbmFyzk2NbHTqSmgQIdUWToUycaui7rZ+e/b6EAdiTfmB5nRgGmCcAuT4UvXMPc+R
jIgPXKlbqxntsdY4FE8Tcz4ug9yajrwkinhqWdsH+aKKV1lmLAoXQB2AGZIQo+K+Tp8SGuU0El5N
vpjs9OwjNl3CK/5R3hdQKipN7NdR0F6i04oACfwxfERhcs9EzUpp1oDB44UHjXsMEf00EMYTYdOC
nJaVa9qjH6zvejVwVZOcl80EBuYbiuwBpVA8lu6OEPQRWRBZEwC36pwszho9ZMOed6cGGhJJPz/j
THUeT70wLWzsQ/yIfLXvVuTopnAEGhKn4+RrCh3WVDPRwsjubD7qQ0C8vPmx/cqrYQogqpfqkOt/
Mhja8T0PdrUso6MAR1K2CS8iaCapxntJwd/o2bb5HhFHZy1DQbwTtmkhM+0jiYLaFCIwee1bIcDi
KhTdh/rYVMNrxudvopcRxsNxD9Vn/KQJHwtEOEbx6d1B+KcWii/tZ1wsd6Q79bKfUEwxaNNxALCM
5Dx8Ar3w5+Ayx+5JiG/qM+MUnLB4ata0rNyR2l5f4PGOssJpH9+elgQQLQd0ovrUQPV48KMyN878
7VV1yOYbjMZhOYmIACFJzft3FPbD4GdGQF3rCopLGewnuYbP0FMtkwTCekQylB9sgxilUtLNb4gL
YI5Jbg3cg5XTH6UZYgSFU4OTmK1L0kYQpEOdd4ahqdYyMuTsRt9Ncx5u7/6QRzUz98MrBUz82ha/
xhgi/nWME6dtk51j+y3ofsW6IeLCko8CqhSV6uRtWIy+ALTpyaofmYOIVUv58UQn9B5CUspzpNDD
ghncVQFugJtVrldOB1Afks6u707Pf+MlaSQ/u6u5JHetlyLnMMC5t9vC/vtPoBK7YwFIZ4+6QJlV
iK4p2H8W6GaA+aJZEyCCVhyp60jjBzF3qqpZkbqrbeeaKrJFxCMZgF3DsliIj0d+4+IqtFlFi1hC
WvWHp0bPOa2u1blP4N2HLmZY/ScOCZWIwYgWagypfRPuxc1RSvYHIxQ84FfFW2WybfXiHtdjGIGB
hgaqVUhuRjOUTYP9sx1d3ZEhL4jKyT/XAaZbFnH6XL+ten0F2cs31E1l/oKqDXocsvV143MgnOsx
yJfYB8nCmNWDq29xGLFtQU9F0A6R1x/Mio5W5iyLoi+bXrlWu1mZZdc2g4kHqb3oX7HkG992Pman
uCJU+5LanqkyWjTmxR4BQNDhMio6EzBcfoHCd41zypss/BkHTEQK7Ep9NmBch0ASz0/JbRoLfDFB
SjHtDkw2HLrThA4jI93LGtqEVHXqFwIHiSYBfNfenl2Fubs70p8zhCSDKhAWHIzHvke9L4m3Kn8w
2x9sokRde8Ddj2gXcTEAZVlhe/YAS809IKEylAJkYw7c2Tj5oL86KXcamSGrO+37H3G0jFj88coh
DEgPcNEFrIEtanolguQe/yK8ghJpX43p3Knxqtq1Gh6LD3jeDqRZfOyER5heyFSD1hHg3AcvM09u
LkoeXdj7JD2gM83x8rDVogBbZXvN53+ak8xoENrbl85cvAp9GI2FF5swDC/G3ueBC7uMz1gUwPxd
BbpL7WyEAxCdYq/wX15gBkTxfBvJT8++XWr0zK9GnMxSft6VhESRQB6cDmFEYUnGEi/Kc5+K86tK
ME0waFJu3yBSef4rXtysUNg2Xxcm1K19P1P3dKunJzO+7yTS/eUz5wUzyjsi+XUseJLQQfLI5VhJ
GUMTJxFYlLUWVuszdSphPJBFbHmNeR0WM0zJ8q0RBJSgXZg8BgxA8iZPyqFgnHyzMztUFoCtGekh
ezz9oSzyDonT6pxVW0RpPKOhrm1oFOWQlZpuVRxAw8UPMcnh6X4JfbOjtS7pheqozTWxjM9K1UvC
7QzRE+Q24ElM190HKh7H2bkE+mEplqYzR1wN3yvZvu/JmxoduI0BWWCnhn5Ibvb+pYT4ZNb9ANFs
Vvdg5FmCu2sLy0nLnQdQSevxlvFx12M8s/SFwoawc6X5hvsrFPnknwnRVIBtla1nqh0mArtWdhIG
+2/dUvSiAto1Iik28/pPHiPrvp2R+xmrlU2F01V+Ir9lxgS8LJ3aCSFTjJtkKxyjccDVeRRY+8Ln
VdcmkKn/fmGAzxEhLo5cE3eXma2kwP5Fqo8fPynjWrcVLuGIME/SxEQ8Yag3VBcdTEk3/GuYcLG9
/f1tfyA/J4ktW8tG4+xUBgktCAd8s0P5RtgplYftPs+rML7N9mwoW6RKAah1ii6nvyaGEtDqPt4a
z6cVdI9+IJIup7fF0K8Dwb0IgDsIQSSHBbbiI7fFC+0Z2FOoom4kismJNcyNK3kbEet1hAUhBcus
Qq5ZwtBhMZnc7/9lIRarjpEZSisANynpwZ6R6Ba6RgayTlDiC7JThm3UMEv7LzpZ2t0zEvNMYpmE
3bs4I5rCafspRQrQH74rY8x9d4u2qaczFA2S3C5gKqxDCXnkkhX1jIkzqP9+svGic7+EMpaiuSjt
CEsjzGzXO0y9pUyWTtBB1kypYD+pJgprgBLyrHfP+vZlSpRvnf98QwWI0rSzrV/53fQvjewXWoXr
XwibH8n7FkOeuonukMupB+qhEIUaHeuL2t/FvIEjs8Rzar21Yi0Ll7K4m50XjU3lsVeNZTVv+voB
KzAJKmFnUBIAWOv0MiqGfsFWxIZ4QR9dmk5hlo8HqJLX6mUveqApTzMsfblk7PipO0DtmQzeLWy2
XNXQwB2zKKtK1VUh7gSbekCvNBfST+v2Cg32mKeAfP3N8iSXPYotlBGKoq08YJuzOCJP1xeJ+EBj
z7zoeMA0oXxZCsAuWyLd0DCzRueUhNDXU7nB2mYqy6skz8sTyqa2ypWqxzRAEHvjkuPsR2XeZ5cC
9kou6aWrebJPawqL6eIeSa1Qs38xfb9J1+WzcwxXS3FM93OBW7K6+BLsYsb+uoyLBiYr60z4FDWC
Xuk2ooENGg8etD+FVZmnFHHtY5THB3yQfLXeiaQ9MfLg1/awBvD2lPP/heCDTHodbnnr0LshfPfS
7B+GWd9MJtf0OviyHC/zptZqLInbpJPjCyeb1s1D4cUK3WCm24hwTbY16N2yTf5yL1epMItfCxt/
OJwi6uke+EieaXJkw/dgQ3eYxKUrB7/O2eu0M3lCnBBDTfH3g1oBKyYooUW+KmughMSBGgnFxNV8
3Z7TafrPth+DjqAUzwOkBesWGlk66p/THp4uu0UHahoEAagKzhsjNhCcgKkDAZ5ai2cHwCTwcPaq
yzJva1YSg1F7g729mHdWNWdveS0YgUMdkEjWe/B9RgaMr6GBJiDyZu28cGvVJTrTq0/0WUbtOMxH
vXmgceHcTZP5VNGoMtMYIP6iAWgmN0MUBi0xWY8ExbA16ZnDnicKOLxnR5VhiMxgwkbMMYM6YlS8
8If1fs2NPYkaCfx7kNJGE2i+SRPkGEoD7mOAKB82FnDdha8yKUu6t7hMq5RqUw4QF5GfbmXUp0i4
6wfR2VmsWjWNi9eYtbVFJ6VN29CmY2zPnRbLfiHO0Cb+8QlLt6As+XNtm5iNtIdkYVQI55siYt4Y
OZNrSlEVhyd0b6SOoF3Tih3QWekhVSuOXvZRQXC2L1X4gOVpUwM/MKfrna6NyfpxivgtZ2HnPejl
JhcjkGCbMQyqbOoRwUpl4ACoZB5t5xMp2KKicAroTPQZWCoSalYseVcIvUG7rf4jbo2UzYBxcl2U
RtccqE4vP+Q8fkCiutnESKnBEO+rPluRuoOcLm/bLnn+zabU7Fa4Z0GrJncJ99ElOYNXEdB6mc3/
tw1K/lxj64wlk6qpzo1S9bgO+50589qCuC+UpZhCCnHg+Z3ZIpBstS9u86FOUlJ8OWZKZyDO4B9q
HYdHOPXm3Fq3P/S/Y1WbsbOf6rW9un8IW9Rl9h4k+E+MtFdOt42NAhLbyV5m6aVAr03YeRKtJw2h
O1VGXZ0aNyJl+KHkoznTSmMHiDTuWKK5TLsKABbecjjoqhKVbwb1U+9cPtott5uYIxJx1I8G/djU
/Vaeb3TTb/SDJrU368NLMgxmvP76U7swhaDGKhGoinljJme/7QhRt1ByykiUn5Qbkv1zKInE0ja/
tE9mmDEZ8neeBh6Pal//NCAJOA3uzmGA8hgIp7siK84JwblsUfeesO5f01Pd8AsTaaLrm/AQtn9u
O441415spdeJrvA8gi/EaUaNg4dgUGRGJYx5c5wP02E4UlkOGcLNWcL3YaE5hSo87Un8jfBjU700
0wiqiusi1C9YzZSNCOQJxxmMjjkIgEDyy+SyTm4zBXf1ExLSkBrTg7SgpxLh/hIBXH0tEZ7eGA24
q0WDfgBs8P8hayhsZliC5j5LaJklNKphUsOfn5PpQIhsDelVfK1dO6MZ1CmxDocxQ0yOCYj25+VK
qgEvnk0/GEZNDYDImjzadi/YEIlth66xrBuRZSfm7UHlVjpJBRt2XFoaaiMQwiOWWij5GVLN00ul
UTJWCbiRN2PdyPA1npkuxAz/sMyGMKSrXWq5BGC6HNh17jfvINEPYC6F7ezI3YtsIXz3iqUBklEk
Nv9G4CsvL0/aWfA8i9Vl7fwM9qwdty+ovXk2kMZ4ETEK1WO24/kffeTFa07d94RddNc6a1oQ6mXQ
DNQkm1+cSUrH1ig4sTIEy810HHTcX2wiDtaLM/ac85uH4FUcgDYEx/X4bFzH3LqFsCdmfMP+muJg
DCAdezknAa2IoHCBz0tulztBve6Y5pT5r1EUHEY1+eo+SfLDZxmC9viYIXcesrbE5QAwAAoYxHMU
ojKLy+0OgDHoo/+TSng1OLLrsrsdABGCHNFBLYaaCJR7HVuvy3xHqQxdQItAkB0jXpMtCS+tL1Qj
xeM4fvFTDhU2qaNaOYTx5xPvbPqsBRkPMLFhHykQnmyqr5j8cWaa2JrPc/w0QXBYSQot0tiBXunH
1j9K92ime8TR7KRyJN6Gp2S8BmHC/91DG34Krzo8TbkH4Lkuh4YZp2x3rgHluTgP4Z80RYv5ivga
KFVurwXw4n7fnqISpg2/DdY07Wmje3/mq+dlQ68pPiobnOt26OKsEUzw2FWM3ZLNbDQfJ+H9l2dJ
zbqlkahM6acaJXEF3PcoHtKDrDnmq7yH1GrjPK5CLta7SqFRRyrD0dPdKpDkOUPAVnkENZuwkP1+
/31E9Fno4cTcjWsyqBLWGZc2MOEdlVBk+sQqHhhP0qExJD2kyGHthNJEqSMvhBFEB1c9amBqf0ec
Hk8uMroW8Obp2wFc5RgSqe0kC0CH0cZIHTJK3hgL3u26+d+yYuvFNOGD9TizwyP34f9cEZq4u2wy
gzXpNRsh7Zxn4msnw4AVU2JdTnoP64y4RHXmV5XT2H6yqAig8tbRdF02Abz/x0mlUQLxxhqQ36Xv
a7zBLCkh4cqIWw9/Z3icUHzYdaQM1ruFfmuMc8uiM5+vrbzDhxnSo8duftgBs4zoJzAHIttwAvk9
Bly06p/neMRnWcxb1xzowrAedrYotJnUaa++Xev9IZpZSqdPGn3QEykqorNEEwOyGCEsDNnPfuwQ
l9N/7F7xDdZ+Gt7/UpOMve0TYoI/sr8Tu84O60Tz4dRhY0dVrCC1q3hRVgzFKchXdwLrg4A1XoGh
7NfUmkKqze6+kdBSyxh8zHr1mxLCLfk0L/BMd8zELA6NOOgZ6Vf4pCE4HKEi6TXlNznUy4TcisVn
pPswMXPySNBa7V5wRgBhfsLPXFTj9df7sLTzX2Nm1W6REjn13YhChbDxhTees4g9sAzM47qxfzQQ
+LCfAG2mb5JZg1kTpYMO3MQSKn9kpBI/Gqj1/as/Pq0cBxZbypGGgnfG0LyFsatqktx1wHAa5nuO
jLwubhZnv/lRC6LxFhde/oB2OeIBFw3cvLgGAX8mKzXLlPgmdbfmT++6m5UyIjgjkHcO75FGOE6+
UbkSQ7NR0pUdrpjRy37wDCd9iSgMovIwEPHUpkRiIzdM/eofYapYAHU9Vsn3xhlqJdgEzjs+AwPI
M2pyJw4wiEwrpboJmXgkUCgP5CTjzhVBchoBtdYxPAUVDcLajxT8TysdJxj0paLVAzN3LobRXXV4
I9Q3pQqsNs1jHhexHstoZeI4MzvHR7o/YR8K43tYCJ4fHuV7/Y7mDa+t0s4vFrp9UruVA2Szn1gB
Tr+VkK3AP4e1DsY5LeLQWKYLg6vfZWARGxrV+K0EjROTlGXfahgq3Be+MnJv66QYZTVbwCs/nooD
mgt5l3DVxK2v801KCqj4lL8sQ3ByDaRq0wenHtQXIG2qLlx/2Ukb3zFC9CAitHVH8J2eeTCNvdEK
4PgA5ppI2NETpkr2e0u3cYyCJAtn2IqIRTCMNJ73n0WnEnCnYu9swukCc1u5ezuc3h5CukoGwVno
7oPKvc2QnTXJaeRXblBaeyUfytdHDTHOi32EK/G9Z6nKc55OIkmunZVUjpQ1fOknnDBxKnnHb5ZA
HsPqccB2rCCLp8s0Ojzyv0XLn7/uZZezeRroV885il5poOc1XxrnmZAX8stmJU2LKtoBIiezj914
yo0b4WjZv6Zn6qB61AUX8FE58bW7kHrEx53W6AujQ/RssZenVM75fwWJZXS3h9B7TB2NiSM7hooT
3N31pjAZfmVEA0+5HBiXmtXp00/EA8SsPz3NfJo5w8FIqCNIccwLyDfWj93CFW+yZULnYn1CdbP4
juFTnAQkFHVoWQ4fdcpiESd2ahpQzBzYZ4gGxeOm9uhwF0Gs6k3rc/eNxr7SfKekRJaJEiyhBabq
EQFbFZbaRJwA4dlthTI2/G73Em3jxKR7mrSnlOdAVAeWFvnuJ+f4Bji/FKau+DMaDm2pQ+FrG/8E
Ouh4W+GQV+UB3WmnZ2js7TgBA7CUfJPs07kSdPJoroFjSk6oit9Abn9jBl26M9klhDeNF1FXrLJA
VFsyjUwPyFunXipMez4kTGgLdpdDXKAvDrdZto4stG7BwBUCXutHosJi46NhmUexQdhEAcu5/pIW
caJ0p2VexyXiCGifFDbSufF5cff4cF2bHmdV81gIeKQjWE64ezVBvrDB4XtXugPLZSgHG4uzunFe
PqaKD8vLLb//k3BoeDvSe+v/p+k5qrzYS5Rspr0oW7mEfrmeAW+UTdSPs6wA0g8S0AIjhe6GPEyd
DCINZlNMUCZ0Rwwqc2Lk0s2cvm0YnMQqGSCEr14aq1a9CerUy2//B0wMeyXarCouuX5L0UnTbOWt
rOOJVQYnMfLHiRa2q4pyYV4RieU9UDhLwKXSVMS8LDTDWvI9IB/4ghVfXq7GcmsKeoi1NyPW3sCw
2uP3Avv3w6Tv3v5LTdLBNSU1LlG2k7POIWQ3VOmP5rtJdFKtrPAuioufpxA4/GXL+ZPR4jN1dCr0
4IPNeRVsV2bb5T60Qt9AWpXvzv/6X9191nAO+BbEh0+JBFbs7MUtnL49Ll4k0oIyCnr0zcKinMQs
/BAAytdoBWoNuSeukLOjHuxhAjPGVPLRs2J7siUvKBi+pnpRbQ+aVP1uKhhgspVmCkYYdKRRjVs4
Cnem0xpe7iS3pCh6FlgEc32/TnMUufLgsLyd8Nsq5VQ9M2hNCztY1F4Ug+UjrQhq/ZWInHT18KL+
x6YSfdFd2pRbuLti1/7sCBPyYFrhZhczLu3wb4fpw6A5HAieN5hD4k4+gFyDdaebzdsjygBki/pP
XgIVOrkK7LyOZJqyoE8fS377U1kirAsMhbABEdZt8V4pacKK0qyFxiD0nM6FKlFthXs39EzzjZMp
h/ol3UfE24oAtgoIMm225gJq9YhJL2GLyiAqQqRrmU2dn8GUwcQXQhazoE6EyH+QTB/9eyVDKxTN
YGuisM9SaiLoNmLq7vf6Z1RlwbB9D95AoUBJ9hB3/lK++zs11E1Zc3tA7817E5kuKOJRbJdZkknj
15xpyIi12n4kHYb42Ca44tBO+lJ6eedN1K/yGO80nrOJq0Do7PwxLV6L0cum0CxAYdWggShpj2ts
rNnaScpEJYzWJ08mcZVB/UoQRD//nGXU1rFUrmWETVe+KsvtoqGtxOzyADxBFmmOx1NmXWjK8P/S
752PT8k28l36Bf3kA8kJ453kYajucZKdPTrMgLXzmMOG7/veXHjuQr9L5XFkdfoIigUTsog9bL4j
rKdTZ+6SlCx7uqVEZ4bQdO+NKbqRlZPiFXnGHek6aQ2e0KoyB1QFYhuNUw8nwWwcMqBFaCLq5lro
3xauIWM/o4L7CV7mR0WtleQShV18RhOkU+olUeW56cM0ggUJFUVg7XMF4LG5DMu1rL2vZht7MxpV
ju7JPeTJ2wulX2HqlGrru55oHKr99Q2w7vPaPG8Kk/mpVwEw6omaE9+Cbn/a+xnuuD3F7WBjVvYx
rWq2HFcN9LrwnPErmyyzNX5K5Af8c5YvNQ4PsreRLP0j3zVcjTLs58583dx9a1K9XjwyncrJ4w5E
TOa2Yz82UmSvfrP5rolYhV1E+SDRz88UnB8cUabDucaeRG9PO9O7kuFQEgBb8KNtwnN90weIN8c7
6wS8Jqsr+diC9AdZXz6NyW/ZuVlcB3CrSs+jpItnynYGPeQMjjeJaAcI9PBi3k5E6lEU1kZZsiFD
tWLza4K5kOd/VFdch8q3s/IIfUtJYT4L26GG7nSdpPpJKDnD2axUWWXKgX9Hgq7x+5qLOFBvTZuA
JqnWKNB9CqGbsx5OnVc13A/yNkCLWF3CUWH7cb34UAQiSqKKPcIZ2YkBs+rNhJPXnN1woKgrpa7m
J4WTD630TJ213WfM3gcW2F+jwzAWhFftYti0sEci3i+OYVQDSEb66J4kQsxaTiDVL4rjqfrrdEtv
JbKtz2EWTZbvXi/IKak4YS79Mxdi0StZUPQOGiGwGm0gxJ1UtilLnd5CcyXvyAI5glra+mTHb8Ye
Yv+EacJD8yg0NhQ2rj9W8D5leUMmgKlov/QXu1vu6Zl0jNXernytdU4U1MndCzb1a7l5GxtCws5b
ZwJ+Xuua4Vh2j5VomRDHZ8C52JS9aARhfpe+bf8HEK18vZq1MgkY9U/XuNO1XqBwvKTP/B8GXbN7
OxpkcbdmADCsYtZmgRrebKr2o8Ksyl6ZJxSwPPEudNclH1R2gl8YcLs9p1TwK4uEY60CZOYIB6KB
I2ktwX06BEMEghz3NZpsMbNoZJnlcAZi08VyoPhlXLu3xrDKYQZhRH95wXohsRC/6+Zs7DMnaUvy
AWSMNc7loHWSX2QffANX+qBMMnT6bCqniXxC6mZpSFMJk62fFXowHTWlE7CVpAkNG/IenJ15LV1/
0m2VkQMnrpppHv68E4xUzrkT1y+ds6XIGrSFUsY2uQaebnTQ7RDdcqYf/iVS1ZQgtJLzQbhNoUW5
gaX3QsXcQN/yBBc654E3t2zUw2jovUCESHEsQ9rDWqWVb76G4PlNEDS6bukI9eD+AheIcJhMthzF
srgV3RvROygFK4S5dw90CDT8vyayjdZR9jdudLaX3E5xiXdCjk3/9JIJD2RMBEKsedDNecdYDHjp
Nszo/pygCH3hDjqwIHJ7v3xeD8DlvUoMaSl+iLz53/kowopwkl6QCpz1sMm9zOMmKK6mQJwboaLS
AdmrtwUIXld8RBp6Dm/8orlBw4e3Ctztutq8uxwPQty8PPWpp9fExC78yshEfN+xpR64xP6T4TF9
/aegEMmh2fxH8zHctxiuyGbDjbjJm7EPBaA3y7+2UfCD+pfwopDNBZLC4JD2oUgOIIJ/AjAu9eeW
Hq1yi8DCoQM9PgVY13hnI7OdKdXCEUABbXhcM3dr5Fi4Uy1R/1+22RDnDnLOGiMBrpR6tfeEiUbW
PwJ0iWUnqUFzEUpy4myltCXAwetZHk+Y8LbMSOtKUDHLE/owHuHiUd7Grwqnd0HEgkvaGX1ihrwF
s23dJd9Oquk6wESAwuw6tCZ25ES7swq+AyuK1yQoOotuR2Q1VetjHiBbQmrFOLMGb6SBZfEG4c99
ti7QgVzaaF7M6Xh6QRBq1Upv7p9ThqXW7OirpVQo1HZdrv2drXfJkl/9x9H08YknW0ELJ3jZ8mBw
NAffgX00xgWGmTxgF/AkAbENz4PQkzMOgp4lIeWTAO2GfSNd6eFuk9uPW0FXBTnHv4x2Nz3jx4AQ
MwUesM2kMGY8S33yJmshF2DscU+aM/9FFVpH8+Bxq2e2R+wyG0J1gcrK1s84j0Quh3QPmwk1ZksU
hvuyRBY4FRRIypPX6UdhRNT9OcY+sKdBZil2/vOhuj2J/eOH/pOokkppmVivacDt1Psx+sfBMCb8
s+23676nRcIiFcVe+sDNQQXnYpflabI9amDQIAopoQUEwCkKpMFePqxDF6Kipen80ZS8hoxToP0c
p+LLPum5iYSLwYlKBdDQF52F+odWYefHjmE5Ngy9iS5aimvqPyqZT3iLIBqU7z9O8l/EWpbUc0Ru
d5sHrPfcn0qr76LIp9EmqttwXDdMEAtmnSt/si/4u0RZlWM2en1GQYao95BbfliD0r48YFibYm3c
R/uJbPBj7i6wGYu1CcGMc7sg4HDlxaR1M79KOHxF7YpPIf9Gi/ABVPpoAEPwAGga51YWk3jZiPl/
XLcu/z2qFbkicedIAiJg06FZNjsSpUnWcDLg+KxjRxBqjhVFo1kDywozs4c2MvVlXbApfHK+H+5k
2/xg1YSGKswa1sDFKSAj8VIUUzbVHkpnpIeHdXoQ60qqMJkM31P4Wq02yWRzkMiwR2pDL8hfYLkQ
+sovfXcneGnNnSkhZTHk/zVTla3ObrpDwPoadGHuwnWHrrjvdgsxzMCqgiZqWqz3/W46C+shvowk
nD+Fq/arv7VnWavMaVOifpfRJDzsvDX8y0D7GgJpE+Lu2ENFhrHtbJkVyOI7TacYBpb91KhQsMO2
txJpFtnsrO4sE8M99ihz+D8J2ZV+OrinBMhEBMxxJEtp3Uvtb4PtjAcpF8w23ufl+e9eLV5ZiR5G
9NqZ23RWQqfXhtczvh3iwAMZ5b610TIzvEYbMpomo5lTWidCPhTU9lONutkHSlbKJXJhRn0mTKof
JOoSPU8JOAwrKVRZ8Cg9yZphzjBS2MbMcxpOnp5BDdSFHRZTjigIPENpN2E+awvQ0NPoQks91BI2
t0z/a5KlQ59LbpKlmWhreCskK9VohWVnsPSQd8flVdYBgjag/TYipBFcMtCCKitshBVHGzVvuH1B
JGwIdUkz3GEIvBB/RFlHTOpdf08x13sn+HHTZT8OZSoLVP3Da5R88PzjaIVEVSwXtgUevfEH0+BO
eOCbQOYYheNvLCrx7qyaBzhuKSBJFLs3KE5FdJNeWFjW//z7cceUlJpKi55bsZtdU1GPz4MvWg+O
JxY+zQiESE5liD7N6qtG3ccEYGe7vtnjNrYTQ5KYMp80XxiUAjLMKBT3tGhz69/Xo7UMiDAeGK5C
Cn/F75CLat1bX9MWABrpBFeXs95uVq43yuu7yxCKohq7c56Y4jSwSDknoULP6Uz8JYOCLctWeiO3
Q9SGxOUOwSEpe7ZWTbmBb1zcTNGgSo4bkhQJPvPYzbS25rRkVS1RgbR9HIX8k9TZ1t5qjEjmpOlC
b6zlHAyvyzTtnuF5IcbwTEw2CxOm/O0q6edLdG/p4TA3ZI6gZkbae8zatboWnVyx3uPdgFB0A5+S
Iofhj1ir7+OlZVmYI/xEavZgm20NNd7/OUGlHOmkv8go8EzJyz6GB7vnTEAoKsQ60SAMiGRXJxDI
5eoGMvI3BrTELgUZDMqqQgh3BQsLf/uXXCrQ7Hcd5IZwZoxHewR7JFa7RNbA5dbt3ZHRvfKESScG
Gw/o0G1P/eTw/bl3/F88Fg+ukBG3MbgJFoCesd4aUbKvmXyP4JSDFg9rXv5HlchwPwoJKLPHyBLg
ai9Y9Nqf1reK4pKnQ5KbA8rGJ4GD1Ac2/UyK2Ejc1IxdhcL2UI/GQesIGr5OhfPIksVTvd0cDjYD
BaUbpLahGaaAZMcA3/OD+KMqUfW0PwPbUq+jeSejBvy3ZnGcqTDcgadyK5NJ6JW5dMi2prZJpMAc
HeeKdLCxKqfyRjJrfWcpBjJrNcW/8mJYyfmG+Oe3i9V6zDPtuU/s4EHZmAv/x98VB/nYRpmbZQDl
QBnExXnO81i6y8z4RNpn6s7R46vhrkN3MBGReC+F+U1OSgF+qg7Y0+NWXxHaka7uiAq3T0xtFG8o
fEv1QHKBrfB9EajoiVideWk0evWMUdZo1/AEGLknyFNRTzIfKvm/pq5n6xhRaj9rsp3is385r4Sc
x6UlJGuoF+H/7F5etq10RLr8x0tR0MqzTOrUlVZeQYThqEdl2xown4Y2eFwg0MrRrwwKM3bOOucx
KIGwwxKEyzs9fL+F5aCaWcNRmCsCdkTxedWvWzZYIjklQOd/T5NYRJFCctE4YvcljySNOOHOd1nn
7zMkn5B3MobFRUysrzCIPyHnCsLvY9AkCuw1OzDnqoaPi9QP2F7u44LW5DhE4zE/vremsgCDzxLB
vGzRKgTvkXYBat7o0lJzTE/tIU6tkVcSBeQe8VZcag+u4W9Om0a8Rm9UdUrPuV8Nto6yj1eAnZVX
sMKFgkoeqX+CjKcHoPCiVSEJbQzDmajIO7Z+24061HgFTE4zH8/ooFM7gs3psSc6DP7tLczk/rLX
CBLTUKOu0AI4mGwPEoloIwHqCxadomOEhDUlkjOBxgeoATE67fgRfZtHf0Q+ZNaDYlxnBWQozgmA
UfbXQIkfxDwPLcycoiGJeBdh5NRhJYVqjHOttvyNTKinfW+U4gGvPyFnPfjH8PXnBkQv5DCdZMip
TKHy0h2IG8Qk5oWZUHM5J/Ju3tPwXy/uDjDGu7tnktkP8tna+oPjILZqAWXjMwyxwf5e+4cxdHim
5dZLVmvyXx7i0vOduO4ht9u2vsbKMDDeIAXdnlU7Z/YAKQKUm2Sw6Re2PuqorTU1nH4ZZqeTACLK
8TMr68k7CNndcwSIx89QxX1WrA29RkZDvKOBCEdcSLqZyi0jiqVaXBr7NWhZCST9H+iuzuhzA7LV
1P02FSs54G7Mjyo2cpHiYCV1AJQbknnf+pWoMxAQB+tPpmirO6DnKsPCbQ4nRISSFfRbh+R8dViX
+m6f62RSBWOItV85oHdouzw3wh/TelrUQpi+pgL97iRHhNKYimeeY+WE9/QlmMb5ileDBu1pl7Ia
bk/bTFfX91leip8YdMUi4PVo85wQW3NsnUsZ8hejumAaMGK2pEflIPcGMte9+9QNZzfBmIxdVgP4
5iSNRhORmjE8YuOelFMg5x3lCiwZzNIb/i+Hyx8x+4XalrhCpWrmTAzVPhbvXLWJnoTBZkr6vor8
R2nDVcwfDuqxWSnJx+lOswN2/+G1iUBRHGdll7N2ENASXGH4ECJVYlQ20i52GqVfgeNYlNzAh3xV
jKO6F+9JRc4tHsOZoYkqXoDSjFvrNWo1mX+0p6xclP5N3r+qZwtxeqHYCc1HMSeCrfScXxo24izP
LroWX4ogu4u9qL69ZwFStU8c2rchrr94LGCnQapRqw+WfccXqH9AhRvXWkgqSUY9L5IPQfufW5z+
24/dCk/V36cxCo1nrKtI9kmP2TurmlGS1BEQY9TWcYTaydE4R2EcpFztbTPznM8VFFboVbx3Khe7
xGQlgQbA9dX3LNVGjnB9SnQtB/qnCaRZ/htwwY1yt0d6Tg6eYdgw5QYPmT4wCErF4PIw8HkrvgGQ
99HzcSuoHznY91LEsoJcR0ujTbJfHra0wq6Kzu37XsyWjVTC+E/VWkjEqWrvBS04uXDo8LfTlAJ6
Q0OiwyJhLd5+Llh8q5IA8KrSJoLnRQw389iAvq1hfQq8FAKsxb8hgD0e6Jk+bgOR8rK0TUuh0n0K
RNuWO6Zji7DL/vsZUOgBVQOyFGdP19pQX3/zoOmoHP0ziw2GW6IT8vXxX2xIXKF+dD7TZi8xX4d+
luYSVqY4y1s+a/iRJvx6PgU3mLVSO5P0TxlMhsKs/bTgPu6aTtIPYWDCjDN6PJkJMQfntZDye89g
EJdpUOXuh+NUwKiphciwC+nMGtJAeDXqv03gYzj+liIXu/vUNFX5V0cvmhYSb1goKQJJ4mXKKomR
2694IJCh5W1hV/cv2M60WP3vrIGQCt2Fdql4IgY2DZHjh9aV5X7dlcCStvtPd4BlcXqhddcCN3nA
x405BsODQZIS0Khd1jN80k2/KbH/I7aqOBnOl1UkswTsQsCX1N71nvJyyNW6z3N7E3VIjSof5BqN
u4/cfT8LmxmqDVr41l16txL6fbhHWlAEOMjp7S5Cx5IMM/tvOZxsApkBdzMdZBvMeN7w/ToZePSs
joxprrHoRFWPM7ACaYUt+Yc5U4lK8M07HKOIbDw+8lLoES+uXujatE2Ge3hEl3884ZFtCuFrF18e
88mSmwhHljRgXB3XG3v36/RNVQSNW/5817WrInsKLwg4vJ/YzFwd0tOLM8JnDotVQAaHRVevf/ac
XeF06ZSGleI+/ZuC0zMykjD10E1mJgL69ZzntT3+zZXuW/gIgGACa/ZPNsKlrlXYPa3hpr5zWGyz
vdp0OtYEP7V/2cPJ4Kt6pxpuFVRsXUiA0eFL21JSzc2FCbThXIk/FYWFgKZ+6w+E6pRy6zQVTkdR
csLYUVBaTl5u29Qa6J7MCla15P378B1jhYdvgYBCVMxLkJtCioJxel2PvmUVcTAGeod4h7+Q7CQu
6yXFdX0WlT3DiNK/IDqiAX7lxXdOexT7Z/L7pBb56YMaI727aseN4EJQfA3pgxDHK1tYWeQomMsY
KblTBBnlTQSKoW5whnyhQeDddTSgx5l2m99/NN6D8I9Gv2zOKLnF6qyNose7JoYWfnhuF2g46CS/
6fl1jw4dJZR9boVhAHNBIxc39pq1ltIeB2qr2OpKjV3u5z4cH2yN0PPhQ57M1o7OY1Awc3uRdHvf
0MIQOFwfqUc61LlM20QrwxFAAX/Ha7YAK6rBmZbphdTxP6T8xxI7cMDqjQHai7n34WNNJj+wN+n3
YqHU7ROfPyMWGw7+S7IXwTqaKP3qiX95RcIAsGZveOKrj/zZPFM8rWb4UZiEdmf3qQu02LPKylCP
ABda46M3WSkcY6v1mW7eQesk82prWdrzCVtK3U0yZGzzy0mfjiS0eKNNjqnTY+tejOgmt79e0jVO
TWtMHYORSMyifBx60oXOZkUT+oFTkjz4t0TWTx3RHU12aC2uioxRb3M1Lx9SdpPNuEBgnTOyLhPq
77zA8TJc9VZRXtHrUOo4rYewZCU5ktZ5OdHGOTL1P928XYnBJQGbByL8XPeLYE4xfqLxqwxj3nhd
cQVuRMHngEhgtGGX6Krbjj6zOiRNEKhb0De5gGwJWUIeNF8KMIjKUdGjEUMgIaJWfqXVr6y1E37e
ggxgKDUktPfkOnye5tlrW2/2RocxK8/SIEytNWFaOARyknki0uAu/+F8ejFO8XWpbCSW/nxVj6ps
If+WEHMcfiUD3Jp6yPnGfIz+4btScgaBkqqkJJtBkJJKT5WlL0nadh524Foubg/TcoAFLzEQ1lPF
lDJvo90N0nzERr5HPNlnj/SnVHghgFyyyQJlkRWTWOeH2P3IIeun2R+/3cIi6WVnZ8kggwjCfsLa
do7WCLuu80scEqv9yXWTDMr4Prk1AYAf7LvX1utFUVaBYTuinoCYA35IZLu1CqF2lJdHS1/iyZUy
uuTNjw1Kq4BB2hAb933JL0M5Ahu+7uBCi9jV9VGRiao+L75WFoEe4biWWwdZSEDpiO9pVIT/E3Cu
jCISCxNfmvPdkk5EPJuRnkB6nw4zgMkseJ0Ndj+5x2hbjwJ2RmNAhZNHiLBnJBcl9yK3HCILIzsf
nYKLGta7Rs3kaCl+UevBg+e/X29+hG1+W+mZdIML2h9xVoF18FSv9bherp8KiD5KfA6x4I/B/fXd
XNttxzfLHaGAScfSppOZzB9uRcy4JFs3SvHt9vlI/rFjtOIkjcZ5CWxLjrQeqjhpeSL6egpkWmFg
guoGNqcciWR2UUID/UgtJrOaQ6cIV84D4ysfhKMgyFboFbP7uf1NpKoNYz9iydyCiPlf5VFGxOV9
L4PjwBJPsINNjLsaExMbDEHsp8W5+cB6B1EXN0CBqJXGVcVUd97mjST8FzkLStOeAOLd8XKqK5qN
g2rw0s5W1WzzLfqZW/3s6b+HO3kUSHQ3Pn9cU1+62Rvu9mIUYvVdsA/ZcxM8R+Qy2DlDZ01hRkQb
75nclepWQSt0HDd7GUv+iasqE+kwHXRTj2iyVVzTYJkvZAXHGdWHUYCePY36vu8/yj26BeaQSAZZ
fN5s5Swvg0/QWxplSncb1WRZ/cmf5ZL8Ar6rlhgamq+YCJUGJcAPuA13vvHEsuSsJpTySA0DcAq8
Re75niZaDc4lc20qUkWhrT606NjdaK3Qm87xGLGx+QXRohPdhLYFBkjNfMHWmZrGIgw0OL+uqE0q
XkTW32TaebodYRlS7ti/0xBzqZKHSIgzXEpnqH1ybDWZ5sHXHs0dN+ym3TTZweBWALlyK9l7M7vN
dTw/WberiTp+j882pWo4dgxYRUY5BjG6wW9IdZVEfZMaTtW+5Rq/srVz6QWIOgbXDw31j3TfQQP/
fEpZi8eAv8fmUrapZK7RPX0ZOfzGoCgOZB4UaiKuvWXNH3Mpo0gLoYIBZy24LeDDtB/3KO//NaEr
k9x18dvxNWElms8RF3VNHlHgkpbacMN7JmITsp8kyv5UnAFDcFqFrmEq59OvB3avheI70Jy6BB6S
Y/86ZvINBuR0blwU/LnO5qldOKYTa+3D8RzLXFFAEH9vrUNl0keNigklIGl9fxjrO9Pkhsho1Fad
gPm1JdDNzA1D0Dbq7jsxRTAg6sdgt6JkNNjt6hDGHmRCk8xJ2RnYVjmKnwYLaAWV5/2tTbXGWDRQ
Wc0gKK1eeRpG6L1JAd04bKPwcXXiBbpOtTDsbV8uaHusvYE4CX0cZksMKrSpJdAl+hWkhzSzgnza
CrLFheQMjY8UOPB7Ccib98WxtV+oCscdRrOD4unSfBtewG8cVY4pxHKu6I0k+Ej0B2jNbw2XdqdF
BFiKgMZ9lZt+mMUBAmkBJJXDtHgtVRE8Wqewq9ne+jf9OQ8yIpTy5zf4CpU1QKAf53Uc3zemJ5R4
i4d6DNt3hCL8d4tvW/Eh+ww/d+dzKIWN1Ctz3Jav0wIrgrQltz1o4QEKEKEA+EN0KNqAFf0yuC+d
IlZ89CXJSMUz4bK6uKHhmxToinf3/S087TrFpWdbKuWJOzWMd/qCyuUOpclfm7lmhR0KvyXTka9c
lQg4WnKNBGj5tOl731CrQBWJyZHl5yUG+Ij0d6eCJEstT/c/9V6KIFP1WHmaF5Ln6Nqisp1KVZE7
tkd3eKMPkuOdgN51SuBOka+oVc43IPvwxhMDHF7EHjAaEGnQKuHiO7lIuHdXVlD50LO2pHi+qv10
CgkGb3p8I11Z9Tbag9OY1dAquoHOl0wYR4X1Tz8DGwPtWwrSB8Eq9LnfyV65Js+vytaqUGdh9jTv
pkCxMTr3BuCilQHmVaBuSY9GiR/xQzqPwGMnIrFh2t+Ne6bCy3QCz6jHHwQtPaKdbja/iGjxweE0
FHQT3TqxjC0VsbWivIbEj5jSsabPu7xVI9suUTPvZYrhwNhS8XzcMWwVyczzrLT7tVNJOcTvOiYn
trHNj8ktQz5WtoHurFIHXjLK/0pbdI8nCmpL7p8r0ICT4pvwe+3b/Nnvp2+nwF9s7f6NPB24ycEM
oa9aIjnIlTAxYPwlprNUIN2puMyxjPEThdQahH0sfkAn0N5oPS4ktGlXhXopRGhMTqyyviWxZN9F
kfh2KhcAMoh5h4uS73etRWJDxrhRhGApmeeS5VEOWezP+z+u6JgZ2szThiI/Oz5bD2kFZMvexNJb
A+WWjoxQmoNjZtrNlVHOcm8V2WNf+IceXWcLqCgSHsEiDEGOi3iiNQoXUGzHCirZlagVrBmnxoEm
qSy6AJ4yqwqJyuFssVMZg5ZmyWhnbFa1wbZhTNmrYmtDZb30zAvOekfbXrorXf8Y0Ov6P3ehyA36
T/NcDIEdMoey4iFctdPHEPoAOabHKc1EkBkVM9pW27tbJeGEe41RwoB/rwTNS5Y765/TeErAh9Ea
9hg5fNInyaXkyGPLEgysRfLZrzMTeIJhFBlqOextOzcLzpNZyJ7YU3NBl42LcFL42RVbq9YwPpR6
fkXU2r6tTEVaUteQ2g3I4mfRneZKEZ0GlvFkCcjKkIuABH7B/9v8eF718w3bUX5ElPSEdhraO7ug
qVsG13uElJCGzkoeqDp9LWZxxKmsMSxLa7UcZZFh6ep50qQaNfdBOjJXHlMX8qGanrdepmjKGp92
L49bDQLc5Ke8f4aCEF1AA+79aAMUFAv+hr78pP/RnGh/VHuJIm0Z8s1eu5BuKYAJVfBSCkdGNngH
/ilyiguiu72QseuTpnJbf1JUuIjPHOy0aGTXDp9aKwG3Epup8d8gf28d0oMefllDNgMXsgj+/Kt3
bTXbbtiJm7fKaF6pfvcTKZPGMgEla/QSCKcLf6aCKruihBqEQqaZLLWOSGv5xCWBkkJV/818dJ1C
n3Ne9bcbCE1vZwPtNZexl4G2un1ksPb8qPGtLH7FuLKJeJdFgv5mhUEHFyhfpou9lbR0MLh6gatT
F2OVrP8XdvnY0X7Vss9Ms9rtEYpyPBy6A83jVZeK8ZLpf+v/bk29jWCRqnrCsiK0NukVM3S0kK1w
jFxGVq7f1iuAIfrOLkb7dJ6VxnI+z2A0GmMzCvzNbujtHUUOfSpS/1ud3/jYDOZ8yXjlIc3eso8r
EC0/apKYoCxauJQia9TcXK/Av0Mg7XyfqhKQ8NUTslwnWSII/DJZLDWfDTT3YXGCqTswy/+ov2Zj
MfulzVSjy898bKj9EWsBCjoK6B3uwuOSA0aSBe/1bj6hst/3cXao9Ez177wU9/Chw+KKaeo68g2D
Xz7Luhw9VqSDqPJwjrTazqO6RRZKwjX4QNk1fLmop1Pnv2Lz1nKJI2RCWPn8TMreaTTPWfCDvOeO
aiIXKLD/PGVWzNxhGkKjWKOj0CsSGBcB4SJHaccYzj7Lr0TbUD9ysVdy+bBQPmQ5ZwAukLd1f2ug
drMvR1hFCgDCWaPl0chN53JnZmD34fieh5UNuYd8fXOgyPdFFma5ALyzZM4KvFJPypa1E/IwCtKB
PR3tVxciD4AtacFN88LPbvqwHBpxjlXK/cpRyY0K2HlW/rHVxFKTy4rgXHIGSoFC6gZnegEwx4g0
83JiVBihxDVtA/34iZb30QvP+6Zsa4dddPoLTGpzqOk82Uey39AVoFhYG6L/qcb5wB64epWYz1xk
UJoJGm6xHJsDQMjScEUOxFnUHxTM0DZIWQosgrk82CGx9p8jAJrwqr1P6p2x05C+Ebwhs8bk3Ddq
i3G9WNvXMkws+WJtX7aqdfRkb3AGUjP4BP1dofox2My4ymGbwSq/GnehK1pMFgfvGhcJhhiFitix
QkpO1+VrEpoMmyh1DOBdCvlSKI4aDyZp2MXWfVm2k/WUQRoh1jB9n+mXmiwMFfnEshlo+2unmGQ8
cDlOTO0HviKInCdlDWVjS7vl2PPR1sBG/VER5dd0s1GBc35PrydfojZgYrDLvJOfhoSWXYpNDl/D
QYsh6wCpZmeq7yuQeRL0JkdrKTzneJbHebbOGRukS4sVTAKO/5EhM+Hw/G81l7PjImQb/uzp5yxS
8Bp0Clj1LwPkbbaJKizbbqPC0f1xFztpFn4888GF6sjPcGIHIN1BX/AO2xB9IEWQnCIBCNtmRkvP
DdAXc5PGddYme8uSONeqmbOBu57w4rVpsH2ksLJurfbDLY7u/aHTRjifgZ2lKGakxwX8gKSAqGlB
sdmyHT9+uOL7yKuW8Yq2088JxS/uwKPAUfZhNfrjtaZ+0ogVq7ImyGjulfutFsWS917h99eVRJtY
oYsV7SCEpWvNapE2RQavPwJCeNm5iT0SNaWS/HJIFaW4bo5rYuL0/maG7ogRgMFpLi9aB3D4QgK5
as3ORO6cOTlBbEo2bEXmghXjpxrj9zsDXLLte9KKaBwvhkgelTy5K3w//KC8BXt66zRfM66OHheo
LoPOZDm+XriPNG6jRAnKHifqzwNfBkuWm7n4/wi7+iLSH/exs4WtU0JyJNX4gfNKLIBnbpz5k68R
qRnX632dFIFIwTS5/CkPkyFDLvwIp367Mk+C09kvXwFtUYDQ3Va2GxotAwPmPYq341JGEX5tJW+x
VwRsMsJ9+3ri1xRX5yLAheWeQzMymN84O2bwgmow7obSPvoYdgSY6ZrEAOnnfA/pOrOx7EK+CR5P
4wKFv01BTw9S8g62ISDq++d2QDc82v1CKfsyuh0arPuPrqOkRlLJyBbfkoJkPjqlAo7fO4dJWDOg
XETYBWr+hIEwdwcO1a49pcdpTJwy7n/dE/DfJZp9v7UprkOm9WOs8XQ0Vcoqh43EcYYKvCdwC2DU
bIryL5GbZaafw3oK5xDeWaQOT8u2sD3hMQqYHzWauvjYVvtZ03EX3qOszo06JVM/J9+dENbeqGSY
Q3NL+/xwngZqZv1fYp9ah/PAlP9YrJKBoLgLBh6uyZCKANLZGbIbY/2Qa2C/qyMsVaUqwOqtg6G+
JPcuGrIqvtYF2HhdWdH8qRtI55MeW++lsSOfVeYJsA3AdcSa8RoNKYlIzPsgrP5pUCFTEmJA8X4e
bx6fV616f4+rFlZtDKSluuqpogNALFZUdXV+2SQQWG6O4Y+pVqJ6/DvxeK/b47iLeMibos7l54ZK
EG0r5F9SdPAvjF6+yOVbQg0TZxqxxsnuQFTD5U6XyfSdSGXx4Dno4QvCKHWWoNxOQ6D0iFBxLp1E
YEK4pUa8oL2H9UGvFejRPRfnFKvV1cS1LbP04xf5lQJ60FHRLqw7nFIEsQp8d81Ref8V0GLD7Z2o
WVKSoKXVk43c8WxVRt8cpGgBSgBTfTqRLz7250x1usNgMBjjM8MT974inDZ9AfNrrEgYXn6hyQmL
ESJBoSu8jISmZXRNcMK4LuqS3EvBqdix8k7Q9XJosfNHCof10BTp4leP5mGktk97Qopb7g3cwc6c
xyyt0TAjSbmfmSwmjRa+MhaOmaSONNgXzHPZBK2fO7qu5adb9R6BYRVXSXH72rOMYijsQiswI227
j9/YP5jSn3Ir/3wCBrq6SAn91eZ//ESsQPUetrqPioSV/vwSZU1Bnh9BGMu2mH+b4IoA9rsi9I5B
FCHe6HWQEGVIuJYcUKqTrjnd6lSKgjPTzqOCJWHmaJbqmsziiWSnuu6DKklTEfHTB0Dk8V+S+XA6
iGN977Ve56b541fZS0i2sD+9tVCHi/ZMJr1HDuQDpHHF9HEhMzYRSD5WJsKcLXDrIPE+8sEPTpBO
FEoySdF/eVZFbOTGGJ0h/I+GMUB3FJ+0TZAuanCsOGqXk9LPG5NllxxpnWZ0EBRoT/677uut9rxu
ZtS49UFLtd9yb9Ieu9XaHUHPwoOon6yC/PqF1tAhpwewGtcgFY9e08MKuHdsub/wjA3oINmbvWyu
Rory81G1yFdrti1ES3Xm+lbkOe33QAkv/Qlch0SxAH1J9aexJWn0wpmbb8gejFcqPA4Umyv/qdkK
nniz2rSXS2JlSm8jvxrd2pnDXmUtLkQ8o1rmn2QsQxn8qZ6gtSxliPmlbOsNpJTe6/L1VEzcBwiZ
aSbKKs5/y2taBJXZzTwKnuXoIndpIXlGktOw5Q2YakGtwr2gJwoYif4umrkANZbA5yxoEzQhinE+
D8ONiESJBITa0n9QraL75nPno9TeNwj0LNZg79RBvUmTi8Iah2h9LYMOrtoYkT0lKEnSfg95mF5G
nIxiwuAUsKzd+s9cbqS554MndFJs7aGNY0A9Y2czilE8bI1ncdPyfD122OAivdQ3PdTuOoWnXo5L
ZY7GnpG9JpSSFk2c85WDW+Ha4ffdzQnhGRePifZgcDwC1pmnCFdgiRv3w8mFxh+MmBnTZ8DFyh6o
Hu+IoAclOnhmiFuYCt4iw1oR5DTDOaxWp+XyuijhfcdvM37Oju53cRQqziOiDwdTVnn2SSdx4oDA
6qD97+L+5IMjNpLTGtyFGnAmZzuHXhi1t12KOxIt4fSuKXCJkvRiTSAKUFXB0DLL1SAVU8Hy3fH4
7hZB8+809rQGBn4pHRgljdER2T6+R/PDtPBldy2kY6nPaAogkMG4ILQ5IHCzzHVqn4z8ep2MBBd8
YetbYMxStzxL6xG/HUVQlzOVcjc3Qg7ycYSEWZEnX3bCJDm7iESLBRG6p4+p/0TSfIllmFhmUQ8e
RZ7thyE+VWuHQzXhrs0U9JDHDMGxWwkMgvqdbcLQfX2xXVChbzClwafjUuIrEP04QKusz2fx6Xpx
2Q2HzxBCS6VJi4zHGzPiRjthy5U/qU87xagJD49OdwkRLHQxDDxEHt8t6VO26ZwgN1+J1kNSP7Wt
T85VjLl3u/ymKBwUYmL0JOmBHMw30ToPDksTnYBrJhG9bWmLRfUdfG8fKCopSN79GdwyNTlI8+c0
YqGpzD8fc75iAje3nIISfzcAKR64De+TWchXaoM4Y/QYvaxJjCPKxg+C+7/S6uMunLNVfmE2fWKa
KS32OlTq3QJMfJHvjalsfiKsq9vwV+HCsvVDm38LIxI1/Sz3O26UHg4Dns86os3fLMVTfXeeib60
I3yTz328xJb3VPOkg2lFtvxZJnmQH7XOX7P0GAcvu5/penAtb/5dS3FehsL2e5A5d2B0He5bLQFM
oOPIwwsOI75b37gqF4Qx9CjCWhs8XQ6yvBloyQOaFgBjeffFXZhQGqZxuDTuQGm930mNAI8YWQL0
zkQW/lJI7PNVQ03oNN7xKsMEhXdEdjcHGPRpWFrnNeSpAh9idd4aMs4zP/rEt9CRrzatQnqapqQt
yVjXy9R6LI4R8B0bg5XbhAvettTatM7ssYET+y6cKQpLVpadb2/NOPoAXJx+2qmw1Mhv/IUXHYkb
Kw1Ou5xEUqGy97ZPy7q9Ko4wVRX+DnHnXM68mmnxTU16/3gi8FCk1ss2s/d5RNapttLUVNmu/3/m
6s+hRJZbkdwWaxcTWy1XyjjyRSeNM1VKoXaCI2SdmtkJbxYu++3gdSZenakRl+ozq7TFkNeJtxsp
+jos2wFOAQk3tg9wf1T6ZNTWCNVgmPHEWOlo8JqQQIeBe32eiy+NJr6TTkJ7siJeF5fZaVT12iQo
cOEyNebwXCs/IBUCkoQDfBmyRFZT6MahG4kJEutFYSr8PN2oF6uJfzo+EjHZF/4nYNkkgb9Fe1h4
cBMmm8rYlxGdfsybJBzi+kw61xjnlU73KiUh52TVc+I1TxeqiKuXkVTp1WkNxDF4m0bkPXq73byR
MWzOWsPliDSNGvdeQMcy88guAxowlm3sucGEQHfUoDybBRHm8qe+FS9APmKxbyxQquiFbMA1o9VT
u7L5162AXcifkHr8Xv/tbn3X0Ra2CXQFZ2q13wIDSAfN0JkAjXMHoVAm1V9cl1bMKqGmzmD+VPL8
IJMxldkNOSGV8mBwMY4blwG6IlGYPZ/N+frPeK9kgIcMQ0cwhrDAbSbkOgWeScgMtyZV/OkObOE0
rxbkKUNccR4yXx51LEZKcIN+G4AR92MpZ9ejm4eT4dP1lIW9k4LWWdsFgy5yrHTHaBE648HjYSMa
m2OwEuOaYXhFchxRp+GClhTVHBYsCATyVLP+HsdiYHQvfjYbfwGYNeLxvpKGF6+QuSFxZVjgZowL
dx/vV8BAQdWhiw/EN4wOogJX2JDR8ExVQxbvW2w9LQgcAgsLwIV6hY8j9u+XlNcp850oy/YkASEW
H/noaXmuGODmtYqasuTJwvv0Zyim4zZ/O/WQBLGMlvSRM5uwrXyE+vtgLgF51qJJXdcJevUGWDkq
WaLxgc0/8OPykmsqhO/oYsLmUVr1PhLoPqHnlPASfUmtG3d4+07YvgukYznnefjd6HdbLtM4Jy2C
7INvci4hun5hjPHXKT+b5Iq0fMPV3hqjkCq86OHTySrZwQOAjo5xNK90tCNZN6hpfpK6jZHHA342
5OR2r/FlvMWOVBeqaxEjvPWwviWmjE2T5dRS3LmjiBC3+CMdIsqC3FVWZXN6L2Ft9vY9yU9snnno
TGBeiCoC77epYWP5aSiKzHodtrS/JOEJy2CtxeGZpxIaN0gL9ZiARTs/XJw1MBvJLjkBHJm+aVW+
AkVItnqBUfpmBjO3gOurP7T6eS/MEB8csa2udBbwRHe6u+aa/3EkHPW1irjETz+bpLAIoXaxsioi
dLkMov+OPDcmiYJAruJllC1hroeXS95y+82e3w5AxrmTTmCeOjnkixmQxPzkuwnD705Llb6frJQC
j56N6zqwOnL0HLXxPTTjr7HUp+4SRSb1YBxH319gvQ5xcQTNMctFpHT+4ouzbSSYwDj4VczP0pun
OmAu7YFlbaXMDrmAQTOEvwN/3nU8ruZQ+7YhqjlHxXxB0HGpSkYB4KK3szyYjUK23AqHP0Xjs++l
JK3qyIVf43XmRFamy2xBGyvugvwDeeBqDaBQHt9Zl2Acd9/L5XBcITQCJhC1CBtrVB08HDq5TztS
hF3pf6rurPCrDcP1TRa8iOnyMAQUjI7TtoOdCVPBqibia450Xos16welMD75LTi7+2z2YDDIyJ2q
laXiQ/MiOBSnU4ywuQR9z7DiQ1+AIQRkIIyTjoQp0PgCKuWRvI/kyIpX5wUxKpjTg2qMRTtpN5C0
tYpKBU2/QEYv+hZ/xQN5mXkY5fiiJ6uDSfIQto0oi7t3vhfTw/uajCHUAEIl7YpYZsiNE9SBnEPV
w2QUP76k1puyVfVYqR1aCbMZhuHtge9s2Y+XRuGZECOiN+o75U0NMHEibw0iIudBlUeGmvrt6NKM
00bLNXyG0G029uF0gj6WHycI1MrurkTU2uYa3VzfH+uxsdA1E3KZSjtlumUjn4EfT4XTpi9uNkWE
+PIddEtnoaJ63ULBrWiM3d3znURuTRodo1bYUOM6tepSHb86a9Sp68hQp4AFm131qyL8E91BxZL3
80yJutjeBQPgzgllkpzRQdIk/74R7VvyBT6h7BoswHHJYvcvznIF9lN01wkTRjWlgnvxFOIDd/Rb
mV3TtbpZ1IhFQwOIz7xWLiuFR94yJ6OfRy++nfreD+mNKunxvyH1+el7R1AyMmuG9zHKKNnhjp3l
JWIlqSm1Q21EPQ31VfkM1c+iLVgx9Bjy+Y37FDM05RnGILzWb9M+NmPRTzWxd/GR3efAkMyipdYS
2mu7FVQ9r1Q4iErH5f0/JO76TGuVAelzufP7H/UbkrwTmY3QrdMfuH7OxHLn/JSCjc1YqY3HaIQ+
TFavdzVic5Ih8i12Hgx+HsgWXGcqWVLaz3zwidi17b+60uCXnwpOb5ZhFk6Si9nRfIaNHO5r04mp
zMf8y5H3M6H89d+/WQUP9Sh7Lbq/6UVdmgimvlwnb87We++CmK25jvtHay2N7yE/AZXoYrlv9ZIz
a+KAvBZ2PJinMjm/xpQfUsj4B9Ji9lIiYiJeE6h3905udF35r0zuymlqCbWEWh18qzgjVHN6azod
4Zq6xKlLQ2fG7lVogh6FZrAdJFOQkH+dq/Es5mNG6FRJwjlLwMgp5j7+p5y6v3MF2xR4FgnCtVA6
qkjMu13TsvZLZOM/30Wk4/td/w3rLlMxeCWT+7R6sZUzBlZe3CfKe4Qa25Rebem8ZX4God1tx37j
QRjYKu1svHUb7nl6HnaMdzeWhZJi5xOFBaWaZD5e/wi8Zndcyi+E7gM9Kd/H2DOdc54YEgFuaW7u
64j9rOuOp6aT9N+8W0QkRcVTlfMQIFj/qklhnYlIC/OBN4SAx9EeCy2liDF0nN4tcvxyCRgDIDVF
XgDC4KpE8cYEqnx5iv3wEsCjt0VWE7SBK1mNEj2MqH9Bvds11PpxKhudYX7lyMdXzZwZ9eGu5Nml
+plKt/gA632Zl3uNVCQDwts01e4FUuz7vHRSzIarf6d7pnlTZ+Mnie9U26tJ/va0vmtVPR1V0mfc
Ujxs2UaWjO0RjYmND9b8XtOfX4JxdUY9ARswAGywxG4pwlskptmCHsTFL/5z71kT9tBkgwsSYHHN
FfLQFXp5oGH1PZRKG73vf+qcN0tFWOb9GEWnHHui2XVCEbB/BDGbXs/YTcxyZ254YkBbehfGClWQ
0wBikJXVWRCkI62/uXg9O+gN9nlvSAdKyCKeKvc3hpYmsHae3L18ftdI3mPqGyqUY1tI+b8poirO
UdyZRmVRT98MIMzv0DD9RqdoXhZrns0Pzkx78cpqN72V7Ub9320Pz/KRef+7wCTRAnStBLHadPgF
BLYmuvKCUxd2KC8OVBXwynsB2osZdzsSSXHDlh8hsVqpXeaJAqc6pl+v1ZrJw6mOEi4XZuPMu36v
5aIusA87pjFtKJ64m5xpuImOWeIVdvo93Z/GINS/97GhfQe8IMznEwXM0yOh7O6MVA0QgUA7Ae2m
rHQbH2Rnerwh5+uI0X1ZMFW1fcmvZH4ACLTxVgZoob3Ku/WEkpvco3sEyZFp+Uo+2lDaquy5A71D
ENddF5eswch65yDABdu4RTLwLoXueMlTu5UT96keI5AtjQMMsBG9cRWaImdplmnboJTgtcLN7alk
Khx8jIdZAxCNEvkxJh82Sjcs6XIEiiE/UEHJ5v7PwTO0S6qWXP2sU4SW3u7lRc7B1VvjxchtxagY
vCGs/c26QpjJEW6tZtS7G5HHwSD5c7mAx1TOtesTVjwVQgfnrYRkgdUimXqFAnxXEd/DPXPu7jBP
+gzOBfsZEqInYqq228C6JtLoVMle3rSJ1uB4GgGbcpoFC6DmTpQPvb/Vn3kBSFWpklokvN2TpByZ
lwp22wj+TxOl6yjcmPL3aLiHmyBbvs+FbkKs2ONKUa8WtwS0LQbbPnq/72lLOyKBpwKSmo4DOInX
gy7QYjzRdCetRVflV+je+VNWnFZslfF3quhCNpqPnGVUjhgRNGFqiPh1RG0rt4wDNnsNqUIM6812
pz87KwMnk1SeDXACTOMOuoOgq4E2M/30jkmA09n9UvW+AkpfkqRJRMAIIOVjaMtsiOYunDfQQp42
u1QujYRdIrg5cc2s4Qwi/12UyFm3IjfhwNRi0/74jrVbhXmSY61ihrj7PASREEm6RCrJmTPPVtJH
6HjlNaJ77ol4zVmH631MkQxB6CqzJq3JDLdH5LIFulAIE5hCU4e1im3wrLgOIX/kwxPeWgGYDwc4
k2uqjwG/hlZbmPp2wxWaSWBLZVhF90Fnrnk5JCK9YFitAlhHHAYTc0BWt+QTpY5iofALm+EGqFmS
phJ/6YsgkzG7LbZhqXwowJ9NOd2AOJv09VMLm5nEk6Xor4rO9YnUK7l5smO3iDOYsD3b77A1Cz6a
d/x7b9AjzgIT0ifRxkTGGGvB2yPoOIHuiNVv9QE1kUGhOG4TwEIWUT/IkCVltVYsS5lp3KI4UsI7
kS73tudBKBj9yhvvI3RECN7BsGuE46UVEdaPGvTCK3OFW+/kiQTfVExNjy+TI4sPRyavxa2uyCbJ
hBlLsfAlZ4IurbYSxMDjDp0nXIMZNrgHGVuZazBsWyT0pxyi0f7dThxvMI31UDBLgwoft7bVemuk
9K3sp/E2Cz26a3GBVAC/LmA35cmz6TF0v+dqqoOeCkIEtMG9Fg+qmVnsZJzJOZjYjltxbptHG7RS
vp5Fm8dWn7gbf1WSlNDOvi/F9KbABa1eLwEg/Y3iZaoIjcp786/YXsRSlfR3fkq+XYX09gzzA2IC
KwJyF/ljZe0BGw9ahlZqM813sVM5+2xDhpt6qJJeYmDfF86uqL3ubj9S7EPemOmK8mrDSdrcbhxH
p7iti2vupaU1b7eOQINct6th/S5xRrol7nxTSAFkjY9tlPEk7cADccxZaUdYBkeUewvl/qOgICPb
WD6qQQH7EnWVExbxg5Ty1yMGt0MIZ9hkCeL+QODIWuSrR2TyP8IjMo/kfkLD7gttxVen403yuM0K
0zeQPNKnAShfKiaYaTdJItnbspP4FLYG3ZHNGwgRhS1wMCnJQhbzc6xa/rUC6qbEFcjN2AXWralj
wKA4SA11jy2iwuvfMfwR+jN53YWix+qZnSFnoOCzB1kNTnTAG5N1QJ86ZouRoONWq0PDbJ8pGJ2J
M/JJ6Efv+fNe2FIMqisrFr9B1obWbxGdFR4MtVelGmOj2pt4cdNV2Lxd1kbscK427jX1YBncIXP8
tho8/DmVkc0Y84zbcWMrsLNOpIL1rS1gAfQtIMQ8Sk/Bc+2rRewkYc2grA6tEaRsICfY8Mhj6FMU
4MZ6q5KYVE5I4nsqRc4xC07VxsMgTAiJbsE8w/1Wp7adp9VRf+mT/nPXw+qMaOnLJI7QYSC+0Wcx
+MweWZqlhR3yF0z+dfeB1wHqDEg+4TQRR+xLusKV9siSB56oaYwfbruMw648HkB2XMoFnquB4VEZ
pwUVr89l+t0fK5ePWpNRf2Heg923vx0sHTQM5uF+rdb8WhRLIsRyHaJKYbSBEV6YjYdczJIGVD3M
IueeZ556BVaaxR2cimK5p3tQMqcM6edRfgTQqeEBK6+Jxo7t0ahplhlmGdoRVUa5nzVrHjFxru86
2F7veeR2kIw9dXRNvMT3j3PpbJPcsAvxAPQGyhAKIZtIvfrwFJru2AcQEm+dT38tq5nQTx+YLYwQ
g2Qh8dcX6m7ONMDc+y18pRXjOToYxAkYhR6xXbAAPK/G6cs8ul4+LxESCMqVDhm3QdNpAEAfvj98
oEOKxxKJZIJhyupg2HEAL9zgrEoZEe/7KnYUwZgGNF/S+R14vz0NRRElrdi8RIVjj2bFiDYbyjBZ
3N98WZPPbueDUBq5/hT//yhyPCTFq8J0QJXef6QYRdHuCH2UihFcx3faWdID1Uk/dnAXsxQ+O1aw
ycfWy0HiG3voKtIRbaj4QLdBGZBENv222EDcPDbsxHavUTiFfYYX/PPox5n9lfYiF7LB2zWCYemE
NWqx9I0wQnok4LZPuXixEo2/2s3cyG8tLLNGGBryOB/tixXu9HcPHrZvMd0YqhWmIPzQiukalDIT
cuooClDqo4/sMrEQyDtBzsm4H8+eok0oRY7LryssDaEgc4hM1OL5UntRKeuiP0fMyeOXPuoj0gT/
mJDPvR1oDrqrnPUNhLYtloJBaE06jp9usGudUDmO/Xp8jAwVSAqnNw+/IWv/M+NtFmm1yxXT9Ksq
ghYgLIU76y7LQcFh2Urvrxa2RbTm23dyWvzJLECJvNWCOskVySLhESkCIiTsvkK64u1rVCSzwtF5
ab+t+dpJEhwg0wEzZEREVe0jJt/hElqPmk0IoioqG2rPNs1Kxl8XQeVTV/aD6x8qa7UfEhdPMIYe
5zegmRw4A/OIwEuYKxhSMfQqJypr9tm7bAUoRSRjRPiPuL4diMvI+UYNLgllIFVRwAs9CSg/xvuu
T8P1h/9rPY9ExQAdttpTNntpwdsM6Fp7gOoysZ32sFqO5F8P9fVzF1gjwqrzysw9JvdKeR5ch/B9
97GfNoDB+M+gjoSJcgVGSxLwUReR4qnccVZ7iHOB0t/DFOLNTQRskC07xG6OxERZ+0WVF+PwfeuF
80vfMM0WpS48hnHms5JqBYU/WOnqi4NEb/oprTCdNyegl7t9XVSwYWxycRf3y0Q/AGYqxwy+0EN8
/+EzsYDtFnmYnF3BdnHsx/2UpbH+xS3YU4kAgttPVmquZwWBdU0SV/LCsSJuPV5CHFJPfvHH515r
JlFY7zNn49qtlHTEQIfZn8hBXdpuGi7tfmndoWUqZQechM52DdQ87qkwaSg+w8rMQRX+W9ZzWR3E
ylqB78jMYoXAYzgUeSBBoFrr8mrEU8JxmMzKiH3JYGu9WPELrvlsdr9QsLDYzEX417DKmkTlt7xj
T4TdZY7KXfZygI88cYHo4DHwRDwWyz2X84lkHncfIYq973MFAkMr8WYYuJqYgyI0TwNznPS53z4V
JeV2OLa+M7DpkJtlb6DtECrsPs/uYWXVcPo47mS2b8+s296L/wEbtWxzMolsCU/3Gk5csQlNu5lo
AnEVn0WdzBXikqk1WXHcSvtjR3VYjgjyiMEm5IyXqLj7T2WeN/WkuptA/IEiYZ8nSZonCkVl5fpq
P+8On4S0cOJILmOOVeaes1mqaxlSwtUaPUMH7YTbwZLwfWvmpUyOAZR9WC+r+u0ryGOzauJQfuMY
c7FvLSsPFzJlsi5uLsS3vEkhNHyY8j8DlSOT5+hCWaKk+vURj5NDBX59ZjgNRKSkiJiKf6hINEJF
MyM/akXyhe4AvOwEQxIvWgAcpvtOfW7saUxnbgQkEjYU+Y7Cx278HEKD1+pD0K7k13V7obNrilLs
b6oJpPC2kXOQ7+/e7014ELNxU3CC2dzNOM3N/wbCJSHRyUzhr5nkF0nbUENg+VPhOGBzE7sXaNAS
N2TfXrYzND76NV5/k4o3y2cN2eRottY3RL3eZBziUTWSmoJpKptDehddM7nWmX3YzSq5dMC4gYoP
6oGYiI2WLYLpgxuhJo2s2tR+yPzssQfmx5gc/OxmX5T47x4jW+Zca6OphiaZsZqWDTTYfI3rBiNQ
SVNukGAV5LYsvcCzuVoahyVYBGMATPRXaJCiiT09Kkbot9csJyImSnpFe6BTnGos3QceM2PoZWH9
0IjwIZ5IBoqBP9ltsWOZuH3mxSI6YUKh7N2V77X32KL1tDfxj4Q2KvAqmX9FvJZ2243NBZhKnTb6
rwIpFwAwbMgTmEEgsa1CQBOYJOHvFpni/1bKJM9o7Pod6QHvPJFm28Hc7EKyHnY5TSsUn/nub8jm
YN+aNkglzXnzYiB4Eu3QYb26EvX4cwwMzFqXj6x2k3LMkBkY1lObun7s01wp2dB9IIIMyv8JduXY
nuMh6d5qRGKtODhn6gfu/0C2NoUC0B6aRu0WbxtdE2by/k22dmxfLhrHj4iSEffYZeteh1PrGjGn
wPdY+uE04UMri8i3T6hArL91GO/BZxAA7Uqitq7a1c3iy+/eDfxK6lKs7DpgUlA2Vw2K8mVyAyr8
KYy2V3t0qXv68rcYdVPJGUaqzjeEvYGe9CM6c9eJm8wrAj2xrxjxmO1i8N4J4NHPh9mqWYGutEUH
3dTcHcAKDcaKt5j8NP9wDLYWZIDFk1QK8IQZxV4zv9bGdt+TG+6BOeyUNboI4QqpvQ/QPS+HJyUN
I/xU1KXSBOk4zi2ycI15YM1/VvmoJeAbMGaJuXu+PHSYRNggn/43SPz3iQLYVQo3VuGElOAk0F24
L2UjLpHqykaTTeSTAVqvoWTBT1/+UUHMRNfNPnl4wxSi2G2LLmE1KLkOQ3BXx2Rxfd2gq1CopdrD
D4VtWTpDGHgg0+lPhXDH8NbbbIqvAhpFzpm4KEfsjgRyQxaLdLQQNsu/ZgBqqbcVBuxg+WzBVRTO
5nVSx8IbCQea24nl6TtEbcAGfYbPbOUKQm1ZSt7PETKfLr9TG1Ylk1x+REuu2pxpiA4pmRgmW53A
JQgrQq+iduAFRZ+8lMzjnoSeW4RnwFLO/Q8YSQUHR4jj1HEGJU/XJqiAqHPuhV6mcXr/NCFMDcis
tnGL5a3pTEvcRubYMxXsXp0dQkyrUG7gh5n0cwPcDQis3pp5fq3Nc0U0/U8l+td13NjhHCIhV+Kg
LS3uBou1gKL5NwOllINJkz3mRjiVxEc+7aNF9alkKhh8ja0DqeiogdzbSuA3yo26e4AAnoy8LVvE
mHfAuBks6kP9uUG9fC8imJ7q/+ms+a3BBHBslR+CxnXlCnZCnyOS8rRaq8FdUzu4e8DEzJWrlF7d
wPvlEoYlHTqKksqO2c+h68Fi1CyOzM1cJtw4QYxbVzxKiI2SQwqoqdUesKTowTNAMljt4buA+jmp
tL8sxrsvhUPuoSJCzk6eWeKTZnLgEXjSYfPyKRGDuGgSluYyiS5Mx5VZVP/oSO6+/yJ7yfZJzDzx
B1JZeN1wjZlV0AFEi0Ba5iinbL8FUtI3jE202BSo2Pu3nEnecieI2SPNT570NK8IATZSpx0XWe+i
5pWZrqXWK8fjBTNQXHGI5aiasy1Y5Qu6xS7Lk0wtxzdPFiB8BIR8NR+S/UXXp+yM6ouU3vOA/J3g
ZS3XuDlUkaIXh5AYaAa5o30sqCneZEn0xDakcbLPhJr2M2HwoBQgKZjdgvaT37YPvBYVe08fWgKH
aGhKk27623O0OVUY7W4FTrUrE0IQXYkoDnieD88IHrjAGGh1yhZeVundwchHzC8jcMSj5/9L9ZCo
U79e5efP7/HSeLXKqCtBNvNGvD634tw0j+KqaUMZLtIIp0VKqAtLxoAtvxR2zQNsIgRPGrUWUNrS
IzN4ua2Mx89RhOpjfoqSqsH59povATC24xkUNx198xfrtZkkN+p1cVu0uD9rtg3pkOiF9QaOFcZU
Goq78A/nZt/EvT21WLa9mbzetV2oN4c6f+6/XMWJaYFHBUMxlihgZHClGyFfmJK7puxnqG+zsc07
2fDTyCAOP2ESLz9fU0IC2JCpGLaO/XK54iFiM3vHXBEfHN15bKIeMD+y+gbjeAA0tKEWLgQHsuDg
eKCMIyZFYbLcETBPvnnZTnqJt8m4suENhlqAhmLdSDSIEdjF3ILCvGVl0HesF7V+gjNS9MZc7XFl
sWYQzHpdXXAz0V1yAYQaO8zuYi6xOzU0gpUnB3+jFPPNIi6F259MM5l+1Z8wfqzJDTKsBzRagRWo
MECtwHFNKiii4A0Cy8bvtKFuvGaHqfRcOPGVHHneaE0MEDMagzDR7p93XmfkxCNx2dTl7/n0irJr
NQb/KD0cF5FnL+T5fIaCg6Q6+XTtyZ4x0nw0b4vrfOymZ2wwI2weUJqJBtfDPeoOyjUWNwoDWDv7
YA8ONntzDZlTjA2CDM0me0Yh3Z35ST1GR6gYMK48Q7peAtZKcmxXwiZYHF7VSE2SPFg0kmq7fKwW
EgAPmskJE+6jelQElefr86PgUvH4ygjnUA5a/UpzYeIe8p1G+epb15v77AShjA0KNQEbFpBlk7WS
/7xAroJIzf1Nf8lASFYzpdlbZH1S8EKdKRrrlWFQEaGfJh0ct33HR0SwrmvI10JFCzSnIIR9APSw
HKcJXY0DNmzH0WX/c+KIyGA0/iUPYpjn54hXVWilRdggmLawlAto2iPlheH4TUpVBsxjJlLH4xLk
ZbQF1q+BIxWQja4nesZ9Q7Ed4F9L1rCbfsKn12UA8FsgRYKIrVBXPRC7JjnbLGX8iKw7Rweenoec
kl/PclPKiPQbKMtuV6ChzhE/LjG8AIrU2n1jG/QjVZL6L3cZnVfrz6jAKrRhAHCuD3mAPG2Qj95r
lEp4OMVx4Oa21lO8UaXxJ4ErajeBaeIdLLDbQdsll6VP0GDcmFFst/qKjqhcYwh0Lz0sK2xnaVKU
4UcfeNuOSu2hww7thMjyPKgals0EL7EWIK4C1IS1Tx+8NbdPcQBDHKEq7IsGQyhc6Is+hdL3ssb1
/RpTVKagIjd9JpfQau7etkwT0iOd/dOaN4j8YdHGFkBYRQcj+KQnl89NYNaEC/EK/a9de64Rnghn
UoDNJUWj6/OXDLMh6nlaTaZHsSeb5vat2r9AXWBgjjGQV1xI1fN1AjBAGKxMtGzwSs57e256sVb/
F0V2+5KYkGxCZG9rm81wLF30E7nANg2hSHZP9YsKILjWYEguern6uzgDxQKsrsNN/dBpmkShNVx6
zAYMRhyYRzF9pmHoY1+zIFYnH3QxP9YRc9njDtrW2ANglq3E9QjbjJ0hq3joGRXiwLt0CVLpK/z1
eC/bqhIObwOIXJGrtNnfVC+yDhJBrV6huvee+YgtCPFwK/9tuX3T7jlcW0lRdVJzU+ew/AlT2iQE
ttErlFiNp2KyvpWacRj7Xxq7HJWTLYXvVuE8XTh1RJAJ3wcZ31MJa1PgKq3JqQEovGKUgTdZ2dqD
jzSjbGKUCJDc30qrIFJ581M1uTmY+zoY5L07WbYEGpFRRhebNc7Mu81cUDZDbPXYgSvFfYmf4n2B
5Uhcz7Z9isLTtZycggoDrRunCIPle+wCKe5Rxk7CTxrx+opsFlCaH4yGIi2eZq/kDYYEqeXkaNAH
VrYHQWFBOxT8mEDAs+p4PBvWiwfJvpZw5+4DBd8ibhRzFTXyWwXgN2alP1z8B+cORk53NTwHLQ9x
AKi0Qc7VqIYzOxPQ9OIIcMaFzvcR8enuzyme5nHQL13smzHiFVkLKB8VsjUVmoCBPxlwM5mLNeAM
B+1E3+kzOFkwCVN3U7s4PqUsVQZVhhBc2p20p7laNBNCqMHIukAgMr4b/rCAxxTzpOcg9mqQA6Zb
q3voYyfCG0VzRrAcYWlhYkKlTSO4B+eINgKu4wDdU2Dd5mIgKXUh2ceLx+QWTKN9S5OlIObdqAbF
ABtxRU+XKZq3JfCb+mKadbse3/Z4BQhU8bDDnooQhVQPHwSm4tFy2OkyR2e1HsCo01NKCTzcil4y
L+AvFCWckkUGPQqNwshHpL1OlSCR9GY1vU6DU4awnqjcIBgVfqhVD75p5Qccc6QLAEcBv7D2+HOW
ocEhBNjGD5ioApbQ1bx2OX/QgDYIJJqeJPrwjAC1BdZaw90vafogluPOnUTr7GNF0uDC34Tux3jy
R2nXfMLsNY5JTk2KVDpfmV2OjHGpheHa8XH27tcY829+sN1yUTWFkK4XQCr29inqjoJRbN2ZDnpb
OAffFTkDSmP4Bg1zK6NGpq/W4aquH5c35oldcdieQ+l9MQPqWDDa3tUVzX+lAfLXbanEwEO2Tq9F
RT+/JnrszJMM+BkEiH5GctoFFD+Efj+JEI4hrGdtNsVuTQKHVFVqfwExIXcyJCeDEoBjzMdJi48O
+ounQvWa4d/9bPEfMQmYvoG9TvOk4ctrbi79nGJp1xBo59gn2obZuE6AicNDxQTbb7fdzPsC8LKb
dnA8tDrbfayzWb0Q4oDmz7tbw3AJ54WfNbJRi08ssEXr/j6gqAq31+6krRhSXZjktcyG+X6IEddl
S4nLJnnqTfyrISaTjsYWze3sByV0gbezNRfk2KwH5BBqcicYdL4DH+ayEkdIUb70q6A67YngmaAx
cyUaSJ+3bFnzK0eoDs4l6RcQh3XbLaioH6owrO9Iz1YWXJ3AL6jSOqKg0rd48toJOIE/h61fjFAW
6kI2HKG9gTlRnG8heTVVbZLRjJr5Zn880JLKI5WIWhnCWJ7A0CpTOvR4VHL/2mUDvCYuvRdDSFau
pqh6O+bOTHwzkTAGYE7OQTrFjJOZYJukWoo+wmVL5nrNJdzaFnhyTdTjYUN+0ykKuM69Ybe1Q2Ay
fvgrjd1If9oYe4C7R3BiASfmkCoOYl7NiLKPLj0xTgEUaxuDw0/B5YoqGCivzYrNg1k040fOR86B
OR5YuBV43Ca+KIfE2SVkSSMCPWGNivaxKGdOG31/wm2O/7JoK/0q7SUV0AtBCqjZYdNDhqQhDJ6H
APBSMUO2nqypz+GwiDdMa81uCRcnmTSlD2ZK2XMphdGVqfsX2zSPBU5/kTbLe9eWccSQdxd1tLF7
LQ/bsS+UyTzXfxbNvy4A3Opo8ck/xaDJNX5ad0aqNldON6p3vaq5v8obqJcXaHdFawe+O+5vLqLS
2Z6encZcG5nL2i6qvBaELWhaK2d5zkRTrOWVA/pxtbGUJ1YNjCD8BSlW33CWuBpCTFgahY2yeO46
qKKS1Lx2OOt3c+lt308hxaYXN8evsQEhnrvMj0k5SJ8vIeO3lgb5Odt+BD9QQn5IIm9RXRfCSNO3
WAdRB9ZvaD1JMvoJZvRhuNwU1W/CWFFBiz0pHf/RPjGAoFvX54BqIvaApa4FaKPyeVGrv4Q6Dhjp
yUTWAPXy/pSSh/Nrizetza3Y7hSQ0rpSLZsN4ncVsQC8MgW832HH/qnq69X7cYq7Miq1D0uxTscV
G8jT5l5wI3Q/28pwGKrJZb/Jc4WYyQbfjTYp6Z7o3Dsw/KHAQpv96HcMBsbG19GUICsFFpH1zDQX
ovhJdSt8XhtyWHfOatNyH7JxQdkUXyxtiLCW7f4cdEETr1Sp9uAL8KQFHyTxeEV6CPa1oXJmQccn
mKoS/OfUbMDrs4EkqZ2nRFWe2hm5ZJcu56u9Tv9bEyqIXRlGu/8CIQ0d98Vu1W3AmWozOlxWTf78
UsGs86sHmg0is4xpKgA4911v6aQ2q4olku0xk6fcAokp84q6XCniq24OENwFTlDPgW6uE4AH+3Ml
uTWjlfJa7eia5AyP1xTsmhHEbBa1HD/EA3AVQamTOOEJPFyC9aiM0F0kpjipfdN2UgT3rAga0rY4
BOOFVmS71cMnNk7UaZ4mnFQVHMRrGRW8Q5H4GWVsoXj/0ZK6trCBiWPWbqoclYVRvwb47qKZGc+L
pmGg8KO2ECD/pO2rXE/SV12Bzm+hERiBJo0gAPpy+dLkrLHWzuadfD2wpkk7CNqKinPzq0cPPMKr
L9a6RaEIRfgGFun8+5v2pxrnlRyQsFnEvRCiNbRrwPwm2dCSPONIvRvCv+QGvghar332Sb0CRcGn
c6sXD2xrdB57xK3N2CvhMuvbdqlK1zWb/qUV1raiQigB11H90fXyRnmfOdv2b6IemwZjCl+eX+O4
BoD781WBAZoZdwGFRI57UP/7KSSc4JOs+nX3Axm+G7zK/z4sPoaND6EjS05oi0IzWpkSJstjzeBy
FSK2+10gqldvJD4yBPOoU4GmIoR+0p5YvHAlFZ+MbGv3TwJtdqyG2Em58ojxPumElijnNNZaIvqz
55wF3YqNAto3u4CQ9TRKo+zJwVHHw18C1MDVgwqw1OKd4m7yEB1t242cP7iIjLCzKapu1lfLV7Bw
Lex64uAeM593mY0pvHISupX2hl8KjFp/jNUurtmzjXRGXyvPtxUgFYDrCvDx0n1VbMc7Rv78S1zu
7TGqKxtoNYLBxBJ3GEppSnNTAzbpDPDzAZeE4jwFpH4Jd1gsLEbv/IJAqX04XenOPkXR0LFrgvRQ
toe7/hz11FlBF7gAernCSJlVAgzjIjK9PficiQSvWUCUOeybYBuW+y7vNvGlX8kzodvgegVKauGt
aP18IfPBu84GNmPnXWi1I5rGp7xqR420Wph825kivKnyU7D/rNM9vfh2Yxy8AAuZr92lF8c7vjhL
DNFC9PgCpx0pmnKmRO/6jyj6CS8NACotHr/EmYh4+Xh69Khdq+6qeiASbPGErG8vELxx27R8LgGB
qf0+v3kwStk4GlWLOcbQWgnwAl9Q0pqwq3gKR6KQdwg/21imwUCSa9uhaJtURyD9qZA42V7lzvZe
rlxjOS+61kZbadNhab9TadNGOVAGFQXzBYDFxe6ivT0I/UOYDQC3V9vyo3Xr9vMtZPDA2Md76tQf
w2EU1uQbRG9UMntYHPF4oZIIms/od5k8m8S7BgWtzfSlNNgLP9WeL7hgjkDi9Cb57RTFusxpMeOe
apRqS9dvCbY9bpOaH3TZMNp5f65vV2aszgXVe8vqhoyIcZ7zcZbG6HlPhx67U5krpPEyDIJXk6NW
1OuvVQ9UtMMt8iGPcAi6JEXm3Pclj5TVQ8R7IAmulf/lPglRXEppphb7a7iu5My5ZcVZipZV4wkM
Cb4s2lc/Cc1n6s16hCQLqmoviMeJtFLmrMEIusloZRtvtv5T8K97cdfVc30/y4yowZN1K4JyLkaY
4ndMdYnJOqveuoNBCx3O8qyrajYQ4rWeThtJUN/jNAPF0UpyDQkQk40LI0kGjRJKSMsst7rO2EWk
1bWbY2nHAc0N7jJPyoGtQt0dhHUprR8GNW+SPLTCX+g5+ZMVCrqNwe2YHQ+EpDad0OxGJ+PO2Zbn
esKtwd+a+RzVJ9WsRuKZg1o34c+qcKSAdIlYsoPnWyxM6NaHJN7ZoHWNhdSlI4QjGD203KAFfeEo
D8iV7E0aQyNUsxGZsVXyIWrTMquUfcAfvgkY5rjgLmii8jNf52EdutD0gtj07IqRiB7isYKNNecN
aWwQScMiJO36jfca25BL3D0o7HneT3DuajWijwI1Njr+eqc4NiD1W+2mDgLR7QEIhRqZ8C5RNn/a
wSzLu4cpS/Hv4oJSaMzkyqYes8jq2ZGVn48rWkwirzDLT8SpzmwV+v+xgyJoFH9zLhlgi2oWzE5b
23D7njy7BNLrFt85LEVmMSe51mc1YRMvQN+h0bojH4YVusup7pnVI+AIYjbG6yxkB0HUXbyumreT
sIfoajsQhHhBE3msCs8/SvND6RCWcBjgnGfoZZKCqyVZ0QhzJkMzO5JzH/L6cvcUHvElNfaYz+G2
suygVk92AfefhKjJgLEX9V4d/TcMde+MHweBN0naVk06X7FUW0XUdS0MGdd7Jggt4OHUryGqOt2o
p9Wko2ufL3b74L1pyt0HfUU1bWupp3keRVyoyFWSF+U9f8ldanAuUQq90Zx+fLIMVqbjA0POkmB/
vTTqjJwD1eVnvXc3ozzQzmS7dKPjAig59+otlF8x6c9gHrDgC0rGnCnEHiLGKuo2qTCFDZ+e5FH7
vSrOa5MTgzC3n6OoDo9zHLpvf98Kku8QKLWG8OGilHXgpBrCmeJz2jgjgxTB5EvkGzvSb3ZFR7QJ
zg+KK7w02X934WaQQTBmTfoFtdXzWUFCMs7nCkQDFCvbE9UTiEB13FR2FePXPXQlpn1sAA5oMbpy
molY9dtnkS7vlzjIYXnqFdDY4S7XcWjb9K7RCNoIAQigX+krg3jZeL7fxQ20NiUTA8Ful3OUwKvC
I58GxWc14AuOi1i/szaN/HSH+SuZv4SNxKYadfmqFQKFIKG8D6IM4+VwWVWHXQyylTPRGW5MJ0Ah
X2Dch2HdRFf/SX6vMsyVJdzu0pQXpthH4sXCwppAN9sP6xBfu46cMYZaoSGSuB7/GvbeKJqm6EeM
rfVidEIzTGwbT/8bCChpMCbVA/5ARNCVl1KjiDAFFiiD5V8x9/02g5daTgva+yzFVB1Sx7vsm+Cp
QS4x3RobgrR1tugh+SnS/58y9LL0qQF0HZDfTLixwqfkouC9ohnP42PFWHsfj/ptmhvcL4G8gQA+
vaT0w4LuCB702fdeyzPSkjM+wRHsesO2f+Fu4H+SqnN9k4bXh+QN/yh0LP5uVlEeF8RMZfMcwzm7
0KikOmPk2/+HIrGeiUp6sLX7FgjV9nL3yt+EQ/4H84dSo0SAKbi9wXSH8K9aBSv4DwbYoUZvdCzt
zBM/BF9tTChS80KIPYOefelI/P8wJz6mIgE8PiKhbRVPtHH+c7yJKoYYIPL+insddOJm98jbHLP6
iXeWtl8JQImWkQMZbbf7NW/pht1ewaR2LZYj20+aq/HsU1sHZOxwwVqI4vk5DpMqjvevPgrE3tcO
LzHIiCk7GmUF59T3NKWwfoNKqfhXE9rXJH/Ik8jMGPZBEE/VWMysjUt5o6ThF0HIUYHTIQODEgAK
TCMJMinsCKBicBngPz/njxD/tmX7BMKOklIGDWWh0LFbhTEBjxdIRhoNXYMUe+TxYywQsC5TmdFb
PT9rzRTtBll30DUwqZLY+ujNH5PKi83wMFL6Hd87YGpFGvwmSagBCOTAti3EjVkf7WWcgcPKa2Xv
CT3dEOAazqvDCTzY/q27KjOhWijMbUC0ppygHZY8RbVN2DhGKN69wC+XkyZRJLFQcI4sPtRrWvfT
MLSMqpbGXJea+7ls/p8pgrVE39cncXHN5FeJhDDIUuXKNfvWjsKvcErjYhornrZIghTEgtJA213D
EfN5MT4QdW7OwHyAXlCKp8W/9nhWmRw51CPFl2yd32dNDzatQwUvJNRitz62+NBhy6UPt+bwrgpv
3Z6hML6KPuOH1kE5jAwyyP4UKQiQj7Q3b6Z02gtBdAcbnQF5Rs8/BpWE2VwWvlrz7Sux8Y7wCyCB
V5IYOF/bq0OfJL7JcmZ2jqadLEhiLVoUKglZhXD5Kksstc7RmGMtMSq+NM0ajGwsIHDHVAzH/lzh
5dc/P37XsC9M7FoomTre5iNT4C74//3yKl6/rsvYZJSIOjS/o5NeMtf1yhSuzHjIVA5WjDerPfzi
XMtGf0fUcA9mLPX4Gja7CyFidZT/F++qgE75ipjjO0VFuyvpfUmU3aq47vendbaBV9cTwqLJD4HR
EHO6su+VK6gQvJ8dw5KkuW+vis6m3S20SG5OpdDWmXDhW9DeFg36PQymZw/tuQCDiyUaVztH5scF
VrqdbHJC/6kXwnrL7LMVGaNKtDtWT0B9uGmPFV+bWX7WqrIRxqzu6qjxHuMMjITzLb2okwWAqb2U
zw2CRfZvLcQoNUFO4KZZ0aSGHJd8PAm0A++cbhkBP9U0MDSC4swNOLZfrTIdpgEcrymCzRAK6tJw
xU6ffJlxnzsmCytkgkwNPTdBULSHqrYDyj2usMMa+iAkommyH03tIqxLyhZUndDUagFpCUgkarwa
vBukp7vzkNWip/p0+ogwqQlztd0GhOhlQMNzoB5lR4h1xH/aZcUleXhufdVpy4sC055XkPIT+z+4
p1jhaSc/7UFnEeBQOLkhFMcYVg4sK8rUWaSddQLZHxyPu6Dd5Hx1eKb/NaVYXukYz3135XOJJWtH
/xkI5+JOme9M/WanoYhlF0z5Mh/aZWeYywelqxDbFhWv9CigBYgHqTrfbs4FWgOAeKrc1Oh46KOC
91Lt7oFnWQghth658b0aKeJEQh3v7iH4X88jQ8iiQvMHwKfH59cw3TnMbg26bGfxA53J7MTD6nOl
Ywk7rHngdVPdddVvvIMBzTvt3XD5RdW+OBx0HUpDcLyJgRDo7wpXUStQf0NWpVDE3aDUpdXW3XLy
Iy/xPDzQpYmbano57GZ++v7yuqRuosWt7X+oVN1BJAX1zXMMn83HZdYW4Un/fxscqkwTl51aCL8R
jQuxVc5EtxZj2oB/BGCqdvJ2oMXPFNIjtpznzrXuqHPh83Nuu0KDDkPx+gt4Url10bhab6Hzv4V7
Bw81/QSIxB3Qm101dfDfOr33xCrKpFnEEeTlE3GEZxu0iyO1EIiceFwfviu6/Mw7nM9ah8rHOdav
jKYE0LFH0yPC5iS8NcSpeHmXPSN3TeuLdKG4yX4aTt2bx1D38QLwmdsihnokBRWYDazu6X/NnCZM
GH/MWfDJf3AoVQrxGct0rLv5LA7Xq2kwRGgE9nLCTHAL3DwPlDuqoJCFbiPa++d0E/Nay2f/AmyE
L9+u384ksfQuzSLn8gpNUDrHpBy+EGbsO/LC7GzoscneTw7bKclQ/gJUO/bpApDcYkOAnNEkjAM0
Lw3CgMGJLthElN7PNcWaaw2uSDjmCnKwtfNeZ3hhD9RI9j0kyOOMfnS4Hf4VwoKB79xUWRt+w0PH
0wKQWdVLIIvlTFer2z9CyJoygInnBKuQSNi66j6PQAwEXpY2JuNNWItWgk5uOCgQJiZhsR5La4zn
FXo/Ky+93Jshz86HKuUxDP9KrSKwtGKGvYeyR2hGxRFIW6SkK9ki+Mk0+TeDDP5NItvMGzZblwp7
GZEISCemfE29qpSN+rcgF7GRpma5ZjNXWD2XaC5lqSsqeIvaG6ySKAp8FRzWmkiUacqJ4zH/tIJk
ZZcPQmTvm/fzM2HjhBWeBOsTN+F+NB3NZwzBbFktbpbU+9hG81uPcWlvjKPvEPmSjgtvaBLWicQ9
U9lWdGiwPm166twEvdcHlf0qkOoJ8c9wRL4+kiI+DTdu3/JFvo1sVj2SSKpYrVAwwYz95eiunYIN
kLe5KEeNiVuVuWIMUmB+77jdbo0/szHDcjtfKomlpgmqIc6mhNzjDolQtI6vUlLrLBSPjovAGhXp
1dp6DGyIs9u3cwGy1BHfAUtXViVf8YCd3dS1EGKKpXGh5DvF6Q3su7z7+0lvyDVvy6Wr7RmEsSr4
dHGVNyBMQr+7+DI/l/1sYJV/ao/8QSWgVfUco/3to+5bn7fr1+4pYKOw88iraoyGpGPvKv9o4sLV
eAfqmKy74WpW3spZy8ukQRed1iraGn6oDsZ63s09Q9/rxePv/u4ZQdDi8mHI6n+4kV2OEhpZMvqv
VOs8ExLzVr9xfHWlNhMinU+ECaFPNS6fBjN7P8h7Db0X2zzgOXsccZ3VHJf4ku5piWkC9nBXXF6L
EZZ1HsiX6NA9zZrLLpAeMROz3HMa44pViJ7eyqlDipZ6FZy+nEx96q96K2gl9lZc1SBJzyJd7O6W
mY7uxUok916WxgsilKSzwloa9co6/cGg3OtnHEZOSsHy/UOoQ2PmpBznTC4WPH426alIoG1AYbbn
jd+uDGvDE2xk1PYDfl68z2nsW1QcUNokZnYCLohZqgn27679PKum4/6tky01RNM3E+IVGJ6kT10X
a0okkdj06thKGSDb9lx2ZuskR0pnhh9s95HFxWzMii/X46C0g2uYLc0n80NiHTR3ldqpYD3QAQxa
EXa1aQ/9Zlx8QQcA5J5QbDiZvFkmw+OVxZoIWKRuWgJub3S353yJ3LtRvuPaf1ymhSahyMRyH7Bx
PIUX3i8/pZELDn4X0sAaLsb01GPhfFMPmV+92JYVUCZgwDxVrOiE+QR7YJuGqzRJX/npF+vvu/b7
HQ4n9Ss6XWJ9J9xNpHJzYF5kXM0l1QvLsqOJYNSQDvToj9ShNzWNbdce5YjCdIs1vwsxnqlXiFQj
HM4u5so+sBOIHi5SQaDBvISG1wJqbmGepM7ToBPyC+OK63IrDURM3SKuvVd1zoWlli33fZH/xS7w
jHmLZqgvpAdnYmv66IBAiKDeMJDKaBtEY7F8M/Zboto8lEABhcY7ZuMuvZgswwYlEvYRWtZi0WdV
WHm8DHPpsXzcocCBHcWAUcibMiXspLpKBSahOebE/Ursj79J69yzl44mcG5Y04URLoJT4pR/TlGm
oeVrkX2CjjY7p63G9JiITDSrNXGjnNCPDOvANHc+qqWr4honoD8T7oOWdfmimsymEgSrRYQyllRc
K/0G+um8DTSNesZ0uNcx3ekbSHOCwVYp03u9vNJvaW+sOlc1RpV9/4BZpoEunnDwNOSU5KUSRVc9
D9pO41vtu2kQnmAaZzLtCZA8goRzPr1zUOY6sV5Sf3imkprb9+jOcskM5vUOhVoVx9v/o/b04Kxb
TFWTYdB6RR+qyRfolNbX28nWt4pi/u8q0OmaYUnOEdOms6+aLLPQMELMxWcM2PouG5j6uM0i6VrJ
kYkJJXf0nfMuI29045Oz3z8fCdIhd7pZ+/uXTbvo4lP6lld3939WoHM8M3+35JpZ0ntFpVQf6u2s
DM6ZJF9bmxhOju7IMSlHjM2pbnvaopKHGoEmvFwt+xMHoUiBSdjBNj8IhNp9VGjiJXKM8hzlbSA7
IjkPF8ziAbZ9FrJD+KqOrQYIzm1hLL8hKbNmdLoH8fd0vlOzauVdAy5v8gq2YP6wusN/D9n6bLzm
rVjH6qQdaUvK5NBzeGkrgmFMUnpSOtfH+I4uaRdpseAub/kITBTTVLWvculhYjIbjj0T/Yfk2i5e
6HFcAmFwAoki+8JTNJEzFSbp7lUOXp2sb50HkDB7tMpdxRNdleDkIRwj8PhXoL8YVAVFUlBsJ9Rx
gywP5SlnCk+6intMg1WOP4Vvx2eygq6H0lN8O4C2eNVh58jIL6XD647yY1nSddPd1VhCKAPJq9b6
xF+kUsaItLf2UNk2q6EUTj+Ub/pyzBV1rs/j4Jhwy6//OeB81HBFifggSFZ25AngYhVWjBk4/QD+
QrOzbWCnwezfM916T/OlYxIJmKwF+QNwHP7FTCHA7JnKI9vGCU2oZ5/YK5udeEXG5InW7WLgP7N7
9zOCOSS9esnUsFNrTTGjFRepASwXTK6KqZzzFVUCQHuI5rTlVnrS3vB/MpKrXdVwCOxZUJLUWy9f
msfW8BPUFwxqHHi2SpIV9ZqMogVi5mrTqZUY3K1GA+lWD5u36pOF4eIStNICZ79hIfpGh6JsmbcW
n4onPOs56yAjcgBciy8hTkCBDmBFMf3PKVJHQ+v8qHHAfYy4EzXgHc9zvtpvqTGmV7WYjkTePaAh
uUkrCK7WqXoHDCdvf9CPvuWaWflBkmgJTtmMx3AwCYbACnD3PLG/c01Bn3a3HVx+96nv9erTM+OA
JePtwHiLbYD1XmJ3I2yflaGzB42mQWWXFRcy6XbzSVz2hU3WycRlwPqK9p+2zLVHoZbWdYu5oIES
vs2Zr+e00/pR7r6DAhKovkJiy6pSeB0ONpjTMznD5aF75zVx7MAPPTuAvq0vhrbJAgiP1RMXuNbU
EuQbcvyfmbgLNLQAXVVHAwtfoIM9n8Mdopf+RihzrjRA/UfHhpKbpBWD7tYl2UgZxqRHtyZTtLfH
7xAoL2MSMQ7LwdblmYY2CC6ZdD8sU9pnmzJTigHBCZrZjV6n+xWcdeVe6PXzL/ExE+Ko6qtsKDeT
rI19Nr0Gtxu2WfcWE4mnVutRGN3xnQPO9U7c1Vuz/6vAc551bSc9XPapbbE/jYxTV4mO9ievtMHU
hhM+GnjmbnhalLfWQB6XyeWrB5k/BCgyN3RN1WXseqfIa2Xn8e0kVTTf26OzdW4pFKzzgJSLoKg+
IzvTCwE2LXsHBMwqSBS9dYLc+Za0Nq2rGdt5iAL8iY/4/Z03apWF567eydnM/1y9L6RRuYshqE/F
v7NmqidMuS1WQTwmqS1Zm/vxlk6qgVhcJ+iR0xfLaTjerB37gDupKllDE3hJaDaNPRUjZ7TZAArF
G83IsbYt14lq4Ehx/ofrYTTO4MTDPb82hCcVhWpGhoFbZYRrVmkE1+OKMZou/FoVGKz00tMfunP5
J/gvRkckgf0DVVxcEx8XQtFUE+nR5aH+nPKRUidPz/ga3APgUKJcpAJXFphXXthaBBudjqbYprdo
4BkXx9GR178VFlzpqgSVMc8ns5q8aDqWyVJkmeXj+rFyc4pWq7bSexPFBiXSthBTHG2sl5UH52w/
k6bNJEJNeF/mTMHDEMqtkKcls1DLLUnpmAgay9j1MHW2zrcVtm3Z0u/iBhJ8l+EpY1VQRJSYtlyD
5bkeZjXixmO9qyb5+eGi5OmBJ98FQeel1ojOCnmUQ9AvgR5pJnohFjqV5V1JnIkQmDvw+8NXzbRo
wfDZg/HaTaRzC52cV8ypJiDnlTJQebRycueAOo4boEwu6FNsCDEaasXtFb1YwswiPQs00cLkFt5Y
UGJ6YSo83T+oFfWSReXeo0FA2+A4/6K36/JrtOeDHxsVmrMyTQjAXPD9NTe/W9s+UtEQe8memH9D
/E21KdN5O9PeDpvZLZJ7vxauN1SFJ2XfRURM5V5PMlzwBdun+kQN4vF8lQSbK5kQsJJtauvyHd2c
RZ9Lz+T0xmCkas4KT4dfBckloc9f9d2M4/Mddxd4Wmmtle/zOJuH0oYaCZB1E1slIDKJfpN7KlDz
T1lguBZ6X2pcrPM0Q1WuYJRgM+WKiLV0Ga1d+d6wHY2LD6UWAbs6P+iKebmxoY6yurVe0mFuChCb
w28c5/IOUOvdgsV3qgK+IkiIaLRv90wuy0XM3GmB317vr5mEhzgzJkDU2nCHudtPztlzf37m3GLF
Ehxfy26E62xCfFgF6Ra+Lh6kHHlcK3Mupc9Wh/hay6GTk7zbPhsewuZk3QEUiL/uBYh/moihjEUa
Do/rhOQOsvArD2HmWbDh0ZAc3hkw2cdCfFD8864blBkuAt0zB7HVtb4ChUXvjBeWGna955p5v58Y
6RHt4Q9niDFeLHde9VGZPL+mOWv7lUW+hWPjdPAdkr63IgRW6PAdK1XSzQFvgkhi4KhCWYtxRHZ9
htuVvCG2cWCfmmSVWpTTU06QDKtxUKdvgsX5whXjxatkmy2rmtXNCUyYaU4ufYl2rAejwudYYcAs
H3CEfvWrKtTcKSoRkCUs7/bLS0+Xos8P7uxkxbHxTteB2ogalnHpnAhrgukTClrK9RXbpPJ6EmU1
BajoC4kNQhSiUER0w3IvTPF2JjQxoRSNfvKBPWuExYdi4MMpg7I25p5H81fnp/+Wq3Rh4/BgLAl4
yZGZjSKJLmibIv4+k5j2oWJRAX78ncZr4mNP/8s2fv2V7KWOFfaPgW8hR2c4iVtdTbdHeU7MbrHK
OkSSPVArJQEp3c88DX0Ow9khzYHQG6CxFVLupTgh0Um5Eqx9bXrxBCHyc6y6yRQFbV7zaPBKPL+M
rakbVZQWGRkxWdd7VhqV/hqAy6zY9JPtOwuGULqggUsBWcDQGP6KQQKvFoGYdPjwIdrR2BZXB/S/
VBzrpNz8Coi8L4MZ8T/2eNleW6b9oKfzPMsUtEOaeC5anYrhlogJ9Kf1fj9B/eooL+MAK1yFIkKW
ulb4Hr58M48pgxEJTqrYLRLbLjl6HHmWYLSMcSwtOd1eEaz1S7kx0LFX5mkLRrVQdYThN2CkR1hv
w4diiEHSDJn+R9nkaPlGhlGtMDV5osu9H8Y6BhLJ1nhruV+sn2m3bMiixc/OzB10hz0BOL+ohyLt
AtNmpSPuQX7R+tWjQ0qAbqvDTzIf7nFEUSo1xq2wBbb0g7+h2xJnBuujyqCdfzx87gTjnKAWfPi1
1QRbwzDTXi0U9h4TfMbDeUU320wvfTjTbw7h1YQYiecnd1MiKRSqjsJtJkLFhVVzlvVATE/N3DBC
2ZqyoTr9pH94cXok5Cj4ZjyVgVCr1z2C+lSFKC04rKA6FAVm4qIwa5NNpgd3/iCnXbOKriL4KZua
b3+VOo+mwNE/LjqKGfYEPXTWd+r0xPHVfSiIuFhuQAcpf/j6gj3F8HAwVf9T1K7RkoOizYLaWP7J
gv/xRQ2Iyrs7iFiyrxf7gxrS4txpYeZLGEfsrM0G3cHvUdpWdJy04C6eFzJ+nOqE3q5eXYwTk5rC
AboBHbrndlbGslFUc8OaJG0CzLsA/GvLtnAPerDoWg4gNdTc3+SX5acTNevTIp26K+JtsXvwDHIZ
DoALgBL5LNAXWYBHNDL/QimAM5m+N8wSRM5sIkn/8N0WtWwqQpZDhr9R+cowdq5Itam2yTl4zWiJ
PCJKAfxLtjn9WctwPMxEXYDA21GDKAaQQtyKDqRduJYzwvW0ANEeS8IphLBSQpq6ghNgC1EqE882
lW6JC2M1uF1ulpd5hEIK7RFpmI4d9Nry7AzD+qOnGqvGBA/M9dxnW52ZXw3hFZsEktwmJ/1CF2/x
vuhdCpCWK9mglxs+laJtPMAE5f8OUOPe6QE1aW3+Fmw6XOPfcH18gWApKtqWAraInuBH3QZXjzxn
JtbUSiFp+BvrSLsh8Q6y8gn2fLkof+8da3H64xhhHtRVZwkQDP62PLIAEcuIPRkMV0mCa/SivluJ
DF0ewzRIUga9zO1eNAE/dVx0jPEmUfjOEkfRJT+PUINkIU/EUhHJaZ6nzbis08+zWRlmQvSwQ0sk
YlqVfZCjV0paS2YJikXx1KZICiuT5ByM2+OzCjqD6J3+dbw46OAQhUbmO3KO+/3X+Vjken4oTocZ
5gm3Gi1EkEJ+6gO76MPQZxKplmI/QcqJ/J21+6Q24jb0ENEq7MmIBhCXWXBkxAwVrWsAxa84fYMJ
nSNeJcMovBPfuK2joAu+CHBSv+E05X/tRLf9cmPdPSURkABOGD52dSbbAq4gR8ly7Olv8lJFvW64
eEP+8lO0ICm/TEMyWq4c0Vf4MucWmPRY8uU+jvUQkSJ7GPjjboBBJKRA1e7kK9r+J5swjFLx5Ynp
s12C2dsH4eTe95QNXdJaqcYdh3pBzw1nFwNErJINhhZpryBl0l4FKlP5EzeolB9zj5Vp8a0aWPbb
kdeRG5vIAJi+YhRQxFLke8YCNQOsd93+MwSIPLsrxGx4l5+tlMlRDFDSi1cpxQAD2t0F/6xDCwmE
ILpBdCFSgQJZJKF5ZpUR1vNfUwC/YLhREhB9i3wgrRHH5pst2VfxhFDPKInIvWyjwrzBatMsFWXP
0V1M+bgR8Ygq5X9SvNULyHtL8si139YmaAfp2/ESqf1LZOv5AB8IhYMB30lKDVE9Ys5jss0Ha+dt
gtjfaI49009pY9gk+gkStCmSslyTUwKOGf5Y7aFbqhlHLh4mdXiw7PbJnDtlKKlpt2i57wc8GaLD
hgFEmAYPs0/GRMd2bWOTIMJlop3ALb7D0OBxkEgRX6wFyGQcK/0swQCRvLUxjfhiLjpG3691fbta
hTuq3DoZJ3Rs9lI4klL7ruAZOiebZPTR+oO93Wb9x2Rvwjt2RwIjd6MxHKaHzTUnIjl2FbWlWcSz
cgncqlB49ZRhdUulLzFW1qiPx/QfxscRaDgc/JQgerOsPcyS+RpeeBtY2eO8feiILSoV3skaEe1E
nq2UFFxjPuXdGVGd16Ye4/5VkUvLWaOtlzDOwCbm/0jDqarajOlX4wYcOz4v9fO3STIQ4o0y5XER
fMHAzMJylnUXGf8xpsRh5lAzwe1u9RCSdSuusZkegvdfgYBJ8w08Oph/K2jzhm3JbbgLvQFwm0a8
HCco+G1Ux7oicQcTqK7vsuSWciUYKG3L6cKUoSh+FmtP28L0XaDyvgt//nRKmiu/h7kW8YlOZ8ht
w41NcX48yp5YNBVjddhs9ujT4MQgp5/loNWNQASP1rc6kA+sLZ9ByR3rNRnLoDnOb/xtWqEil65w
zcpaFOX+sKe3nRItY6Ul2fP+IfuBqMzzZztMYAI4mYIQjPpK1nY4qEgZ2nJON0RCy2ZBRLDd46De
D02gEqcog+SSG9MD0AIUH+V1AmHhTxzWNeB2IZ87/1sVbFo+0i5n7GkWwe4PlEcjAP2FVfvqdsKr
LtIrSfF4WR6gM7rQMhJz82idaCycDLRSNIHl1cPo+y3ZuAAqIf4m43mRUhiVlf15OlScoJszd7+t
kYvevmZes6qtJ8D5E5S/d6jlcD3o5ib5An9xgzF2g5V2I5K3N/M479cYmF9igHAkgqDoNynTcPAg
5GG52CMcSagC8DMiX2RqEJFQn7x9SaQhLwVx8Rm9pR0pWVyq2DA3FrLFuvlxlGeSxoEi4n+0Jgdj
BLL1lLfAf8BM77paW8K+xPsl8EFJGrf02oEPbS4DnO/J4ootSAdh5qX70uSkm57qxjWECXVQ5miz
iLb1YSV/Tf5KZrkODeQtGU4QZtkhCGWavsv1JlPNTrBO19ixZ0YbY93orJGX7av8U2MnZPM2q6OS
K8y15v3wIyEfK4ljdEiR3RsufZOEJKkSBzB0FwBak1NZJvbYG0iFcIfkxFpvlmrMXli11by+laq5
oCMaXSL7Zu+5BEMqWdKxMNzPjJtJZbcwyRo2PG7nlw3keZ4FepSwlPVCqYcVNFFRdrHdrDoD/6dp
Z66dttwHVHeL1KSthcJ4xi5F0V4q7NbwYaMY++r0K1QLLJDFiv6yq4pi+uoybosjlTT1aJg0tGP1
I9dYuBynZiUTeXmXAyMJKpph9tMlbBHogwDeiQ0dO60w4up+2czwg5U3/3CT6Ye40ktbIa3WrVkH
G6e4aaqO8tJBVfcf9x2YHxJGLDbf02FewIn0fVHxkb7nRF9nIbjcQExvVGkbh0FHH/jlDlbdtl8K
ahxTs8lIbEA2Xx2nzyne7TSC4i1UuGsMQGEMZXSbs7fcVJtvHLsVtPjuRxjdTdsyVoNvZIpqvIov
iUNN0cHmMnHvTz0n7M5RZ1NYa0Y5SiS+6t8hu4BGX7mc5uWYQHloLBtxscFhOOb0G9eNk7DPhJkU
Th6sD3GtteEBgezJnwXKTxzwB9QJ5ya9EUnehS6wthFFQs9tW1Fb4v8+ZvDC17oIwy3Kdympmtou
pDVGJJBaG1sImwNIX42KAGiIzqEFL1NpMf9pvB/ri4VZwKaS6hoGMGnIB7fdSIAVkBC194L+0zLJ
Pp9+U92H2KQ2H2ijiNRkk1DBRdwerJuui+vud92dObhwnIlyE1FDWndYF/u9njln4NjP7wtiZVgK
xzOakljDC56RTCr1+luz5neknV9pXiLPFRdKknA2N++93Xp3rJi5sUMi4xf0Jpe7WqPH66TE5TJy
oQXHjMjsGdzZxhTyF2qdzojw2kQmXhIjwrsVjL6RsAFt+HIwjZEUlAgzYt4wCl2tcD3QGYYWIbq+
YWL3UhSQuUI1J0M2wLz8WN9GJke8XKEAM9vHKsQ2FrquGza9plG8exZb2TmgB4rYqdVNyQdpA+k8
G3pJcg74Pr81auuaJRm6R8oygA6Pa2QOlTh+jIBL3Y1iWiVPJv8eHPL4t82GQbgwpO+EaqdpyyCj
OlpJg0nk4VkBQY0YFalBksmMOr1rEWI3ZlzHRtnRbL07DUHCbVCPP+Vw1KGEEeUgBZlzckuGBXOh
/Jzq4H0Qt5RyqKPCM23lZLOuMn9kdtphtlNm+lZwYwEkXa9DTiRqNH941jLRhIYthnVEq3ciYb92
K0S22o/NhI3k2zAs2s4letBP4fWYXYcja4Yx2mn7gxuPa1WdRbIASwVfV0lx5dxgOm4GIFzXUFNA
MDtp5YZ/qtFEaaLrg5Ek4ZR69KHieKm+xqB8Wb3qcOs22HboA9msvfegapPU0JcpMuqkGKHWWpSx
/YYJ4xcZJ2jC5raysM6hLfiewaa25bYX8H5YjSET6Mfs9GJbekFfHBgEm4AwsZ12JqMGkAquNq5b
3iLXDk6rHDXDH3IcPQEs5cDdHHf0H0rvkw7d1KsqrE1MTA18GBk6qsummY8+ueFoR64UYrMa/bd3
8tBl03lyT4cAeW5CeH9s/QDqGnmT9jdY0fZJxCKl9lOlnzw3zjO6tJkQuJCs8eeWNqO4UhIK1Hst
YpotGgwF/r3y5VD090ztoQTqa7RJYNJij7T0OcK8YbTJNXlILZL+VIfp1zS64sX03RquhoX9zfdv
Dn6QuusUyea2H9JSS6gpMZaEiav5wJZpb9TvqlOdNQXoJSnsBZdIOXndMoBMT02tPqIHD/GzmDN5
fUUE2bMR5wzTlPojxs7OkB6VRF/lMb2stYvB8G1yTSI+KD0WZDcPySGvU3gpDSIXuGXzLGbuxirF
d2Iij2AhWHXUNYU8tRtlvtdBoAT5QvixFoq5eTkUBdG2hk+L1kM0DDyQ/hVcCQ+MeJAKKhQzHwzV
8k6aYJyv/oJWMLqJiyDj9YYtBmoIjO36YOflGlQel0n/brsQe0myUzdCGIoHTme1eJ28fFGesRLx
8VRGUY/E0v1ShkAmLf+FzdRBdUMjpGaQ5OqtyPuNniUH+f8MphTMV6hKw0zuuL1c69JXIrh/4JGH
LaSkMA/2TcVsfI6Ea7mdijpmPZUMxGMANxwJM1412acrbx+XkST6lLt5gnufELiXHuuu/9PoRYsK
OFQ2CH7s92vebSu/cLdYMV+t2tj0CBQZ7VH50IOjo6g8n+OW1JWm3fy0U+151Zy0Yh+kR0N9NHz+
Pc0aSOzi0bPOdcm4o3Q5QcL9wZIhAq6BMc1XNFuKfTg33PVnlMbSI2DxaE7LqvuCOuxjMyLW0MDR
gVk+ZBifZ7LVAX+3RaToEhAA4s1zcqHKh+G7q9xemckGVuaX0m6VT1BIKcPhE/TS+5utAL/IP8lk
Qq3J+Ew9f2XDZ+rbZVsxYsQH5/yRO4ao/FIW6NdNOt68anWjrPV5woCh9l4V23fKdaMkgJiHGQPN
3fnIqf0ii0ivlGZxH7FNph+hE/BmPSUy0MchUJndftpJ0lCGg+X2g6Uv/GOhJj2RHqlDmhe2Znk9
snI9+IRNnLF4gD665Ec6B84lihphDsUB1ohr5AApyWf+qzHwd34PMVz0G4oL/aunvzR1gh9ltY6P
6N94XV9Hwc/u2vAeAq4o2t+hIycZb3rWX33eOR6zdqL1qvmp/PB19BNxGAXso0cf3t6SAUfpgBtT
E/Ko/5bYoRCtF0aFZ+X5b4rhrOm8DNDojPoJcnIXiPwhmPcJt2F6GzDlJneGBa0yQ0i5++w7UMQc
6Bt73Z/jkb4VcnodrqZhexAQ1zSfJj/DlQ4CcNSQoJdeT92BqqOHOqe3OQmUwBtFyDfbn3FiXZk/
wTyfVYXeAP8cj9mrZ9NT266t5QEv29QkIt/D21QIXaYeLBc9BV+7yJIZWC520yX6oGsU0XeKvf8d
rSagRgTWu14F8za+AB//3rEkyn341RlyLkHgazG6kFvDGtk3pWZjm8czNE1M1RTz8iKa2Myp5oGt
rP/OeCg2DYteJjFj7a6wbFpAcWVlnGJ0q/zQohF7pHHT6gs2vNWr9jbWMPZnsTW840adjbP/DCXW
nzJXH8EZEZkW2QohbnhlHFdMdBr9SOYMYyRUfoEFrzR4K6HSvHlN/21vcVEZcPlVH6CzsPiSTP8g
5qpSrdQ5GE4NjTLeFvk7a0N8ex0JK8RZtjwbO24K61zHNbCvNU5WtuOystk+f0F1TW0CFkBAe++c
OEmsmuJP5/zB+z/5wVk2BpiKc8zVfU7MwtFckpCMpTe0LruqAPFHwEOV5xs/CZqcVsMQB9zEiliD
8Q6+XgogGf/tSzjAr2ssFOzLSPyYyFpCWhvIhjfO09WDyUOrRtjOJCg8n1YDD4Ir8qGOTojwUPaU
B8a9gLFko4ULd9K9uikfmY10/os4Rhr4YUQ/wyTfZL3qyHH7ZrNjZbHSlIqmuBT3J6RK0lh0kFz3
GE0wXKGzAz8nhI/6e71d76h/DEvMeVXIk0vPutDS2h5KT0Q1fBG9q+OUHnXu+fFKnE8ML5FGPQOP
HNzhrIoLzkQZson4WlD3qcBV8iRiHkYugJa0LnJIgyS4VptFDc5f0h2kOcyD2C90xxH0gHfQRAVA
/rBnlHpJ+vsuZZTp+jyfuKLC+NSpb/hMEt4rEsSbbzCi5BR2BU6RuRw/lz4fCtxBfooW1HQKIxN+
/XD5aKMPy496qLuwg6M5/furIFkyvFL8fmiS8UuQXTcuXGoVHL9nff4cBxWPa3mLaoujnoya6hAL
HG7RYhq9tnwxFLvnU42lrgEf9YMf/85KdgjU46oEJrfoEOvF8eMCB4vp6SFtSaI2HjJNBVTtSq8M
waq+XFOiANQBcw7RPtCnzCkTq+WmdOGJrr8OOeNnlsCcxxpWuttEWlb8kqSEItAgqOa4KXJpXjz2
n94qmX8NtfmrIwTrT5rMpzFpBlTTcrt8SqpQzWqUsGerOuRSIobsD3gnxaSeWQ+ricqCKUvCG/DF
nEvQOVtc39uQH2OuZNTa5aaKG5AHr5hOskuUAesSXr9MGzkh7tdxhXq9OVScEAWCcrQ/2ivv/ZoJ
u45Mn9VPbeKzuQgdi0uJw3a1fb+vW3NHAGt7cfn3RHMwoodEU3bqfqL0bOQ5gnJ0ArYKhJ/TZ6Y0
EbF98VZAX2hWV0z37JsTUrbP6ovZaOnxFjSV3UdmTzGnZyBBZBPdDmug4Zfv1Gk05sxze+O9526E
MYDdtgbXdZED1wkSveMigGsfCVlGnOObMFwMpsS89tBrM35IYj8guhXFrjK6HXlEp82l0YTV69Qy
U+74QhzH3O4jzLtwidCU1ZUqii7ZUwIYZ/UnEV0tOfwtQ22xAGCFVnHv1P64TSX61F7Nfzzfq+rN
uJs5fHjU/8KwOOlwUITQ0qQL2xuAzlhJHxn3WdXU32gzsjuyATbMxAr5F5QHB0QBUvyFubhiChQ+
83jQI3K4dOGPuuU+CYNihQqP0KDYnO5yuHjCZ+TtzszFWYJfIdk3nLiFRNNqamfIz/J+vAz3SDyH
64Yajdg8W0EC1IgBnE0U8U7mcXXenzSPsA0TNFHqi+IR9Iy9A7UmBuQCKqjG7YTIipPMHQqLOmz3
GRO1tpNzem5Qiu22xTtWQB5MyXPsW1zSGkjMCJFaejXEVVHJZcMhUhm3YRgjopD3K17RTshdD/xM
YGTXVSnkynZE+dkG8fcQZdqXh8IToqtRiBV3ihIddp81mKAUTeXmFIbk4QrIRXaIqBpnkutWBbqO
TV16O/TOPUqh1353hCmqhjgTW1CxBNbLmZGQKk/4u2irOglpapEd+fmGyBVF7p906UcbTXI3smsN
QV+WvdJ1meMwBxXj/alBeSZ7FmXZHuLOEaV3MmFHWAbEYV2iWWEsjddYw5Ao6/1b+bZYBQ7Juw/m
b4O68/gFukr2sXgFlAa7XZIxl+28AcfkmmA9gU7OEjXZRJ2kyGOwCE/E5TTOYMwKJYNarD+LM9rU
Od8gW+d+GMFD9D98Is729lPYsUBXlazJFztgwyOE3GQ4Y0w+mIlx41pB6m8l4Ag/F+wf1V6Ti16S
He+WVbOzgdUnbxnDR+O5Xd5QVcF7dD+0MG+KYaP5A12M1HHIYQI00uAMptK43V6ZzwfYuc7DW5j5
8Yu2vm/kmlABSPIKkfjpXUGZxTvTwnAc/2TAQoKMoJfuD0h9R2puxc17I+GecPafYw/KCu6aE3p6
KqncTC3mmPmV3vc5xf/sSuQyWOSpLgbCvkB/xT4UPun3sUgVNyo7p0SnljamqZ0dnjWhAcT/PKZq
b1ns8zV22OdRephe1T9fsJ4wJPAZdInAM8Pghw5KoWopJNQ1zA8DewUxinf+tMfRg21A/rRWH8dq
nJfU/boN1QWbKTo6FTypBHFafzkeWyqwfcDN7sPNuz5F2zX5K0rdS8ZjDcdxPNR2i442/yy90ZpD
riRaq2XSIPmhfeKZu3fCJn4LdgB8BoE8XgGFrct0zZfx5kWszuuPS1X6958jY0nc8oB18QRguVTz
32Tgp+l5IpfIlOzqEmNM/eFFGcX9QnWDBJyF98laIwxqx46uO/GRyD9jNwpsj8rNQrLaSxuU1oTP
tKEczjCZP5vTzR/pRpIlRtgzGX7SZIV825Hnzeb18TzacbHz8nFGBbiC9Jv3AD+YReprqvAUIdah
yyhQCEDMPIILl5Y7DGNjTApywYiHJJmoHoJ1f7A409fIIbxgas5EwBN/7LeGEBgWl+1X5ARuEmNO
hWkwmjLpE4LE4QEjLE9msVuFrjI6QwsFOGhxCVc3sJG/adqi7B6LDQe0e0bvXWzqxFmwUuzCM/xK
RGLQ1Fs0BN2PnqW9thSEjRbuNAywghGoifj8ltywYktMmdJv9qFLgaRqrXQ5RSe1L3t8jyI7oWpc
yqG09CD3XUrVa3/JZNUAfnhR9XGazyNYDTUfJNZXf/yjtq9J8UZsZ1B5pZmsZTEvJK8wveNkc8Jw
0hpa74ouVCduWZUaMp5mgGK9TNL9XWOMA/fuPyo3s8BfuZUVHSDrm9Wkp2AWCB2mk5Di61ZN4uTf
Q9Hx9e1enCpVVWuhK+1XvUjTuW27+FYx4yRMptKViawd7v60V/AVtDpK0ZDno1xcfO4DgR0J2Srb
mgZe4+HyW9Vl4U2VTvi0MhTdQfbFwqdYk46haKS7kHCeGt4j0vjyIdTINBt2B5sTOZ9JqyPYGVMG
tWz4+oQ2HtJQPdINBe+jH3bVEBbZ7vIQN/maNCl1SzluxYqN1uza8fwlODG2VeAiWVkuEsDtO7qc
nW0/vxRIdcuQHG6HShy2kq2AAF+okXRHnV2buIKrIhVKCCkkoAWYqE3x/XG9VAYE4YlA73OBM8FE
e5LNdX6MD4iA4Eg2+B/dL2N706jwmKYky4MiB/Su1bz/qlg2P72GmWaydGRc3WHnGHG2hkjg1F3D
mhzXa9+7YgJNCcDDoWo2+2OpC3c4l2HFlgyKtWQ8SDVNNAb+sPhS+JDbwDZk1LzLMIPbn0DutV5F
F0i4SDQfAENp/sowsRGJjQX9yN8col/ZSugT/ToRaXtNDRoA3wHPal1YwhCqsFfZDkildzb/j8lV
G5udm6HH78qX/sooOiskPBiTlXqtC4UMaPrrO/jgSNfjjSqzRVdgDzVdIVop5kh6/YqH7PPQAHGS
K/BM8dVPCMnxHxtxnkDEeywSRjkVZ4EMJchejnvuLjsmbQPLgqxZkUe2LLRqvmnmWhahB9+FRthu
SR/sNcUVtYSWmMLX1k/VMHbNDJdqEOn4QQNJLAQ7UOjLZmhaKD939SRBrRzBKGCD1pyopt3/uedN
ECKMJfWsW7y4Bwaq4h6glW3FN5FelyHrDYcMhO0IZj9UZPbiLvxCy/zUd+8psnEnsavzD83KH/gS
pKOpGGrNntlHVZijtoxooBUksFtFsD8/4RMxH7mbqzAYzWqlQ6zlk1PsEhe5/8+b6Z1rx9U0aq59
l1Th+XmKOr4G1UpSROO3tyt+k54YtvwF0bRZWizXIGOv6WjFFBw2n81+xLpzYc8PI6NsDRtV44kO
nZw6MRvN3mz4DeHbp6UkN/HPh2iPhIpPrKSArcapekF6nMcaypSgyYij2SIiqR2nckoq7HBQBiUG
bHexiwsvbkrfUO98XW9CBUSN3zXJm72xlDcj1wXQP+g5+Rb9ZKoOpU9snHXk+PEOTk9Q7WTDKVxB
a3RIccgvaoyjVrIIKiHhs5PobvEPGXK+zqsL5Wr4IkXVOdYoQnCFCts0SJ5vlSEVScPZiJmlRf89
gRR+JkoUoB2vGYacUp0onBlJnXi4BDbvfKAiDzsWSmlinbk3qPBo1cXwjR+F9WwhIBpZe8O+zOrx
9JvDpeoU9C1XTNIxAg4nS8VU1hGTZJwIb8nPrNxtoCKj0/MZ9XSIVORU2AMitpispi6QNIDt6Nam
Z8j7qZzaAiohqD/Y+8S/73ydBbMR3q8PFpp9qjeF1c7SWNtm7mJ2wHGoZS0zfWDR2sJvQGzHgmYL
fm4/dJu35XRupHpofIC19F/17JgQDx9CEvSC5ImcFtxqAHawrYya70Vd8xICIqN6tI2L6BWIADS1
2ywBXrwOti3EWyBi/sIHhQmSv45pNYxGQj8B2M9Te3PvmN+31GMD18Ku/KrGqRSHMJH0NhJqPBE8
t+jDmRqXJGe0EkPY16EgFftU62sEH1DxL3DTGpe9Y4MdOzFJgcm6CIfgUoD99+g9tZ4GUZHsYc07
t9HXgx+8Mb28re0vkzOMXIk3OAucGEGRXLXuavowTpRij7goc1Hndd/mkSYHaPpEk7vvJ4M/h1j1
IUk7G0Dj5eFrFjJltSNsGhQCR0IYEjQmvYOaf96Zd9nMYtJCWnibRKrwHoQGoE1DWOW08iOzXL/W
ZBndhQeIW+zeWS9yscyYAz5CXvhO7id2zOsQOrJuN8NqfU0DlDoHcdABeiTLd1HJ60HzOiLr+EHZ
9i6oLrifeoNVM7RHaP9qsJ+5ZrrFRrO2zQZzo00gNt1n4oSkv9UNZX0e3qWNVWLoKQjM9+Okxggr
3B9ctZRC/2O4hk8q5NcCg2Qqtq0xE8GZeDOu6xF2WRXSR1dqVXjgYVwp+JPs0fQpUd4ozA101Vcd
G5+HrJJMd3xvobTf5c131oIBZvCdByLdke4bkzJlHe7eYzWyxC7aYz6xjaT8amr3Wy3+kqtcCy1O
waNNvqKAg4tocOFmTblI1kfrkzldDX/dpanYD2VOcO+WMv3pvA8UEzJ4FXjdb6a/GodY1HNw29Sz
/eomfyyYAcmeuthWDHaMtyphCqiqMPrtcFEf9C3IHjzwxyr4aVJqN6oHkNJaMAqBf3uSMvz292Jz
ORcQAyy2epdHtkXS6wLCI6Z7pOkbMN6doxTXNyCyKTPJoILZFaahrrCPBLOCCRCLaZ2W3X0ZkK6/
SEC4XjpWWNrsdrEgmGHuMyFRy2Wr2I4aT0s4xfBa+KZ4YgSA3O3JZhnn2y1cVxI1JR0Lkw4Zn7Z5
uT2jqJBJvlGQuG/gI8tuNMsjzOjOORKQ/JMz4Wxg7RA+h/ncQlWPyJ7ns2puJ/e0GtznemF2t0KL
ZNS+RVglMfN+hJFijrbvjouHvXv/0/ScAXp3QckKjlAAw//33xQJKhOHrTrM61TmH5bYpWojaFF1
qm6pkdS66Yf3MxG0ZrLCBi+tat2NHXLXAilt3JRdcVfDuZkNdmZrOtySReuh/1bazRSezrSVv9et
jS+Nh8bL42XF2kjRbsuTl8qPEHQDAJWl+LMgoLxhQ1y/4D/qf4UQsvWRds+y6yay1gMS8oHS6izH
zeaogAgdLaYsFZrDHFIyt72Lad0AscuY1KL29OQSNuNWH/5cpBa3sGJKtTuKN378jhCaP9TcBYn9
vF5t8RQXN+JttInzOSYYnApMVr6+TKE4CmKeIR47XMVZjco71CsVZeHdjwk5lqmrhoZuzcbaFSVn
1esSRsObz7eW+vTYISNRYfBIdRQ5Wdd2/sj8kMVb8qEuut4+/GXG7g3Rsr/rLLjVWstxfdYOwrN1
3VCZ0rmxSDMf5vFJaQmI5CARO/HH1SnvWTciuNgTiBcRmgD1kXz404zMdmJvHIwmft6JIzXG/kXV
apmADZicalAnzZ7EbgbzIa0YczM0eK9rhtlcKmT5TKFyWl31PB+7RdZksrxvCw0/vQIApjuXn+jX
F5n+nYlkXeX38mZs6a7xHWnEAKHSQH6V9dSOpXJQ4Epz9B+s9fp8IqhUN+fX+5PSO2hT8U2eAc0h
oFwiSO1d1+blYevhz6MrLPsAxz+lsAlM2/0zA3yQ450XD5hzoeOumtd1u4Opk3Z+xxeNjhIAw0Tt
YdjUzBSYuAiAnHvXgq2Qh+qzT6vL/CM9Tjw/eo2bh/OyJSjej8eInSLfl/sAxZirkLA8WB80VWJ9
P89RpkA9VGyR1wPbQVv7QCxhOE3zu7gtmOCuDQRgaznE9OnVbUMPHa/Zz7+qAhFfGsMzFolF5hzt
SZX4PeAuKRrTJnbGU+aRbRIeLzu7HlR1799AvyD5kE46gwg4D9gUPGiD0hXgYl3IJxiQJWvaCBBo
OwB4nwe1FjIMqTPW6WnoxopCdl62hcZGyZdY1xrt0bSv4NC+VAFYNYqh9L2OoADj5QaJ/4polquv
VJ2H2081o4xOldDL7NVXgfGL1pvBGhKX7DxIq9rfHauOPnESAQf8BBIU9ERu+63c+rG3uayrYBrL
H46BrORCJIyuEZ/PJvJrgcRAscQ7MkxjCEJpTJkLFmgqrHR5CBcwFyLKrfLriqVW7TrQzC3QiHx9
CecTTN7kA3m9EGbzgL31eU/WHCKJEU2SMJyULqlBBKz2KTAZ6mfRsWFp9LmLtFzFjfI1kViJaQQq
3lj6m+2NNucxYt5NoHEY1zECF448gtZwybX+yd3Jh+eSJqApztFtUc5zryA6QV39hWcjthS0h/Sq
goETPNKX6frojIidS5vqPR0Nog5nW1FTNzcnJ2M7f/QtB+TQg+zOr4mutDqRa7ZmNsyzV0TwS8xn
aDRtGxqkkNdHR7Chrg8arH8TRNdpW1mxYPJF58c57LZkJac3sltVhzEDUxMtu2BVdMl/YRPkrKlZ
mpTFgMxsl7YirMb+VF4m3MtSFrOQktSUA+iX3NlNl6ywII6JDMJZocOWdQGASUL/cfSilljaEnRi
YRsLLjgUJIqRMpg6nJ6HCYuwt3+UNTeBIZqcpSUJHnTHoqv1hSIpqj0mJaetmAId+3erHxEzcXba
c9EBlly3n6kOliRNZdytldp1HMcNEXpffMJiWn0xlJKe4qnV5aY/HG6ZbPtA7A/M6AvibhFfvbs2
Y276BV3wmf9S92HkoS2sbSuVJpiZiqRoalL0WafJxxxSzHXgPbBlkJ5Ce3t/QGFyHwBOSqAZPKsb
lDDX5fwA/VRuC/yMkFKq1dfv3yl9v0CChqINOwfadhBOXlCW7nUTWOREDBfC7HbidpR4plSewCj1
LccX9UAbQ2EyIC230XuSWLmNsJV1BZg94MugwVu6uSH2lrqlMX8E/jhlJcXFRhphFOaCq2ZyHx6v
QwKxfkIduHUCwproYOq2RmW1yyyY9wyxn7o41qtx+m7rgWjBeKfr8U9IlZx7K1VSCHSqwDmDRpn0
qeOd+GT9I0z1zbTT3oRU1kGkTwWWR8hHCuqbYNDWBKichnDrKF/PhbRQ/U63p6+muqespAgFFKKB
2w8yZd9oE+be3tHbCGwXuFWLqJfMcUeCwsBVzKNwSyXbFzc6X++MWQ+bJi3YmFBnFqo62tx9Ua5U
6lGW6DtgHgirC3g9QO//TyKYryPXaBeUCY76sRwgClo+9qrEOEP84hpGOUUx21AgWKX70q0mwbwX
Uaa2eYFIglUWOsBlGhv0hzIWUAXyVomWXsi4+QeFn+wntDoQuK1bKZB5H0wejrnVUEyCK4wleMpu
JdJ5WUtgAe9pSBMHG0beHJSjxilglQgvcMThBxRYEval+RvqwtqkQgXodq3dyWaAYyKiP4/q23Y0
8dX3i/SAUuX+HHc6u7dk1QWcQgrTOpofpW397HMUyfLEh2hOnlQCeLzScdyjvs63oYaI/21FQ6dC
0qJphk81Hfi9N8NJUmAmnUVPcxYHRP3kPJjHUMIw0R1TRnPQN/7Sm2naAyrJST8rJgOtNXfg3p2Z
c7fvI9G7MreiHF5bXH0qYFB8mxEyZPQsw3Of0MnnwVrJTFgNcvxVklRlY+hup/QGr/EgtMeuq8P6
cS/eNfYQMBBaBJqKksS12+U2UYG56c1hYk+5ADtPgsKqgfTqvOVcZDbmOptuqo0gnGPwW5g5ucME
ZtFGRrx831wS5daAJmOtsysOBKe83I7MMt2FFCjH0os3BvVD6YCVJJ4SAURMGTCg7q4xFfQf3yle
BuG+Jci2vsvFp0/jkYW8eD1qv+2/7KsoxZdfGxftSHTiw7laLlCfSAAbEyjh6cGHpVfV3Wd6HCHY
xmsXjW7hevLxMV3Ep8TDoS4lrMkeydS5EHODXFwaALl/ZbqLra6EEf3th0p30UBiDTDssCL4B1sU
WRkYKbV6YX4wfBnSfxRV2ryBu3U9PBFIcp4MqJSZNvrZ4e25xRzAFu7pnyNkCMg2noRUxAhMce2W
5ZycAB3gNzzFgul0G5o+UKxpAymzUerySKEGpdxz4OLaCGl3A/bh7BLgmGeYbrKAPun1M5Qxs/6U
D1Fbauj39VbZzQZ1KlvanzfHI9+JlBPyX/0RW6yauAdtgcqu2V5WOMpISzWMyh/6MavSJobfhmhq
kRulJGCOBTq2kU3pqNY9jkAzyZSwkyPBXYPuepPJ+JqqCVRf/eIvFIEQV0zVGE8UtabaGjLNkGku
AdH7eDFjXNE49C4Svuoq0VQkRDS4FVfPjVHa4xHmsnjPT1AlNq1ZH3A8uVmN693RgUTDMo9apX7D
1S1S1h/DbUZ4ZTwL+ZudMArRbx9YnVbFgAm5u82wxNGI7EKrn6BCXZ+mnGHHlbBXA3GB0S1/12N3
nVRtpBXEkbTqfB6WL9OYBm3xk3WgWwIBCbj1dUWzrdOqyNLPYtMNVq7dNmK9CY6d52Me3WbBjeVj
P00i1Hx4FvfY7zzIDKwfMwY+FQL/hFYQ6StWWNu2WpLPVCibnU5P2h5fzCtVuGipdohNnEdjJg5N
1KReqLr5QV60hebDcAotegacpOCVdNxBMgWFfyT7KBxbhLuACdzCfLa7nguuyMxeCPdMPnjoXomJ
kOM0mpHJR+C0cxOEFvmH7pxiTy8S6DHAcYq95Ais0BI4njr5HGm8rioY8mPn3lIgo4GAWCnq4hiW
TB8wVlSkmLVbujcjpo5fA+MZSlBslAkFyl/Qmd/cmHwUDamnx6e2s0Rhbt9UYc1qE298pzJz/Q6z
YM25pqoM2dWZYtYleZFe8Ilil8osLjdwJ9N4JpKTpykjEAIikE4LbaAzoeKuVENyD1ERVfoDxuqB
iTuEifz0jCVRPrAn8qtMwg9RRXFViDSK2pbF7NAyzw+zoQBHqjFfejvEZa2Kgwq5CJhvRros0S4E
4lc9rYKuV1XgxtUzhLzOWc1SfQMRYvE2f59ZgF4y2ggTsnGeCJzJyNldpwzmu6pavOgTKUcXI55I
WLd+ztdaZCUwO2TgDOdTkmrdroH2BI35lpRQSm7UJSd3rtso7M659Ak0lgx//xddK15L2rtdupmt
ZSc4qK7sZTJsNPyxcYJpxPoEDMk82qSN5o/Fyy4MlpT8tkK5pip/eP/uAgmVTUCC0MpSxJHNBtBv
WssQkOHjMvxWxOl6ZDudoL52XXCgsV4jRWWg8MPC1zZUR31LgXG8N+4MXlz227QWbvEz4RmIq+b1
qrkHEDx7i/zJH9d8kROkuaeuu0l0CiaMt0uuTHlCphf/DyhQKWEZTT7ONjrR1GyONw0eBs46W5fV
ualWUOEHKJxStwwkHJVL7e5h3cvrAcB4Y6kXLDYX4mIKJ4aGNsDArnM9WKQJHx8Jg77Li4YBinvF
/05s7Yla+yzCakHhuc87hnnOjMkfZlBhvYDaUrhy8yka8Ap8xcDqBDj6SBOtv7EolWoCcm6GRAcn
H1WNa/wug+0g4pEkmCC5GW/3e6gze1rbaeGXhFA2eaWew1Gm4XjafFVl1Jq+F6tevjPmETleEuXf
gWlOt6nJZKSG8YA08A4DS5Lr74AvE18XJLgiBtnno8PrMVDpcp7Dx5x3uaqP0LAJ0xdDvqIRdkcG
7WoWKVz0ylGAZ+QxISWIxnn3fyiRMooCk56F7TQXUCsUhVh1WLas3xeINtT7jyn6vcl3bL8OGvMI
hxzZb/C9m+0SoSySH3vjIkH2cC2Dkgbh8sLL2aJWQYS+PDgz5KQwRyI4Z+BUiuyda+xjai495Stx
BY8sKWQArydCkNOe8LATCsUc30P0cO40qlM/5IIwrMDQmvKmxmsIL6RVjAUMH2jpsD76EHaeB6kB
xG9xCHQjOluBjxq2DswqIfAXDXQw46lQ7QumKgtc2XNxKzAAdZJ4Gq/5OzAA4l7d2xOFLVBLvFmv
cs6Qon1msk8jBqtPfPbudBTcZa032qz3u8aR4QTBBXnYgWkGFBf5qUriT0MV0CxCn4lqSW+rAKm+
1BAeMvUNoCyoZ3Vk8VPPKr+94s7yrHKTD+0IFGFQg9xOjQGEFA4tBfxxPjjkvEm7M9XpA82/I35i
Ep3ao/0QLUWI++jGLhsdp2sIbqw5M0YSp7BxaFBY2sJfv4AOgrtnJjdUwJ4zXqD2x62Z3W+X3pIr
GUeqsnvrAYI7Qw0H+5FjhrIG4t5UmC3G7GD+w86fjN6w5ETJyKrvWXF42kzPJFo9ubtku2C/bWhX
CGI5jv9wRXr08SeaSP0+oS7et1a28ffICy9KGekRHda0rUeSVEaX3RnuPJziDiUL3QwKXCFXzmpk
p/FLZ2npd9hPtN8r2ILBaCfx/Swrgm+2CSTrbH2BRwKg8aSZDtry5+4xev1WpoT1PGTzR/1CLpWv
hN1IqzfU+CnzPiFBCYgmnv55h0UBZaIGoGDyBBdl1mKuZec+pWVFJzH9UN5o1pveZ5YAsxDnsVYM
YACwPvFpev4t2wlY8UXyABwimUdRtx1UMaQLZQU0fI0vxDOltYKsE/dd8UFxyTviEYZPYCeIWQZ5
kyWd8ZJMJvonGFd6vhpJCu1TI/j6T3taprtI9eDXNfj+7FF3pMqQcm+lht3xMFAtLk41H5hXaVkl
wSiXDNF/uxixWcKCRr6ppCXZQO6t21StQsLAfcKWIFphs0+3Dz3RQ/aikxloEASCCR+d/A6YkYUE
EV+eQ2kJfs0FXQp06zwCBNT6n5OS2/gyHZoDPJpo42UiLDkQgMDrsEvkSQTkiKcWJcWSkyRYYMpv
j+f1E5BYlm6OgWYqmDfzTOy0QNHUPFbaTnT5U9iHXGVN7+ctdlraJHJMlH+j5ihQC/VtlSXk1RdX
qxUoOsj/VmPYnIaVWs897hUhxV5yrzyWRFn20l6ujCylrpkgtbz3Q2MNb7f6igLu11kBw4u7HF2j
aeePqmn1rd5egvHh/3sH+mNF111YBoeUJpRb0jzL0oGAkzP6nccksZkwT5EJeHdIpu1FVKitWV/I
B7+r9s1ILtg96ZhnbgajvW+E+ty0ltdRV0NXq/kwWKvjPKbWQr0+6tVgKHtdxKM14OeHg9IOEDEU
qe7g63+h97H/vLybpg+uYywL1EH90Yx+wj8z3aFdWlRECLon5IhGXsSmTzYwUfePDPvLiM1plE3Q
nQymvKwWXXamyPSQkZd2F12+2lp+ekkj5hkgqU37kbW+aEPzPJcN5Uuac3uiok7i/WIdos/8VERb
U+UD7Kap1bsogWTvX+EzujrGKmeYDWWzyZTpsfQNXQBDw4n4zKH9ljsl2DE1XAn5AL+E8RkaafEL
PvKg7okZZB5PM0UcYii7kHyEb3iQBZkK7auy4lJDEyIhi0kdifLnJner6G/dE0HGemMPJ1mw/+vX
vAa60LCuScAH1WwZTEELINZ7/Mz+JWidH7Kg1qVvN/0ZYda71z4j6TfD8kjek/Q8gHRdU7jGPp1F
wB1D9NZCWcRJbHPxJNzH6inFwegGWqr/FXvbGnT+rAH9GTdcJssM6zPMkXVN6q2Ofbr6uZ7VaIl4
Tc1H40fvjYxtztZiEHGUUaRp0QidOzOY3lI30H1ldx4zeZnHazbYbyQddMaDekAbFmly4+AGDfYB
WCmeWH/JyHRKey1Qo/Trj4twMMdriwFcAx1ZbrumAeweSjDbwozV3991KpThxQXMX8bK1LeVH932
L+zOUaYVzrShsXjIdZBB6K3eyP2SuFs2sx+RzUKFuq/MvTZR8CoVc3zJi5KyX/xlGTnNhvruu2kN
eb+Ed6YlCd9T/UVrmSqhV+IgQR2JkXkPN/IvOWSUdqhm5bs+JiHEj7A6RBYFITuGjvCCAgO/ELib
pi+WwC8k14WDsZ+sli0o4wHwy2/Q8nB2+AWGc28oo6w3kjOysXh5T4u+iqtL6eXQCPyioQ7LCfUz
DH/2jLnI6jNuWmd0nLvm5aYaZofjldbH1hlvOR/pgF3wwKI/ASaov6LXxYoQJ2+Ha6Illkwo9jSG
xAThl9UwG5nT0N8d0k7d7Ffc91UIi/rl5RhEU1WGVSmdr7IRMbeQq4H1y1fttEEBO3AOMpX8m/Ho
diiDu6Pju1aWErAyHPI7ReK56xMmIT0mRIla9ov0q/U2PegKWSL8nj+dMepuQ/iYbBCcu692XTgB
iiJ3yJDv8GxVzTTlmLnJAM6BOz+ozXhn8OK5KujIEQIpjBKILMxu4/P+K2uKdAQDm6yFzr4fBhr+
FTMXfuqyzTua/WKEQttrgrgGG8p9/c+v4XCjM5awfCqubjDkloT78mx7COow6Fro6oVvc+CLQgVv
oxBotJ3kfudsMtc35RHiX/wdhDSVrP5ALnJWFRVnz79lq/N+i9mTaUSRSr96/Ic2FNB9mPktWPOn
0XsRy3aUu3lAEFMBGCaMSTVwqvuCrRevpk0yk9dXRDT1Y3xXEL9kW5sUzFz1PL5hoPhV3akd8EL5
O8gTnnMy+V91omS6dYMAnNpJCaEnWG57sdWDIROmGlWajOinSmxmHT5rNdA8p7nxQAysBUGn2rOO
oNkNdCNABTwyRYpfRhtWiR2y9Zks4qPVYMUdxXRBpCI5iLGZTw0MV7PRRj91TmTv9t5hYRLUbzmo
Ap/OacLSm0kCVtAsAmrN/iLxCjgTKS5nwOyry3nF3Lym0pp7zXAjD0LZsEYKf3hl9cF9VXTsM223
ZqXdK/z3deGXmYgg8DUEc620D+4mRyTv+qzPNKMHHghDqSVi6EUXA+4aWIDjQZ2dp0/dqQUVZ0Up
pg+kC89z5Z+K3tUesw2dgHAORH25tp0jo2jFU2/WEqSq74Bhahx9JxKDvorwvno29ptoL08NbylO
vPCKXQB5cyI1C5h4/cYGaZRGyy/3kfqKJyOnxSh3JZyTK0DKeomZmMPetEAW0pbO5sf8jXDuNvmx
hyJyriJbGyud6xgFhn/CSeD7ZvLIzkZppRHGGYJ2aSL4TVSCbIOU7viWxbVvFbtff2namsc9HnAF
zMdpM2mddoDnKbvSwOc5750fAPVbyKrMtAELCC+tGv3hTslh+nvJRVLtq1H80zfitpD+9L/iiOif
qJb8RCVFjlgCegmJ3dri8m32ZqP77riCgBNGIb2yvYgMnOMGKec6Ztkz9Qx6oZGwwP4MaKUL7S9M
rOd1/ymT9gX5PRyKcybPVLWRMmHv3nAetEpH1dqgyw1kF2poiRu+/bB0Ql1RTD+HIn67JBNqBWD4
Ga7MiDlzZKmLkzzf/ELQsDnKp5L23IQGKbS8qSXEP5SyCqXEVHzc5CvIVnTYuCIoVxRzi8jLDv0N
3jkVUrM24WqLD+eZT64sGxASWdSgzMhm4H4JP9wOZgFDDJR8qdOUlgRyJnsxfc4zr1inQnZo0lyy
3ck9J0F3Y5QDchLX7h2GZSFY9IV8CJvjET4CjqjIvOV11OXIvopsXtXRUN1po4CFFLgYzJtJp+St
bDgNnQy/n4ksPkkRikntQNSz4FaCvnMEjp/EeEICZ/GHNWRN1Szz4ohbkdAxhnqiGOX29bh9uK2d
+1N8TkzBNR8H+M6igghLo6z2XzVnAzX/OqSC40WwGhpVkbJ6hIOP68SFTT8l+hvXlFvahU/ytUir
ZBC0biV45asdggW3rWN63IVNijOZdQd+bb/ivwD2tVZwotJrKEuvTTs0bws8Sm3LnEMz1m9Y727W
IhEkrR5RMnfZeCx0AT62vssKR6FrpKPsOHmNp1+CD5F/XJt03U4ZFKSJY+iOlUvuNfWn5Tvbf95H
4+7C04MWgyw5aDIr32vGwXYgOooWlxskQ7EYJvkW/1J5Qs3gikN2rpVCAjpMMmn9HgdhWejShvut
106E4QTpjB8XpIZWWaQNXTFrqsprOZVCynzrClC2W3U6/88XeV7tzTI69V56HFz7v0qf4Gl2bNwm
sSdT+Wfzw9f0FAg2D+kUSHKDQDoBEpyTfKXcj/7QjokEUGyBmMTF79XKAGYtbpxQDxdC22mPQ4+8
v2i4nf+LA4wKwOzlYiuNZxy6+Bp99SP3crpqtykFw9FPrEMGhb+nqHNbEj6z0kA0h3mNKBQqWVFh
J7vOOUQzxEhp4AUmX7YsPJxYFFYTsE70BJBwVDAAG20CndW3URHvWsi+Hd/9WcCbi4uZT0gblP8W
TB26+8MwYxq7NO25fFrvcn68IZZv8FmNSHGS6ODqcQv/6a8lsvjkuNEbchA6uKi0kyYHU2+QiKgX
vMZKAERiHpgcYAQISdVON+Sd+uxpVeXYENYWKjtGRp+qywkngrYlhfkJiL3HzoVC0zbI1txnA6Gz
Ii4wy3l92c2cAJogb4e898GyuZJ2X/aZq48VR1gbcO++9GlJA9q5iMAY1BfAVS5G4gLP3HKAs5zJ
w1BLrdktw5BHcBW1KAVbTk5uF1sIhViRkHf6aqwd6pfoys92w1smPJcpgNzrhNaxxH/nTR78jsOO
9oMzN1du6RpQ5ZbCsb6x9oRtWlJieePx6SJZ5v9u0p3dbGh26OVnZzVDlrhtibKcre8vmlNCylnp
9QqN8g/FGrxDRFGGyty2DYPgz+/vbz1fXUVW26++PkPbKObRF/sgr5XQt8DUpglmsVi5NOE94Bxh
DDS0ON7ajTMOJf3Zvxn+NiRuh1ZAQv/KW9Iq0OEO/NlFiasE1J4/9kebzVU1ZGRr4N7MubjL/Dlj
CJsFC71vrfJfuT1jlKL4CMpzVii2uyoUSf7UIdNc/5eXYvnqJ1eG5Bz1dRcw77hkyp7jTwwePaYZ
oBlXFekXgWmva8krA9aF9O7NyeB5mNUYU000gr6ox03LziibKOaVTxszZT5gY7/yFouIhc7ktVgb
YskVU/r7xTctls2vPxCO0fRA9co0GelTXuVonJTgF31tlxA4jWerXe+0b85rvMf2zAS7yOuMmFh6
cUEjfok03P+1a3irpOCh2NPnopNPthQdN5M68TKQjV6F0ivo5sHVtF+EPXqyW5MLcgfI8cxhVmiD
GYtFaFyL1t2FoMrjmKY87mtRmNthQn3ND0uB85UEnzaqsLDhv18ptX/sAKsrqgOHBw7BCbR8zpFE
klMzLm8U7qqAr3YSi4FR0hhXZtnpwg+HBEzYM9ypN+/BiXlKADeSRy6JEdOB+MBxPiecxD0Zeaz/
t38DoSgrI1JLUP2HbX7EDxlImNNBv2neiAOjh17UU9TxrHbnIxZ+ZkThGI69B2RfnR80nD0T7M78
7oly1uS4MUoEfWYIHyl9Hua0JuXQ7n9wImnDnlEprm6gToIx18PB+g71LIs9Ptb2C0ClasGvHAKi
NMm0aGMH1P+4W2SjqVY0xv8vr1rGHp7EdsAOaBA/jpjNf8H23KCbGc+T433JOM8euMfPCbA1BHFl
5kWRzR2uag+j3dP6CtMsOZZU9cpb0LFtXXXYsR2plDlZnm0SvLAKl5YIsC3IDfjE5Tg4wLArdrPa
MCAysfe+Mq5HIgCkymfZon+pNSYrGuFzuMfrYchJrwuZkNIYAbVZVr+sx0elk0wx7oh89ER82H3Q
ehPT0mtDjUw/bYOhh42yU4Xe3o4OY4PXpFlHdSJuDh9OFCPsFRVD6IO1YqLrOta5RFNzD4LWtVbn
9Thq6sSe7nZM3RW7ykY6Hu6H6O/PlwXqlIhwHKAY64IfZDb0zmHyQJtZel4ZDjbNACjzfAvPKOx5
4gtCH7dmvv0zhwOlhlW678hC8TgAmsI5wRlX8niEeR5j4HStSIr4UuWE8I5G9EUMePEsQF2Ec/be
jNKJYX+0XZGrb8bQGNFJwlQdhlRe5ESCMiVMi9CcuCa5tZ/2OCFw292bQhaEQHl+6qDJzZaDnZ7x
f9+BMepFmsQKkjDwivJPANvuQb7Jlz0uQngl5tUTbCJtjflE6eSJUmZjs/Lt3eWgk6XAy3HSQwxR
1pCGP9y6aXGS1xi3QPhVABsvUvDD9YIccURQ8KRGmOuc4pLvF2fCW546GkbE5rXoVNkav+dDzfGX
34vW06ITOPsfWzjkKzGlUinME1h0G0KeD+jV7to75Nat0vHPTnLc7+BGVE9+vxxMyuiC2+vRYcNZ
fbhBR7SXm6UEnD2Kk77Qrs0K1F456Td+wAuwR/aFe3WpKIZtKec8KJr06Uay93Az8STSi5tdCyMP
CFeB2Qai4Vhj76tjwLd/5iIVohEZVr14f58065WqQp8YUMbLmU4dZqyAejjs2uK9dm5cBtAGZMfe
0IblA8daTEZkS4iOToHE5A3J+gGeGqVhEO1DclnUEb5oIo+EJsZ9A1YH1Z5GxCWZ+yNJHTr+sJ3i
MGxIjBRLSBgh+MwP0Wl+78TUy0yID4/Q4DgmN6q9Zxi0pzVCfOkKxoUfkeNLXzEwC9y7HW51UQRj
9yyXqvCUpdcOD2JtHRxnw+RhXZ/0yg9ULi153GWxzaQMoUD1SgsJJTfpPWUzW3pEgYLENmg6neVp
RlizN8OITsLLnOcQw9bcYXvU0GIrDP0aPRrJ9yj7WgcaqUno29oDeO/FTmf0FuK9UsFDdO47mhhF
fhfagOFZZ99keZ+qbD27bDQqf5JQYyNPoIwbsEIj7FhZMKbMCa6j5A9gZc7BQIReI2i+8MBYg8/V
aK+AV9hA/pLpZxqZu28GOJMEkZ0kK9ivjdVwcyVwpfdQpJBf6n+5hN6mSdLuK+/uRiNlO9kLcwQG
aqq7JPoIwFNJlF5GTOg+obG3swVkX3EnCTsfp1eT4YZ8gAZsNp/mpyXuUVr0Ad7Bk6LyVLfHOEXG
3x+CbeWnN+nzMxTPI3SHhYvoKwkratDGSF/Crh7Sm0G0rNf5Eg00mNhpap2QQ0TdiEeN68Zv7712
aLbVi4QcKPYmNxbvfw92JvGHS95u5xugaBuZ0UQKbrKFjMCgS714CuTmv01VvXEsEKHs/Rsf9Wow
lcYm5C75C600J5dUSpCY5ynPFYlUL4UUNMup3uhRvUxLr7GnntR0lSctc7QJ2vFMmKljlNfqs68s
T4qQfaWTtLkr/pm/X8uqhE+Ix35rrPbJtyuPSw5Xt4KjR2fJSdLV7xjU6qG2YAoRYj8PrCxE3lIn
p2U5ZQy1lBMt+2A0jGyCUnSvfXwkn6F8qHWleuIdLOg8aaT1XwNKI6Bq4NG9B7hb+E+E5KilpepH
AAvxCZNDKK+YUsPpjiI0nTa2w4G5+j3YZsoLoq9fybLVqYGt2IjQ96ZuPkeWYJNwypDvsJd1aMA+
sABQ5xUsgL+PbIZMDDBYDWvQNPHkCJCsavlpGC1MtGf3WGwlYnHMVNNnCRPdHK3lcvEN4mVmr/g1
fXjybUuS4ovavRvIEn7eHTVA0i0FpflCAsjZ1NoYUXcvalcUD19O2MWUtQqVoGMNk2UY1ORDYG9j
EupVoiaQc5CRqW/vIAkqHDkDrcYO3LBkmoYnEkfpPWIgVQJ3lgG36bykr3NN55Sfp8gmHX74A7xM
Kys8OmA6HJKrWecHOS54OH5MjAyLY7957JJ2wsS03OVFM17f1UcVwtB2EL4TI9aY4i7rofyLI8wx
+nlWiU9eT59dxUta/dCwCeeDJWsup6ZkbYp3R/bQ7Ka9Bwc/SEKK29EdkTDTcEXvkQoCP/vihnwc
bLgoA6i83QvVx2Il5PqZLi2Cv2Tyn6AmVksSlR+2AXaCGktZTXKvg+7D82yT8v4f12WRYP6vHTTz
C68iYTzHUvb0AKac6se5Q96pEH/BqiS+UeKokEMr374SS8GpIlyezmafyE82eGQYDOMO9l4tM7C1
/O9BLGzBgJ9qvoXy9FHFk76SIP6VrAR3GF1X2v700e3dECmGir3nt2mj/dHVfByQppzB2wpwmYO2
ULTXObToxW6Bxa1h7/YaNHXZiw6KtnyDclpbaDLSsI4kxHHseRwT20g3KBjgLIZJMuPwD+Ve0+wB
jrD19LwczNdtUPDyP5ceDIKuhWjt3p79bJaB1jcNt6LDebRI469hrmelVqO4xzobIaxKVGtnr7IA
OXtUPWgZVehyMlhkEnDtglruWEha9mTAoGbRShuiXg5mDtdjGMMnZOvnGPVghVN1HuaQtR3U3Buy
MllTYBntBZas3JtHSkv7B1ANxjeLVDvR++CURlphPeBeYM+rh2M8Ns6hG7VVNG0UKcLXbwvidIXZ
O+ApByaHLyJ34N6vDTZgAZbAx/PFEW/FVJdfkFDpd8Fqex7yqsIbX4fBwanbzqPgVp3VNy/l4yq6
+nbTEe6MYL05IBzBkbZQzUz/hM7Iq/7I7uP4JAxVXAbiCnYLLDzSNDLoI9rrGVOfpFhFYdAAs73q
aC9h2amKvi1iJr7rigUe7GMWPKRN2z+Iif9l1+fQfEICpNf41YvYjKf2GzjkQ+rLpsZ3DwDD3cPr
soX5BcfiWCSHodNGzhR4DQew6TyJ6+ZreNfUMs9ZuVAvLZ2GpLhrscapD39outs4zp+PA0z4RNbI
D50DQ0hv/w5TgigDLDddwT4lIq5PWDoy5JakCONktk3uuJZ9/bL6xIY3qKtZSSeauDgZN+7/AYYG
/vWkR8QEvl7Y08GosKr1fcZ4nSgH6OB5rwO9g+R/8AdaxwhYF/LVnJWnvN9Ln+agzlYTJCuU2cHB
E5uzWqMkmCZz4/qPFrJOAASxImnY9Cxil+rbqv5Sq4eFU/HGwQBxBFK77AJI0fEb2ijdbjqMtauM
8H3mj1xEHCaFLqni9w8r83NP63vA0q9LMjuU2E9DhvqeaxtzdpApw0S4EZiglGW5MwOd9YnFMP0v
0UOF9xLcG3Pn+ZcIydGDiDga/KfOgbkuS2j8z/4e55PtYnf+nRCdzy6FkieJC7JKk+zr/FuCy5YU
5vCizmRFlSYmcBzStpWsc2wEFBH6Yw4T/0qDB0rkAd3SMFa9TR8Zxtjue8aFtF/ugLm8eZh2oB9l
chyCR1A6ti1r0QPuEUYzMyaWRKtM53AA5phvmwKZuOwhVTSlRvpX+votT5M3Wq0x5HQvD6WRlqhq
Mb3klIfnPGHEmbu16wMPc7owBH0eq/28WQ8B8VaBJK8t+/d2VNupvzItYcKimi8a3ceeVl26edyM
aOpH6ExbOqiBo/nSZTM4nWdJ1oTvZ+v/OiB4cftB6F81ptmes+FvPC7PW4O4aYdX2No1cArDvL2z
by/TMFM3u0O35T/EgGBjPJufy8Z4qN7kEBluSvUtCO3knGRbKMJdb1XXF8+1L/s7h57UVEf34Rs6
8aAs2vMHtjlasmwu3W3WCQD6WEiXxshGtOXbHT+DvW+iwpcIw7jRvtD8Zmj2VUDfNRAtea+u8vK2
w4SBaUnx0Ys67WOKuRYkkKfyuaDig0RuBjnU2pqLHTOWmtARxJyOmmNqFBHxq7pCZT74Lk/XAUHY
QbaGiZ6udFc5OlLzJIb2cgWDkqKqqM0KKK4aHsvv3CCKW42rjuR79NjnqLzadayBzSkvFwCs0XwX
csv0Ygzn/WI+/ZsQAMx4qyQjQTZHvAdO96OjXiSfQKt+vDq69mc48CbmIU7zUa2A97muwAeRfXN3
S+uxP2XsX9WIpbxteROhypV8TqQG5f5XojnxwdvHHjr+ClKTN8bY8OgPAcPI0XR/m7fh5fUfgpz7
f0gDNhNWNsl3ymuyJYeqrEt+P4l3qpCC+o7HG2SrbJBshEdh5sLD5+NrCt8aOvl5ePKvuq5+10YI
oEjcgT6kkl5uP4InjfzVI3wIwfn8baujtdoCuk48TT8WCT5lnQm+aO9e7RdGvjYkQdghxlr0JCss
9hdQoqmD82/YNy42vY7OVZqhNImgMBJr6X8LW/UVRFph6R8m5AwQUNmC7l5KAa2TuopID40exPdK
vEzLTSAB5O/6B5pMAfjnHQQFv0aHTL61KLU6yRHknkVGT9v/qJAWOxv4eWpghqd0nGkc//3gk+GT
TMxg+mZgW/tR9DVUAQBBaIOF44aY+ryYVrRhzcphRck0iZsaCT56NARBmrpkQwE+4N4so6cO/ByU
ZCekEL33/cWBjdw4Ix7It5K8J0m333biaO4S5qfKNGw5wewgVWbv+2ZG2z6KaQr4IBoC9ErVtBpO
dS97/Me8jtlEnZwijVnSdgHMpWeeON3NwPkZcTJStbWH64ZuUsrPQUarajJZnVarFmUzPytUtDJJ
QW+OFilOZ3/qxwcR7uKa/S89wdFNGfvyxni0xl72BVtHH3o6F3zdcBDJjPk1yamytgzyYW+nbFH9
hOz5C8MTZ6oB7LKaRKlgpGsXwRyDDZvNlCrNtdQ1/S8rY+wqPTxAIUbf/yaodt8LDKWglVDTVnwO
mUVXGnX8KrTerCm3dSDgc8cd/JPkM34jMA5IGp3A9D9F5dXS7XgU3Fgf8DkuJc8b4VTT5CpR80k1
VsklMYS1nwx48cWdmt5FlRMSSulL4GKtHBuR9O7JUWephsX5Wslx4sT/6z4dcGPdAwdsFNYJsMQY
kB4aeP307HOhYHGZwf9kr3Yn51JIAzbZE6Chu71nzSKBcPS9lLUr2EQWfLkG4L6ZhPoxG8o7BgXw
SudGdmERQiQy053KebCIhIq24zJb3FAx4KEOoHj6nKhGwkuNC5tqykiOf/lvJT0LirDSyiu14jZi
gFuqqBW9bUqnhzVJUXOpnlMERsy5JansGMcfbvy8mT2HMXR7R1TpMmRevDfNCrL10RmCt7zlGbDE
wqfX3e5gg1VtWdsMSsrntBctGnome/rxZfhsMcSFVW2XXHl/0EUiorrmmRthFsl/mopTEY026d3e
U72NUPGE4ZroOvzfwDl5Pe/nsvUZdJFxIzI40x/8pfa/mx9ZGzXy0tScGyRii7ThPyhN1W/IMO2H
DIesDfMreRF58dNYrCmeD/sBcAOrBvX9Mr6VXSxNOF6qsoTqJANooqTseJXanoWleDequJELW5we
pNklkobL3BlTi1ofotK+uk807Ii9Whwwl6binGIO2fovoE9jWlQMn3FcWqjfWZVnFR95NilTLjuI
XCsj6PLiu249FHSPC8Xq03pTSXqJWEI8c8dVTrIq3IzS6ysuZiejzEBIqLfA+gG+/Iiuj1QOkVdf
s0BmGKoLDslZEegcGPlRJjXdh05p6YgOXlmfg9nrFkrq3rMpmUL6FZa2CkGwyo5I6vAov2SVdwLS
z3lVfDigP3u7VAokceLEI3Z7gglQMiT6U9llIYYwid6cBAExPWKdeQ8tiGqBsQpx2mey3HMHHNx1
FXJezcm+ev/298LC/qb73qAtzhGGk7te9pTiFk0Pl/t0qk0W7l/FzYWAtshlzPnhoA63SyfsW73J
yq543awbLvJL1+ufD2I/HGAYWTUwHmbq1/bDCOK1sDa68ccZci5jltS2yuUoRvs21khqyFBCTZw+
q95/9FSFiZHOfVCEyU0Iaw7MTE+kSzs1dkTpLVRQadQvF8peGukL78cq+HC/Rs39a1UTeNKXRmlG
H2ANWa+e//R8yqEwO/kUx5rcx3f55Ehlf0iym1e5kHxGB3zcib7Hn3OOuwgh+kLm2rQG4Vtkzqd4
6GdsNjqczh+jme3nIMapeIJNIsaf6FAGkuzEbX2RjQ65Dt0m2Ryfc9+hVL0mbrPmxawQ4yz8AN6j
n924mIsC6qZrfit4aHAILmyA0b9OrNCdUVrOD3mRlzIRSNuYOUPJP9tKBDdIP+BwQ6+P2ZK/kXE6
Zkoqr22Zlpej49UK/S4+1UfbRD/gzONzVy+ICE5a9F6LS9c+cFjsEQSaiCASy6x/eRtY4rpcaZGd
bFBvg98lOCKvcTHKlVdaQRhXBVmXq76NkvzCQ5LhZ+DubWe1CWp4liNf8p0CH3CjB7Hh+wUVAkIp
27CNd+bPOJFQsRvwPZfeiBOUsQZRf+mV9V+LuzG9JJFVG8XCfoNm/hsuJ8TRjZzhBenyfP1PBjNd
wSxuKZUcJiYcbafTWwo1sBR0OEzjaJwB9Y0uc/UE4hE6lKrwB9OJZX4dPv385Ar7eC7lDYURke10
Lo3H4TXaxxJaRwm7vkzbHlH2ehJmKVAk6JDqfxFpt6RFOKu5Me8YoZxgUMwGWmZ7XBaYVi/zu5oh
LNFHZQYJSlXjJTT7ItkJfeIOwdLI4O5DsZqbj2PcjQVr8N1dcJO1XrVD+Lbj8azLnPRRqUox0h4m
QOBzwo/d3E0GX8uwZ8cly5p2fnVEldlnD/b7GkfY95TXV9nrmzSQH1NaJr7J1utUJL74ySFpzssT
CaF42kTSRNdxW7xb/qe6IFurJc/eB/q4J+qogjrSxbUwUVFEC5WvUD/uZlgDXNK2zO/25yBJHLIw
kyQ7Uzj6nz3sjSHdaKxSJXaylWarVMx4uZuBYxgCKfPfhyt6qNftQVjeMK4xbfEI8ax2qM/BYdfV
kldE7o48Fs4htvBvkXCv7OOaEpWRfFQutlT+ZGF+hNuNS40DL5r69oJXv39qKxn9NYR69HQS+iKO
eAnG4RzIh/xzRl4yltCDH/5aKgVQkKh1KlblCoy4RduporxLEABD5ALpexfgIfKgjAg3vIww20Xi
uamdl3/lXQXKRtbCEmusCEMUspAw+PcPxi95rOAhuB1X4r+vG30I+ReDq9CTazosoaaVeLd/VlTx
yjVTXCcdsRHU31cARGnCLIqkEOtpO030sAtz9vnUyn6s/5AuvXHttq/uh29oFmvzPVEhf9zhQtPW
HF7o6TnGy0jZnUCqMtikw8kJ0GBute1hFa+LzB9GZkn0DObaXAsXfIQ0+Ihk6yI2yOJAYRwFZZCe
SDfHp402da4w5O7yKnXoOXzvKOva67fmWdwm1Y1pmO2mwHDMbDjXZ6hN3u1yITwJwQ5xMKqK4+s3
d/qFQN/wCAjvzNqQ2C0KoVYxCW8E+IS2NRcuPtE6w+WJsA6hTndcLe3FKOzRsrUSEr8QNiDii6bJ
JI6n0Qa1UBCdE+MW8uLiYHSU4r5N2YuP7r8BmHBtVGcj+fVXhuqluMHJ0ml5hzlj1W6OtnscnvfX
6uQO3m11T/vW50qQKfwAG+rhmj+PXIuerAjM7sqDy2NJl6Uo8bGq7mDNhg7TUhZbqE6yme3OvDUH
YNTTuMjwvdFLZNsU4jCmbSzaJQY+0jmHY+lSzd+Jk3b14eWQHQMNR5f16DWkv0aHl19IfkF3/DI0
pc1IP07aIobWlZXmlWlaQjkkq/TR4qfvJ+bj470oQGBAgfheRYVB/dvoK7E8nw6uQXX6cn6v+CEF
TZW34YOKEOgCFa8ZPR0yp9cqXETIxwW/PxB8X6NbmbMW52CelxohxSZdA2tbZ3IFU2DrLv/oLWF8
JBkeQIu6NWxYBJtG/20pV2Zc6ocnTvIYH138mcGdhN10/ZQK0PyNKx2jJBed0axtyn6VBt5loaAl
ykvMd/mTmvn9NLs0PE+Siw0fqhL12OXGXGLS0H90Vicf5vR3oeT3As/fUEhD47MXYVr/WNigtLcZ
3Sto/tW9Ntdmf12TvE26ibwEC9gADNN9UkzTayfcKNB2f4azNV8pqATiiK07wIrBDKFjGphJ/DFc
iqffLpWQYnuCh4m2jsxbIZBYPA4S1ekUYiBj8Gl+DIuiXGTBX9ZaPHKxjOJ1PiRsExoKyEKZ0kmP
f8kPFvlDgmTL85Gy1PDsd9QbISkvEtUKMXO3rV7kPXGF3EkBh/jyb644piFnzJIycjTqzBEKDYyp
4Q2XwNlMK6cS1PkhTVeKvr085cPqg5AtTAOsIj6P2TjQVJ/wmiD85d/xI7NgzWkuVLJT2801Px3E
uIQG0tuluyIEM0BgrT1zVGV0FPCSgeASMxNK6o8g5uu7eNbYE0UEPp8kcNa614r5xaPlJax5q7Ja
csSf/NvVLZKNESx6xQMjqJhovR7lUN5g65ydPOlplZb8knpJGzu76vYtt+UjnZsjNny0PxQmNWy0
7OB04dfxs/Mhqv+CFtsugrgjXnCXgMjSqAwrsW3Xmn2YQeGiv2roZW6rP1PQI4NNMM+KK7RZc9es
ifj7qzWJowGALziW0dz2NhOJtEeXCfmEc91D/v70yJAr2WSnY1jvBwtDvYe/vH4MeuVJmJSkDLm9
b/SoE+FzoAw0vmLbKA+FZEypUSH7sLrh3G2rjvWBlNv2Ib9qfqZjuORkLF8M4G70uqLRKH1gm0sO
Mfg0qmrZVy2eqLg78ZZ9IYcCQMbOTxcidPpg6gswgVg8a/sKqLVNe7agMPEu0CuZXSkvcxFJbm8R
bQHng+ywU8le9gvWJGPTJotwlGmFlcP+7+tYK6H9UBAsxSg9M4/59oL11TG5ZUR3oYIYdhYdbzos
QfsI9LX0gXvxKQWKkxQjd9bAkWxEdlSXOIBZPz+7kOb2J5UCesNqLYE//JEoOv8yTUYRqkZ/uPn9
JbPILJKvY1Zlpaj1sxH8nJJQXyLiG0BxxugQKOGyu4hi5yxTKuKZlhwL3Y7onnvK7L4Pzj/YO403
ZEHX3OWqF7rIoRtbppZ1HryS3ISG4wmX0N6wCCHjgX0d5VV6Z3Keh8YX4e8p0BnwGZSHQtPsw6TL
Chn5Et10Iu2gJK3V+B3VJQ9vEOFjLVuvHNSd+Y09pG5oPvSfgjD5REKIZmLpeQoz5akYnS+6dqEL
Ex5N1KHPUFa3dCTOD2p3DYCWkwNonpysKEqFrHgiejHuNbrwdoKBPXJkos5STnOuA6bRnXKD2hr7
SbgEuAypENhVlt7Yc6dwLowZZOYQchBCCJQJZK8tlaiMlJxI64YW7cJ+E+S2wZLMAaWI78ka3cR6
ELm7EHWhgGZdo6HYy+0Ep14+PpYBMhIfRtKbBt7WeetZIsymbl+VA7W8dBFBiQtuIXzzkTEq+pTN
YdK7KwBly6QN9TT/SMyGiWNoZjnLD8cByL2RgRcIYqDkbGvRHkEb4fQ1gY2I+JkHgLW4A7/dYsQj
hbiZcz2dl65H3Fwlux9EOS+a9UBqzw6tdGzgJfdc1bYEQGO8Xfp2gRJcPVpifdRQvhbQr3J6mgxr
iyu6agRBGUgW62D8Nr4r1q9Lp/eDMcbtIZyauEQ/Xa8ncyoSGGEgboZZ6mn/XeK0u8Gh7UbEIAIo
Z1ygnkauRQ0aBUeDraGrFoPwnwMkO9eTn7ybJMvYHMS6orzW0uP1IUoJI4INVOy/YXB8bIsRPvCQ
R+9UanUhakBXomULKsml3q7U3Hximkna4ix0A8BM57MD1vimUbKbG2A3jO+qbLdVwEPzwquSVnFH
PKV9G9hK9D6/FB7xszVP4Z/uqVcKhK3iXmVvxKCH1NTHpwVsTwj55S5Oo/WuzcrDd00ZLfa2TqN0
5zgB57MPOLoODhw6TSTBNIxOWGqxVNWNAEAWd/iA0VdcVn7H4+gSdsvOikmq5n1iiGzcb2saf7+9
7ImK73QKeQqHxhREec7FmXFU2Bk+z+7NM1qa6QVZsYjGJ8wJd2r8g2N1YnzctVm9f9qPCqfDNWv9
5W7Tz5BXpOasWgTh+pUnuJVDhNRDfwIxVIzz1BaOqKerVzMfLaYtcy5/BZL7tsKJQW+FvsAGP2mh
LRRD7xsehRBLIsm7RovK6rXIeUBFJqANXZN/IFSmsJlhOrXVDLLUyj722lX5iSXW2OYfDu7wrPoo
VE/uaYtA43CtDyVXUfmRGGxWR1y2tfc2lMSzKanBBJf5h5BhgIW5EI/vtxy+DRYdJBM/YLYHq+oX
1ptT7yJj6FG+qk9afNYFAXurEepl8MJ1B5ZgLdBAWK60YEI9i/R1guXccxSL2jy1vlQ4dgdU5DKx
LL9Q+ChtqDU+jl6ShHFhVOd2MUmEZ0iFoKOFVFLSCTSIRM9oAY4+tkGsP34qjIeQ01HgOI8ZAj14
2HMtv8A3cNmbg5xd+7iTIqifRP+NNjcRBr6sLWMFaiHbzDjUZBRCQkuwaynbU+mKRnoNqJWRyaEj
LaeGrrE0aQyju8YZ/bsj3dyq4WuA/AXPrf0EA3FJ/btRd893NnaotvXPHB4vJSdB4z2npfI+jnqz
09i5oiqfbUtrYXD0v/r6BYzDRnatKPN8BuhWGdtCdcik/VyfFl3cYT8/mL9IrUcjRINvrPs4zncZ
atAVueJCP1golnBas16Z6ztpdjsOq+oIfkI1gVKylF04I1s2kVbp9doDMkX7tN79btyCcCj84wJu
OfJb8c3e3pc6Fz51hEFyndVQLVefjjj/7OoYURtA0S9KMhIn0qm9UdO62aWZZPseqw8p+kyKs+8X
09WwmdeC9kQjQkMR4NES0QVRHD1tPYxwdghV5UVbxlN2fjCMDBGeMjisssbSk9Ll/fXmEIiHUQm5
kk1651eP9pbUYr0ck/T3jKwStafPWpJulclUZw+0DvtOysAXndwzylhC84v9MaVhlRujsgL48N8i
JmVaWNtdHLqjUq31Xwn7ESA1YByvR4TJgE6DxqCMYSKk1cJaYAie+NaUJtd/Vk00EPchPTzEbcO8
+r8NCGyqnx0dtW63CstyowWapPbJUIfRE3viy7qL4piZEd7/yrQu8S34iHCSeScj5nMXeXcSafXp
YGX8b1dktc360SXaYKlmjdfO64jgcD6vvCqcZ8+++fci63kCTonIzO6T/n8obr2K59M94Uyc2wvE
y21g35aSRInMj9kp1ltkvxd1ztROil7o6rcX4ZgB2fb8mc9/qoy90tzNTqummJIyMRen69pXp74S
MrkqA14h7EDRO7exmdzpFMMpiIm5kohF8479oGdDJQIW1/WD7tfjoV7J2cjlgks7rp9f9+NhwcWw
+HWA8Ae+WqAWOtyf7tE77oC5sAKSX7L0k6NHcuND+uRjODj4UJq/0rW2NhuuMqqzfihTJ8vlsHR3
IP/ZSTz6Vg9q4dMmti6rydZCAdhGIOGjnWAnqtHCwGNqHDGsu23T+ebVvfb6k0DfNrt/0cnNjf2Z
WRy34P+9zaNgXvOCsJdTJKw7vgc47orBJXwLvbHaEq4DoB2kIqvhpMEQwvq2IOFmMpSXZB+TYl4C
4F5VZrhpVfsGIYJHpPzJkqQSpCEJhIIQ5KSxxz3C7f6sqyLApB6tc0znzrhDI7xeNig6rBy1jVoa
7VA8+7gAKGYm6pEGyvkhHK106Bois9v5svAS3zskk44d0kULHwnQcvO4/xrNR38wjmIH/vIX+QmJ
wnOCSvwNMerbVwZSB7jX0wBtja9VDO0wlPYaYHWkAndCX/I4iZrj8EjzFHGj9VtsQU27EBgMctxZ
g3Y7BXjIU9cq7gXNirbrz/kTZeohZR6qdv8MjCd3QY30v/PaW/uH/N2JFHaHMXMbnz1iJefwmq0I
jQk7ueKe4gI1yO1GnrtH+dn3a2AQN2GMOzS6Yj8AEoHBuBsn2yTqlG+riOujV/z+aQanmTdoqwnl
w9UVL7PN4/Z1G/rxLrfBPt5IjnR0tu/hTay0tuAeeps9C/C6wabIXc0U19VKERtGuXWzKNAXHcm3
zRfnmDeoUTxqKA08AaKaUTjOvz92MzkJz9ZfBUGja62GFrCOGavTFltjk/ggeRCNK+uTAgtzZ8B4
KTG/RnH0ns5WZHgwWjgjDMiVCZLc1avp2GXPhKTOiaSrUNyrkBU76PXLF9njQic3VaSsCA4Rhv5Q
j0EB/dLMFJvdvB91D4xP8UIqMsEA6CT5xMlaa4ty3L0GzEjlmSFUQSBHMgIq+q/F7lTxJq0mHwL7
ewwFwtovj+gSuGa9+kFJfiLwo4Q50q8esYN8MpJ3v/K11XWlq45fSJNhk9AppPKNtzTGQRuahAr6
O2BQemje5zJS0tmMPlxcuexnoGgGOWkcbkebuE52A0l19Flt1nngoLhhWQ8u0fN/je5Td9Ivqovu
tbx4DO+cheJoP3K0/Z3bh7lKHjcdOLA6U7nRLDADECD1XQkFtQrTMl4nKITcX+1D9hhqSWQR2BZf
1NAJQZ//u+LFI4JW+BxEi6k7aApZYps6cus2fh+I/9r6WiTjdpHPKrTsUfmShXFGVPUXxbMNZLPU
K4kT9+RVd//42spMtFcgPrZ64CtIIDwxPLPBqA4GqKcVJ/8pXh6ub+0zq3E3aRyU8gbMryVxCLPp
RlN5aa247pLCcRWrfLbDujp/DyFFgLNRg7lDVxa/KdI9ZWypVus/d3cbXU9GAUpdFEzVWLGVMA76
Xio7YCVOQulivo7og46TOEI9OFzQNyICsydcdU004XY4jIin+Tip1UaCGkyuEQzC4QZaXRTHxZsV
EXN9F5+eb8X1Q6feOYk0N5/AE9xsdXRvHNSPSCCMr2HCc34UNWnTxjeMxs+ihvivixG72ggitiqK
Gcc+nVKxzytmvIhUYAMnyrKUVynVaO4ydKw2gpNY2vQ8ym6W3Jx1DrX17bevHUAHU9yKiiWkOeiY
0CAXafisfIGXYmVG4u/7WDp0LD/rd+zvg24M+5krp/LiPQcXKAxN/tJYsPYNojZsx0h4HX80GKn7
91+DcXfNU1EBERot/1x+u4QkdgM0UPsxRZfN8B2QYeFDGuJhGOzlhoOlfv0nn5GkC/FNOI0s5alh
PR+rFaztiYv4K3Rd63Ts4eGVQpCs0D7Mm/jAknMkAgRSGXqZ6anBs2ogUSXvvumXML0egWrp1Rhi
bJwoUMwdUlJ+oMU29FOAT0oSaWh/8bksMF2hIbyVmXPPg1+oB3JVMe4WtRuskMdGdZpdvTnLxqRY
K+W81sHL0rc8YPHWfkrZSLEuuaBPgHIfm0Cn+kuYs6bXQ1rjbvRGTeiJ4sdZbuqsJdU217we+q2m
Vng9ZYeqW9R3kyJqfDWfyrOtW/aI0DoIe52+jKCLH5AaiK1xbbrOCRk4LesqkbWaJ/QK6/0p0RxJ
z/c0TTZpsbJkkjw4EgG23ICXs4qeVbEbsv2bvTj33sqPQLJXstXes6AUkUSk8euIAgebwxqKgRIV
V3c36X8VZt+X0w5djsIK+Zt9caWX5Wkw8piAYj5YfREAx4ChcFQroXx5ZrgQk8eGeEjPIYOpcPZR
KXN5gxO7/LcEHjb2/pzmCFX03QYkNwFd4SYjAyc3SzQQa6oBJ+gTKDGL9BGvq0h+K/aotUKCHFWm
9f7zlJ/eS9B/RyKFjo/XnKwkSWbx8NAq1/KNexlRW13it5CazO9i7Qt7dWM8iDRRW7rznfLmSHL/
GBI5Zs1lUZ/9kUIW9jCvx6Q7FgBnI64LgKW5ZKfzZyrsTb/BeHHzraHlVOAiHbk93eVk33QNIM3p
IASj/i6HU+qP2dbZHs37j475rJ18e7BCA+GEdr4XcKgMImb5LXg2B+YCoT1+7mexlwyBh0Fdd25B
It6vc6SjzHie90Wcps0nOjHrI64Km5ACL0LziffdiHN1pibpUSq/YLWqa84X6BbTnYxISwo+Zf2c
asZ3CtR44sIP3rhtjIe6KuH1mkJF6HJod+6UAhDGSEFQtC0X+VxCTfOHkdawAhuHwXrrQf0a0rM2
O9yVeb2PN3Jn96uepB1hfaGZvAVZB6Yl56uIvWIRMQNhPc5wJ2RMlvO3HtO2+gThTjKZ4eKIQV7m
f/mC7UyWB/Bf271IQkEIMbyxgh49CvGPAyhwRachBgv5vpfOOIuld5CVQeHDbFwEYA62t/TUhNC7
Cdx3horz4ZpvsfRJwwDl1oV5fBAmRpjmslyooNro4ZkZ00XhgP5ofTdlgKVKE4qmUPF6m93iRfmg
IxVwXcTMUwIf5WG2PquWNadQ2Oh6cc0WbJl8wHD0AztdUILvUjIxkIhb4wlJQo1QPvsqmbprfnmC
tMq3dh0IwLDKMhi4E+30s66MShV0iUIgjEEEKuJFJ5Ktq+Drgp17ZrLguW9SIxftU9nDTynOfxqy
StW7a1Cl/ztb/1O+y5L0xQotCdG2ifQddRuI5vKHKxH3LAqOailUJIasL/OMg0hasVRBzTmFg+Fg
4DD2vMwJTcvSB1vkNrkQ2VSKnJgtlVErHC97z68vNwKTAYNevuaq3uBU8L2ciB8XCt8g/IX5NmS1
JQXJnv//IDRp9YqEkv7lheJ2HpQ0++VBzmdvGZmpqEDikOGxoaHxpU4TqYE4kw8ngyGEe+OZgWLa
GX8BmIa/xYKU5+83/JhSWwXI/NetOTz9sZwC0N8D+uACB0l1YC9icw5symVcdRY3k4QowyVplaCx
lEtTBYOjVYn92a4rhzHeQ3vOlchvRpY/jzMwO16a20ag355xt3OcBAuphkcVS8wNcwfaGBZs2nax
a2MTEGM4nrKkrgZsPiRR/GLV1xb8M+CIepfvHKuVk9KuHm55RbV0WTfIvj1lZWPqzLEtFkcmixpg
aBy51e/NMAklhNPEXNSWcdii63wt3Q2SjXKnnBeJmQa29EBsjBQV3b3NRjV/fkp0/NqqCjzYvjRk
4wKKT5wuM/eurkWbUQOaWSw/JBls8vZJRDifTV/vtMGK2QfxCZa5WOAIM840t5Xoep7XYzxG2oLk
CEmCaEywAMjejXnCz/VnSSzEBX7UEs3xMyfugsw2BM+80xi2Vp7rRrapMGPSlwSl5eBZDBqB0YcO
OPyDLuf4iOqbRpdUe2FFAexUBjMNtIFkwUe+zXyO8NcKcDrYtB0hGv6X394dVNufmKHtAp1q1MAS
w214JT4pMiKa7JAK+FFDv9QM6lvLrC1By7S2cZ6UAOueDBm9yAHFMI39yDgCGwo5+LNnV29rZIYd
0WIpHYikSHFnje2WRORiV53v3Yp1s155NmLd2ijFMlQuuYcxzdjfpg9rAR6QWhmWPOTExDUdgugv
q4914TME4E38ELzy26PiTg6eIml13tpETNjfXIFDBA1kZdmRFuZ5Qb89TJUhfF44D51eCtb4z+fS
jHA+rt3v2F5b70YhZaVV+L3zlpXJkz45pqrvduxgi1ENZzIpdsXdch0QeBFM0gdD1p7pjwt2TxFb
er2lDIYPGhVCN6P47tw6ixKXD2bFXFHfYOrjNklIhI50i9v3HCc0rk9uvRrxIY8LDWM70PXBfOFc
1h9H+H0vgpkAjopBTGg1J2lqWOx+cQo0Tlsm8cisgNI44ZkpEh3gn8Z16hIR4ByNEKXW4QXCK3gp
Nvqn4WziPKg13MizwF7wHDmr18hxQPxgxTNDX98otC+jbdLkn/zWCXJVXyCVmFclvU0aaCSU5ZEI
9cJtD+ZFJlHxoXuC9YU27x0BTYBo+PSZqfQ5v21xHF/E1Oqi3jD4R7k3pUT3+yIBhSrxnCIb4VIN
LBhVVp71TXReCaHwoea4+Y0o1jxvJhL++k/Fh7XkG5/xB1RXyQMA9Aguug4IAqvFg9fgE+YPXIGq
q4uOsNjhhT+Lb9/lc+pwERt/c1rAbaup2T4e4l+jbISvA6g5/xozioqgdmGvMyDGzT5U5FynfA0u
N6zI09300oW2kmNTqcL2SuUxKNuC3TOCetECc1vQH22+MLg2P+TqXufspCuMbJo1mAD4OT+2pfGd
3b3ACHbcOiC7Yq9JhGWcnOqyhLDRgQXwuDo7uY9tDDp8l1yXwFT38J5+LsrR3uyKq2W7FSeIjSJm
QIZfkLUhLbHdj22D2QbDCLvKAdRIDJAizVkxf56o9bEw7d1MiAjc+WsKvznh1lt71AHYpYJ1xm5h
/cQIMA2j2ZSzBSgcLGlDS4MV5eVdQ4yRyg/Af23dnM3g6xeLutLApGR2svj1BqMNEn0Td6d8/Vbe
YsDgEii9FlHUHY1GmR+7vQyyXZHqGdX3NLkHn/PloqTH/Ux+gnYnJuHCbcHwZ/ZyZwoFZo2q+gIq
Ba163Dhjk1o1/JqRQCrUhgsM5Ft/qh5Fm/m25Mt1lTzINZ2/h0Rpy/ecHxVnPbptYO+bPrjd56xj
5xszR9qtgAKiHvRMWSW6J/UEpI+ELTbQGXG18/lBDRztjys80h9eWwtQ8ZCLjFvHFHvxJENaVlWE
LGV2sTE1cmEalzFO8C9+1Kks49POXXhjTpu7nah7D+RWY7kTlHa0EC/CaiwcRxbjeeY1BU8sK8S4
46JoC6X1kCvsP0cC18eyJbwdvfrmcT2pyGS90xd7TeH6cE1OBzeqFO8N8j4x5wMBTamg/vv8FtVB
jXCeUAJ+ZNObzxDS0/JPAdTyBfaK8iquYOh7pFBjHKUOjXZA1R6vS1kPzrbkJ3Fds+97fvMH3ULq
v8rNkKvQIM1+Wkpo2vt8V+Q5Whli05VUBxxOjYMoY/2GgUSdmh3LGQ5LnxqSjx3bYspPUrLztdjb
6qJWgl/YeRMY+UbznBo0JWjqXY8MeqG928NIA2uHi5Jwgt3ODztijK4HQvpap1zsYXLzvLrWk33H
XRPO/oNti7e3sOb7bCXo16HQ0JmGQcPEaXED6F3vTnwyNNwivEl5qrE0Pk2m7sVFBXbCmuChYF6H
YgOpUsAfmmxraEe9djtAdNPUGg8QVxGuUTndAihfeOoXP4fC68II+irQ24BS6CxAtmJyxniTFFZO
xf4lPo57pnNzgBkMR3Chbo3ZB+4E/wMj7eFK/j7aW5KAUzx3rCT1iIvxCNlFLLhoiRMKx3q9qqok
gA6jdVl56jD8VNDDlaRZ6i8fKWFmR4jj4/k3MbaJgr9dXsgGlmCg25yOycmCzOXTwy9P5UPdl01c
53sa+c62tMvpx2OlGJ+hDxJijfcBV3dlV/PRqjZZqAEpq3d/PBnJeSVFp3Sd/QXG5Fplh1L/5l8z
aeHkXs0+qiRbsuXScb5wS6zZX3JkA91eN17nKIjgk9tKzG1JqjjIJodcsKpW3uO8X9oilJGBPrXj
2GPq97Q9z/b14e4PYj9Jg5iFghSit6NuX4wKONfm7Gc1vWWeD040c9srXFGbo8ARRfjyLBmSHg+4
EyvzVluqBEOkrYLyASrIbNLQlXO6d2D9C/Ud7SuGwbP2OK1Pce7KBywwo6L355YIhwF3JW3tZjCk
j/9uc3IK4wmRsRQa5GHKfIh/v7t24c6zP1c3py9D15D1c0y/JNTlbrO3n4+GZOklZT/keBT2PT9k
0jnNSx3imiRuV68+WMW/yt4EmDzSPylnYeC5ZtPR94rtzL1iuONKFpwjvj6/QRcN1ymz1fcBTkkV
0doGOZkhs/I5LWTX21PAFVx6cCrnFOYWCnLDN4hZSqMg2xvmLu7ZHdkgZIXwm+MnHibDHFNc8wU8
RbOwMMMqCIl1JTdAHwQvhxPsIe8TezNYbLEIZw0Jqhxs/xowD2OBywjkjY92hHXpLWv45THUxcgw
zO6jte6tOGNtPQF2MVHQQZ47P/JSowHxi+YWs4OH8Fkx+JwVYLUI2JFbcgxLtVnTzoJUmARctaiL
nawDsrvgA9zjFR4zu5jPVYxzHGfaquCs5zj0yX9/SCu9wD3MY50gcGtc8Pcj0NXf0D3YHCjc7kvX
eq8ape26PlcU+ZNFziO6z1HZ+dbrKU+rmOBIc99D+sph216/4ZLE0JXTMvWzE6GXQbb4tNa+FHuN
QFD6vbh3Zzcje/f6TJCCoKXBCWunL7/cPA7oAXX0EHdyLvqyGJpN1qKxW9olaKHgyWb5RlWZ+j+P
CAOzEpoy7y51mBfJL6CvjiunVZzJReFI552dqgXwHs0ziWJZXiGtS7CLxx54ZS6Hl5IuVEaVL+ue
UFKVmJOMCr7HlBVi1Acb5d17XWf0lCbtynMKPZUwRSaNzVIoFRCs8c0HhOsvoVXywGTIiO6NIaXN
16NZv7mTKT8QAXCZAhXa3e4YxJvcjyvb9NJ24OaUyHVsFQRiL0XCye4z0/EjFGrnxeLecKfNR38B
jkAspxaM7IbH8l0SQKon8F8mCER7vwBmR7ZG9vaFdix4Pq4NfIRBUh2uqifC/6imJ1xNnBmvApGP
wT+jtp9ydzIsFJhX3PsrC/7XBI3w/zmPNRFaNx0sMR0n4Ry8OksSiB4CE1BXe+esMSYJlfP/biqQ
wiPbBgjICNJUgptBe88LOKCmfyce25lVHZ94BUOX3OkbsFgAj4TShYvG1IOYTkad6sRN/UnsWnb4
RNTQZvxek2Aa2k8mWQHeM4pPWoR7Es0TwNIsLmuoqdy6NY2BcoSBquS8J4h16JiEXbfoSyfPzzMA
VPCjtnvaol/0PiXAr1qf18OCiXDcXvbgWvj4xi0/eu8gRs/a97Mc8o9ZJQMJ1JvEmcsfVuvtIXbc
qnU41IQThMm4ZfmA48juAuce9nId1TcJ8xHEeWBXNtB5BYu6D5ztl86OAAr8udIJhEDvuaBEad9z
KFbXqSlXMl9ToAXR5tgGmbq8s1ntkugOKaeJ8Ka66rDTRqWJGDIPGsGTr4Y2yk2XWLN04yzCS38t
ycJcEKGWDqWNAVl2pgvxc/PH7JYoIm5igxAlBjSNNPSdTqPadS0ELFy1P5dTrvL1lII+VdVIOQr6
Z0X1nUVSH5wALDOWSVdq4zQV0hpoS/c7lceaoXQ8YWHjGZM/ai3qVJca6wmJRgKu+l8su3fWaoxO
aydK5OLzS1Mw4SfdZUcf5C7vk63fGi+oQZifd4bapXdd0vTuo3TxjCHqo+d3tdXDHF1bKrZ9EZIs
BJUGQ8a8nEfvfF9cOh+cfeKUP2lWk5mcbVmYWa0vLqbbZUdIauGDh2s4yW6F/mtDfxOBuszKLpOk
1hG3T2+5sCZBXD8vvaqdDxuML2OY7jlY6KJHi/+d1cc/Djn+SeTIgBJs6YfE/+82a0qPZUgh4duO
5PWb7P0MWp3lt/ofIIkLxP8nj7A8T+UuYofYqwELKGqdU8I8C3RQ0l3kU6tTprQwJHInXbtLkIeQ
yvQhCLhgQIgbcOn7raYVaBmBHPfmhQfFq5iNWkSLjUFMNjrGxssvSK2CfoP4xmCcFNEnL07xHBVP
ETJRV3GBNDJNut+Ro6MLITb6ohfzEtZHEtyYJLE/G3miVmG4QNRPXWWcqsamSa4R6Axxk4SgztdF
vk1oRmvnqenDllIFFfTXByrlzXJM5GlepjwAROwdfIoBV9KCTfv0ET63uHxPrJYeYEtwf/DKMypd
6PIQABaAYyL0mVvE9ZsvJTPDOsG7eGcrxH8BMBXT1qYpgXrLLaGJ6Ko3+pHgQM0eRGsvqmGcTTrs
IMm2D/YZxbLCEjaVUfCvrxjFgYb/3wGep36L7sxZWoV8aolYbFIoFt1f8r9GAqCXYoVHAEewx80t
luW6rDFijtT30GBz6ReWogV5lhzGuGi1qggjgPZhJ5g1CTKWwu3nIhrGsUFEbx1NyoQtfcHIgOUZ
5Dh88NqRNQKDriJnJzUHVdWqrqpDxGn2qJsbCxyp+tLxgLvCt4yK6PaPLThPDSumh7xC/i9fzMyL
MRWAN8N8M5+apOKoqvzmIk7stP5nGiWQi9Eky1jqD8VWmWV387uUl+VsnkNLwW9ry4fH4WXL8KJg
LSrynVHcN9RWVsqXEi7WBd6AjLWZgUxboQyKznw0rZeZDpAdQTeV2Gm8cNQEkHp1bkfMvLct/d3z
xqcJwkk1pPAreQuVQfbcQEcHWrFp9VTXA9oD1ByE5gHI33/KoM3quZF33MTDtcbJQiKt/6GJbw32
791adobjeOKEhaWlXuoRTZxAbuY8pC8ZgoMR++hT++Xh4kt9BZUwvItMKOWHodGaBtMxYjNtXcS7
IZZuew5jOo20A+csHVXSIRP+B6zKtNWMxnFZVNaZbQvtEa/Wn2RLYoy746+A+u8RKH4wXnYSOwX6
aIYIvxtvArPmItncY5MkP9bs7Uy05MKurJDB0xPNnyLGanUIT5n6DJ4mhx+PyIdee9hjCSsAvDyI
+j3rgFME2YxOVe+FXcrIi53JPGYfZulZaawYBP1+MP4Xj7xAIppKnu1k8+woRMxblIyjGMWau1cA
GImaL8YCetA8slRahju/TiiN6cePjlZk5ubiyp1Td+m9MeUOEHFPtsX9d2nbDCKa9my7Az2KgRwP
p/lnGhmx0sp2wVckRBJxftQ0aM5yLQOyadFn1g8fZ+OJ2vUPfEABMokYF8DZl21XSiAgFRpkDqLE
Pk0RE0qieTSHoQbKU+AOtyoBH+OzkAYd9qEWTeqyn4vJ0gnhivPCFwnDGDEQuqdIgZFFQEi/JL/F
wpP/Jb/vr3ztdKwdwzGBlvZw6tOQ+VrQIen5cNfbfJ1B5W392p7eln7HspugagcBk0aU+zltppYs
aTIqwpyqpjkXqiOKfgSWP1/vTg/rKRqD0fMrHQBdzaJ10wTAKFAuznAEgYlIyzH1ozotR4nyPIB3
Yzzmo95+3MwdIWEgpGp82Qm+JYYBgrlkk4viQ7aR2btXACuZumSF625fM1QFEO4thXo3Txf+X2C3
qugce90M/+FdDwpaZ008KNrAFDEkAtqzXsCNWiyDBYyYxLI3W412UKU91ucvAGbpQQIxYdC2TYVZ
zLGsh9tmKjllvwbzHc46SosfEG2ZRNpjX9HyuZ4AQ30ZrIGRojnEdl83U+zbqWpDQDwRQZeZw8V/
DV0IzyRfdl1OIANLuL4l1sIWBL9egYG3yhAPvdcVBGYY21240tCEFSseng4netSNJgroErWGSljK
4SeoocX6rYRt5/UTkZwz8v2XNbjsKt6G6POs7GXoZ+PksoQhdNawToetEk0oH3fn+CpiO4OwuRYi
Coqte59gKHkk8W4FE33m80uCbdxXKK/ihNaOf790HXBOBj4ow5MaUu1OmVke1BR29B4w8aCBvDtj
AcpOTMn2FZtulynp7iSvFgGrp5BEbxCkgnEXdQjz+K0rt4dyuAgH9cSznZ0ONjgZQIhwB9bdkkWN
1Hd1wUi3yW8X1UdSbXHr7j4No1jUHbsaWE66f0OmTleT/0je9d8Ocz2Ghar9R+0YS5MYJVEjopio
t+KbfIZZIai5To0ts1dG9rqyAwxynwMnKyYb4ShjkwovCBKD++sl+XYOkOeggQApxMQw3k9S6+FM
W8txOwmmluAlUFfP00j5hVfvPQXGFAxMb1BbovopVYcM6uoNoKHUTSBf2IGSbH98LysPVNxXb8ue
IRbi6nDJrWoiGRRtQBU3hRycF2TtD4qEPuJmtCr+b5hwcSUxmIgCiKk1WoWoewz2NDz7D0ltxb7y
iV+EKk0PsNmQyP33LZ+0s9LS3yxmPo/r1XjkkNnBMH3sbQFIaQPlXNpdmxCo+2U9YsoXL+x+WQ81
68QPcyAm53hdZYqpZlEEdfCjqYx2Vqcov5GstdJa9IbQD5Nvq8xS4+8+CkmCtGdVRo+F8kN8Uv4x
loC9lxF3xN3aOqjgVai2WbxfUtxhQ4dNXLPAsZGWfSr48mkGZQ1U3WwS8M0ZVHGcvQyvdYETkZZH
mZx00v0+Q8ykhXZEVb8o8oNii6Ody5ktyGmGKdVDdBMDARAYext+sacI1ja5lFaYI43W3qdSPRth
DiYnrao9JiCnB8VrQE71Kk2arYIgrHiL0OWR7rdf3VuHlyp5TGJR3rHbgpgzpIQW+u/JqDb5ZEao
0jdMzZGsnTboGpDX67+72cFAWWIHjXocWU1wNgc7fxLy8t+RtJXLa4du4xJJKUkidDwyywJSS4ib
c0X/aTGhBdH8090eCVKktYvmrhCe33aChAjxZEXALlRauXY538y5Fbqco0DsWC4SLcmHWUozaFiT
FnIiR+Jt8nnV7VixAHXWLN3JWOpKwYKCaNJvDTfngPjVPNk2uWRIzrDkXnb8nG1nb98axoOH+Png
eY86UfoIiPj8M1oN16Xbnp4+scJTrpQEP/75zMCyXW3hcfkTCqL3DZMbDl4AaHZGgZi9P6N+LxMh
xR8O7yQLcTH0kkxXO8jwwnHhAH2pwFLyrO2uI0nf1T8SF6KTbkx5Ob78UEwWDP4MBkCYTMiUIFQW
WEG8+wrF/EAtIQplUWhv88qJ7i0sOCHhVsKWE0SJ/YaUqju1CGRkXitWn35t060574tDOTytSMv8
8+r4fVbDBe5kEWezqIiWgCwaiDURsBIXh+dwOtpXZCBOGrRcT3+z7R6xk88HtHZXnUjHKvfRXtVI
NzQkn2hDUlr0MsXHeAPOyyuR0PBF4dBd2Ss/xQ6MiqTbCX18sMo/AjY4LKzUmYLNDM6xpNK7Q33I
BxcrOF6VqSyFz6j8XCEYi+ybM51AaI5IQZICN6l4qN3XvOr4X7/3GzW0Xfa3uIEmGQusiuoueG/X
164xYQ6YLKd2MP+UpElp8aXTieCQN2Lo55EniZKPGpl/qO14ulAwY1Ez5Qra7uEphnbi1+rNJDAl
VwReKhbNBmdd9k/P8sjrAVrU3KVURQs0MWxvBubjj4Xre0qJlzwCz5g2q0q+e+p8w1mse/5aOPwj
FuWMf00XG2xpL2tPZX8EtA8ya13LKldfWNBpq5AbG1/GeQibVdtywME4eNnlgMjYDEcSNQ4wVp3Y
bcaHrXFjhKTuIepIAym/TExqvIQ4wPLW3SdJmjWEDBzb/0oNg5/VLNvjK1qGo1ILPum2SUbppXm8
SYnvoDcOAN8MxGXoiaeJGQ98fB2EHOmzSoPPgljqGdcuNwVl8EU/4aTCUvQMY6zdCRwciHLA4M5u
Hfo0YRuy42fU+YAdtLqqoCQ8vfuhexV6NgVK5yZFwKyt7TsH1a2VcCiN+Ay36eUf1KVNgUOWw4bd
hiuHy3J9UpcOfJ05g5cWczKCXj/mDoJboXA2LcIoI0WZZXtMCEGBMi3oFLyQvh3UCuihCC74c9XO
ZgupFYY1ZUiuVuMceEB2v+FhnL17T7bTd8nBbgbkUQET5GzG8GLXIEmdcgt6ZSSj0QiYu/Rdu7gW
suXJkd7ImwljT4FyrJ3oJxV5MFhwyGNZhgkGYuHzcXq/QMcH32+rCErHttlSN9YZVSrB7IplMGQW
7FR+1EvpC2srD6LAAFSdyBLvdr3WseLSs4YF0FrHzOU/mebhqwyherXN0kDWGz97Ht1SHyQ7zrks
EDsXN+D/OEwfDp2xOKFymib6X2iDS17D274BAg4FND5L0P/sE/0ed+XaoGWuNVGZ7R2GMq5fbYs8
AEWsLZwK9y4OfTTdM3gF42qN4OhB2EjtIsNegdHJiSdhiAR8FSInMPfiHfiptl0HB0flh7xzV1qJ
KEj/4kNTV95fNeAVKanwhAwMCcpYM29CvSZTidf45q/llM7GP3j+mtZshRPEqO8CNZSw/avkPuNE
RLe7rA1dLL7XkeQ/2krJmuOR211wv6bsABlsRhKO74/nu9X/M+R2gjdjcMS+W/iiiOVoVfk7+3qo
EFlXEDstkQ7FD1nbdWVF3QEnUSnK9Lx5d1n4V6VuuhfRh7PUHnDGAG8EjU7Qkt9FZerxfaugLw+y
ZkR+g9JoTg2TIxEDC38buWeiXPk7K8jLxHS7fTTp7X19KrvaVfR5gCAaGECr3wJma6IrkE2merSM
2oKg8F8RRv0Dl5hTUHqPk/yZs1jKVuAXj5LQppVK0jhoezosJWbDBO1lqsJOzycX9O/Jdj9NVLFc
iVrqqeaRkNKFqElFqqGrPfopOCpSXkjssd7FRNB723v8L0eR8u6zqFiYQufoBRh8Jo3cafHBeqT5
WjGBbQvo0Pi4l9sapfrhMmsyczrEjOQN4UaFyYcXARI7TKDAsT8OkqqXCb17Myc22pYKOsKOkoFm
Kd8JQtEZf+AdBweUfhc5fxE3XLQLSpjOKFiUFHLAFXcN7YkIARi6kMBAzaV7fmq+k9br8owe+15y
AJm/xPVADDv+vrfdatWLJ4IDg+67iwFgyPo8lzuCW745pzS5mBPBZmaXkEnkPLwN89jqfNfB0AI6
gm57x0TFbeQRWLS+/3obWqWc5Lc1d3BlJcfXDUf9J7viIJ5BZtJPutCSKNMsH6deiaMJjqLfxKZB
JK3+hXKW4JY776SfSYotlFEkjcK7XCvl4Wsex6itwraT8RShHaWq10sKz37MvlyqEb/T7+VeRoXk
gDS8C/buvj55AdFyMTtbqn1E3rOGbammlaX8tv/J2jsyjcXBgBvN8FVtLpc8e67TYAzZWsjWnxFZ
uya1W24tQkduOUbIOE60l6sqFLW3ub/lR5rx7fnhZ7mpmxByHzQsFII/7rRplw7iD5bUItiR0uqu
srMOEO0vEjVGaL+LX7dPVFRWjFr15A7KAO1aDK8Z3t8bxYNOfhPWTmjoJ6oUtp58wZjRCHhyl2d+
wMTCFcMB5LmSiQgm3zr+zEq3UFewWDnj05acy8/iEMIJr95UDL89lFRfJ4AYrcx0B6DgHPp1YqZW
oGFk6xzQYx6ZqcjzjEZtpDWmMp4RpnfGDowuQJdd27J6piFlaelgimzDiyk8fVQoUyZ/7J7spB1a
AZg6enr/XjaEE+aex8Dz2XIIT6vEOyymnVcaUUx9AKb279NDVBtIKY+Li0k7L0iVVughoL1HXSAw
HE8Jv0z8tJiEX0rDoQiGGM7qwC7kxtMqGRMpnJ7JFdgMYp5XfFfof/85cxsP1iaLIT1dcRrmn9Do
NfUqJW4tRhkF0E2tIkF+UCbWte93mut/rSv9ImMwdtdvG/5U7dApHNQCFrAyN+rSM+VEWQnfHAtL
xGpIpTnsW00cYJ7pVNAs6Alb7dBvjbkP098Tgg26YkThRpS9IduzBPz/IqibfTcpki1ZKT/rA7XK
nOcGSfnskv5awN/1CRSJpY9vAGAIGEZLVl5DKJwn6YW2Hxy9Fr4QqQlyVEIdDAFXWTdBPs9bh13Y
OE2NNmVYP5QzPXcqGymSE/8Lmd7ySyIjQmdV2mGloEM3VrfYDFrTRb1jKUvKw9X9yT/Qly6r0a+I
lup7yOz11nvd+R/eqy4LyiWh40e/YgnfJchdb/ZU49Hw0/056pLFOaT8+nPv0503QjgHCqGDoQ97
cfRjiPsiL84g+yf4DT/dmXpb+YuCf0Easo66xw46fIV1YL1acxFkItw5j4y/t+uG4cUTzLzkmw8z
idSb6rm0z8XW9bneYc0Ytpn0dnA2PIPWvldumCNNaJCrPNTKg6vR4mUDMLw4j0BH6L1Fd/Aa0puq
qa9RHCU4f774ufWgtN4txxJmSR69QhvVVaWmnO7qigE0c6tUem+Z8SJNJH7ViOYFf3Cok/OVNYKB
xVKqM3l1TE+SytXtS9UFFOIVBsugiAK9vuemnBm5VdqfQh9jwgVJo1V63ZASHQIXBngM0cq9Mt5G
yKPVlZRaVZJWJrfyEuioBPnWvlhgVJCMpZG7Qwk3jSQggyvG7tXYQVq0U3ayBbKdu87X+q6Z8UEJ
i+kGYoPHts/aRf6P0w1+LrpKU0+oJz4wFPI9ouwGyhuFgHStiw80mvN3gvxQKF1ygWVQJm/3B6cA
3ULPB0NoJz/9tOMuJN9Ykt//vSE5F5tet50Qq9t3VmmJL7VnGBWhkpbCSS3OPfXOZwol20QsEX8e
NCt4QOQ7EsAB1ADmR4sDLQ6iz8gD+6ykR1sOlqPfthoXk0JRpA+PBDkFt3T6WWP9QQR9SNc5zN9q
DO08unuFZqi94agmlOf4Jq0x5/7agJiCjBa+njXA7wdVEVAKA04nuQylL0hZKjthl6VItU+Fn95r
5Rkda7TWFPxPlWNUO+XGEVLkR3YAw4g6LnRxoVlB76DPvH/DlLdH3uo7ZdybrfX2JXJfwK956iRA
1jMNqFn7CVEBDbfE3qBYBthwXDqcGFFhYt6SiazuREQIDS6vjollqkz4s3qK6Xt0L/4xSfRoDRfy
cFrNjYqk0gLM0hslKgjjKpP9ejjQndJrG57IxvcQg/C3QWwOw6VFkS2TW6flTy9xyL5F1xRnbcL0
4YkYh13Eaj8s6TjOYt/evBznXfRKu05jNKrYumecJzQ3M49qxL/m4KwxuD+P7OA7yb4Stt4+5Utp
wTJ/1CiK1RyA0KFb4jRFbVmjOjhOFlK4K6As6T9L5kLOEB79DnMnX5D/D57Gar6Qrkghcg2Z9Zn/
Ro+wH46r2/8msxNvqTZwOkF3i2NFCS7veBRV+g694qABTVbYmS6W1VDU2pD09Ahs71U6h2pajqw7
0cbShBCp0xGXBdTL7r4mhSBXc5CTVKMVkwQ4GeiKbk2GIcOYSo+qH5Baa9K2qeNdue4p05dncZt7
4/ymptwaFWxnowvs7LX5v06OawR6agINELXD7kMGqLijPsVje/Ti9CCS41pFw/7EGkH0PTN3FX9O
cA2wYCfyRQY2KbnXnvnhDwNUoPQQ6nJTuYETU72k9oMB6K6T/S6rTYeDMymynswF8o1Vv1iVxdyj
0nd9UDAwZzWDIXHJ/PApGAdg+VgQ1VzoC6mEfsUGT9xAd2Nq/Gbfr04qxOf/Lxu8ydzQ+UbR6NkP
S1hH1WXruytH0tbnstT5jLchifa7s7pNcoS4JCYQKfq+PkB6Z89J8BLxJQ61DAmGGltZYCUBvpON
n0LPMWNEQW5DhO8Sp7xxfip5a/ZOc1ppBsE1NDIAZ4AvzjmJuCpldvrzOhtJGx+mh3nXDxk42ROe
07xFu+GU9Cl4RR/lFzRfAEw1f8ilTL24G0IRpCQ1wH4AeqwUyUH5PrQdUL/eRI/DtovLj7IUWDgG
6NFJOmpjiHzHsCmLDJy8gzNjbvnLi8DyBqYZajE3Cmdf9JR1hRQdonPd8UYd/OgBuyUl8gQyMwmn
PDVmJoJX/MdpWb6qMWB8idEZUywCZueqqspJGIFJBHlu6Cpxuc5YF5F16CUs6dZLnqIq1VoOtZ0z
8Tcc6YXDBRmV6ytXWAJybVevALPuAQ/XCNid2UY/KBZR1A6wJDWikmuw1cIbXluuEzp5qc1QGhU3
A864rs5qOOWTdbZp+7Cwp5vLpnKUwgaK2vQBozWHPP8eTOyuUHB5XOhUuzs3IAanRjmWDYsaHkMX
WjXOykoPH9VJxlV+5yAj+bvC7kRTIGNo8SiYitAgRfzBKEq3BkugkgKSXotTuFqyBvHDpPjZ34VV
a/zEFHCNIsIgxWzs566tpwwUdANSddqOlZFLjCAZDDqKyBEVynWcjaHIOuyJvirde1SVyL4HjDD/
+XU0FIbrzOUrJFZNjLw9tEnMtOKcIuW1BKl0x7fnfSm5dSXbjrFurdew6skBYCam5zOm7FpYFvhs
FtNlN5wgzjZHoERvmobNRgzsR7fqwMxpf8/wVLWPirMMceRSA51TiyL02I2V/xuFC2HuayT1nVbp
/e0oat9A4EvS5+Q3AcuhtcpABmPehVXhnu6XVzkC//JahJnhcEapayznVwmfwfHMiybpGCuQFppA
gjiUJElzLN3T/8o99tud9UzK/j/I/NBCnXlqTIE9/QpOXETloI75qcA7O5RFikwnJKPn35SnU1MF
/lQNttS64+IW9jBaTQq15cqR/M79jEXqaaBcYAWua01b2AcmCKe53o7xsF2DhEZZfVrHz5ja/fzR
VGP7nDE6sNi021CkWznrJ5UAIVDRRM9SvafPl9nMH6Yg2j/VWftfHrLnKuZECkomezGhkIGKOSzH
r9fV8hHcw+ZN685QVe7Zc0A2wrwo/T1NqxFDlZBLxQ5iQNp+lf3usImOB643CvNetLOvY/tnzZQi
l4gSqEykrX8oN+LDjmd+a6DIY7CKsAmJ3Nl+6ZrjEgOq16fc3T6quvmEmRO0F3xsXwRyQdVyHsRD
MHgpCNu0hGadA5nnyvGINLFwKbc8B/h+XYDy1eE1LDeI7/DzNHuGCz61yJtZlbgMSaTrmeGkWVTQ
W7CMD86cEIjXZzUu8gHAxPNpOlvWBSBSnSMeNOR3fbOzErQN85fRtlcAX5bcMiIVdwZPL9bOPyDy
eF0RKtpNs+i/gRGYvJL9MwFaTxldX595VrvWvEZ7Jql54dKY2VUgZKrUhyekm+WbBljUB4mLp5zu
0oyt0EWAj+vpFeKNsyaIGxnbzI0muxhLhWFXg7HdJzsUa4fc74TIkLE14/5onD1RCeusgKC/QP3a
xNIAmPnqIwz5iizovXB+NeDibMXU/TzMuvApkXa7Xm6lbQ5R7aLfC97eTKho6KCAofbV2AIyw9m5
psGo+kLkLQkaLSQ9X4hLcc+r7GgGt9CenwazoASPhx4+a7H/4sOpu2Tb2XigigYZMThqZJgzYdQ7
CVKYddzV/WulBEllvCwCOGXtbMUQgvUPKRL7/+4PHyMA0mveDsmKZd2sNKCsuy7bdXAzifGXRoXg
M+4FHhmwRrfry24Z7PLZxTXbSbpjTCxShIQs2FyxPM+b2rQ43atFeV4qCdoZ3PNT646C4SCXUZqZ
h6q2Un5hwuHOKrGaw/G/z4uYcrLeSc/CiBeSONbyHx+NtYS4VdOL5j0ZYnxMRnCVVpmvKcw4/NES
JWS2gvxEPjUAUOHtr0BmEbsECzfdkiPPNaTnuFSfIP4PAvguTBOd+7724ZpYlF7FRk4EJrAQKWn+
vRxoAK/0eqX6SQhJN2+Xw0JZCZfMdgUjbZ9J5aKaQF25XmN6Rd+z3RtninEURDcJ7rzH28jXa1r/
wx5M/l5IRrwBEY6IlO/6/MkgHLDyvpO1KW/ZWAFsdCaedqeHwaXPumCop2koPNF3Eli0xlbJkD1V
n1AHLwot4w/ydAHC1qjorJe98+TE1baKtq4OUGgiGQGXbDNn8nP6B7nu3v9ixDBmXHaLVOUTO7G6
+faDuRW60FMDCmUUJyNEMm8TRinVbx8D9Ef/z/VU/q4tM3czB4UPxJ2Mb4ACYQudg7wExxe3X8Z3
5gt+GFXRdFG/0n68fl1wpHpn95O6uW4gxi+ChEiQRVr8//HdTXw8pZuQGV9v40SezYEk/PhopG5R
3bEJ9eMy6WgtHMQ/WikzsLJjuNUiCAfkwrxQQ08wC19t0wQyXs3hKlGQo9Qn3HSrKKnynePDQtyA
zA72doGXsjM0mefJSyGfY64U+h5U21zibfepmBjPuRMMG9TGHz1h1gvhBvca/uAiMmdj0xjaGp09
P/5eyIeCBFGPduPR68Vr4+s7AVtA7EuNNvs0vyjvt44T8ovD6xw1XdB+pK6Q6s3A5NIycttGedxD
UQk8hREaCPo5OzPJC36/7lQF3YTw2xd1YVLhqWrfWtHhphw3pSYUCd29iw86qWCYEvb1lYpYwi9I
Nqe66+9YF6PKyDIjmp//4GYX0GXWm3Oh1GY8nvXvSVdVoRpSknoJTMcXwK7cmSGFNNv8f6iPjCTD
pgOWHXOvepgSb7FM/eu/WRoYOwBsnkW+pCl+bu5h0zkLx1vgY62WZbub6CTKXWi4enB1/L3Lm0ap
WClsNPvYUI9cW/C3rfyH0RrYUcB7GCi3GYfumIuNuN9GLZi2CG2IibyxiuNHvS/9cevYjK9aktSy
iN6y2OtcVcHLK1ervG3FLdvQrbyyoMxn5QayLrVeMKnZhPMp/vGhICM81/P4C05emcqU/HpYdVrg
w//ybezoD93KBUIZQn+M2Twy0ndxoVa64KbHHe3B+L/+jPOZd3dBSoPYsobKmFME/s3DzzpL6+St
cNVPsEbLrZA4gHZREnRX33KJtx7zYE/bqFWcirglgBMdHwCMgHOcUL/euHldYbwej5Yz9fs00cIV
FJrV9H6ulnihH8SkeJSeeflEyYAoBt2xUH84XQzDkquVPMRMSo6Mk7+0UoDt3bKgoiAFNxjxbEjz
2l7IZJuxK1h8KAHBpio1dEW18sCJFPEWnRUIZUGK3VCaA7YSpmax5NVvsMRP5lcEgXJo40JBTf0/
O6fKKv9FUMCxWcDHd45BJPYcLc55IUGgBZAzWRs4hwqGp8XVefYAbbOWKLQ7G60Hnp10F8UdAVT6
BvS3kEJGADJiqAvrIk9s5MMVwjadM3+rspJgr1u5TnQyhmI9AtL1uandw67BmPG8yqBpP4NIFFkJ
e6VX8NFubm8UvpfiYwPlIXw2gPpXdiinsaSd8i5agRme7w9K5FeKpPVPGiCXZ/82jpr3aBC22yAa
InjwMkGvQsXdDgPcJ2oW6TvbUxmgGoCWzh3oZVcCjqay3lRqOo7w5XQimYUTcUszzm0dFqa5ix0P
dQZnrsOrk86Rbe/1X4LKNPXF3QCreuAR7N9tSji6ua7IIsMC2BK69CyZNHEXGJYCvjGgG/m0giY+
8MidOPEP9GnIdn1E1/QF+vWCILBIikkQ3TrnHvLdmtzKzQ3HTqhUG+nDNCEZ5asAr0qWv+tqIZxf
kG9kyNkoLRwUbp4H4gyA/0HDqtzcWG3aVQn5l9i4RH+7TN0jy9oZFZ8ijTsYtRKHWPY5KCQ3OGvn
mnsXIlWPZgYxYHtFKhYYaOsrE3YWXacL4mpo4D5u+2y1/8ZBlYAE2cQvn+66ihw/OwMzbrnmCFI2
PZqYDpQoki5RAMAirtjcjlpAFYBO6ByOdJDaowUmTLwmR4QmD3/h6Eh94R2ZBGy3HGoKAH/C7BAm
gXrBBaUTEEF04UQjMTNQvWiHeQmkFbJi20VYVJU6jxQ5E4SoPTp8DzLGPJEqzAK4k31oko+Yc38w
43vAG8dnzP/5M30reXOya2nu7sdij1Wtn7n+6ad7Om+EcthEe16NkduZfOlJiWuErKRYkkoF/8Dr
Y/HFYikH5UWpNVjunlMSQP+LIQSGyb1yGWU9OOanKom1J/IrMs92jJQCshrCuABydPRWGVd4cA1u
Ao5TXOfE5KZ/ah8NeZ57wova7DABE0NundSz8ieZZEocSUhK/pz0qRvUeRLjDrycuT67qp2AM2ba
zVNrXuvNwSAEeC4iyW8ee3sYiRAltF9jSovgbR5vR2MJ4MVf7jzAz9pKW9HaRwo3DepEUWYArfUY
91ggCp0mFultEk7NRvDa8zGCtJ8lKwixqD7Z6k3+6+F7JYBHCv8bWhOpJCapf+wWuFX3iDhHd4e/
ere/oKqzlDLeHLi7nXtXnqyuaF1LGELioo8bhXbI/hX/p7DPZSxnHHYvd+tIx/LY5/EzyRyKptJL
SdaMMUKSQ9MReqKExCBLZ96KQNBo+vLrdnKqHFE3jNThUfpnwIm2CoYvdTTnVXJJyoSGwA8/llof
MSgS0EmIDRhFgzQfVZa5t98W+jRTvAMArD4LwZy34j1mvWdrxUCpYVTRHhbbiDLzq70gyODPAmHF
molgx1aZspbAz1tIccKIsZg4fzLsAi9TIkb7wrYMdAm0yx5J9qTWRvWAt8UVvVgT0o57qzuACtNX
YOfUhF/9t7//DWZ1AxG++/Zks51mYVJ88LX5i7nE0PoBlc2Fv8KEBJPgIsl3BDotuOPs868IdT3o
d9tXlzRaW4DZK6bo/5RuULScp/vF4G6pZG+9fVjw/CxQoeRYELRdgGvsIqBcO9doRuKBoeiuktp+
zwYUPYcPViCCUfy6YCcccnrDmVp2Y4XkdDYF88rstMAZddGQ+oQZp1qGDSHghTsgAjlOxY+OFVS1
7z+TMTvgdU6bnBhnAJlo0UEVQ7+4wDNKsAaXAwhnxpdolzigSig7FbDT88CU95UNCFfVwx9kXWHP
jLRh7scx/60mK62VO+Dey2KbLBKHUKZr33gIKKlutnhNdL9bEjAbANvTRJL54wuU1e39lIx3t+9M
uVsSveSiAQbCgTvMxtd7y+hCa4k2AQE+wyeowZcvBa2f7DjTg4j0bmy1jn9IBF6UCYuz0ij1CS5d
lP8RmecgblzRLSRxCgiGLzUAD1XHkha8UkXvptDovHnzcpn5ctqBoiewNJxtRQOl8hXgiTAsAPCY
IdRAARy00PUeZ2z1GiIRi/qZpXVYf+TEA5CwqGKPz6iM+V0WgG8t2WK6fpR8U2TV5dKPu/zj57eN
fxC8ZNGsQe532aRdiW+PVIhsy/3aIoj5b4F2KyJ+mw1jjHdyEkioDCRByLoMc+EZi4BL3PYB+90p
1hkrZ5kiBeWM3SE4XQqEktgC8SuxXT+9fCeMOegRFifMSf+WWtqkOPfKhWowYHjvg8cjmshiPl8b
D9h+/FeImHgvusk3KtLkmx5xDnwlrbGouV84oZrZO1pye+TQfe755XvKO5prkD0G6LUR9HUZt7hI
XfbvAK9wRMKtaDVLGNdBvRvxZT8a/AfdbqvlQTv5hkCXWdEfmUO2u0QUhm964Y3YkT/Zy+9UQIXZ
ngAzBUJ/sXcTnP6+bdZW8FjHwdKAkJjOQ2veR92oIQXiQ8ynGfMBSyFEOEmnkrfiGZU6S9QSDsUm
wIk9/t44LQhu+D1r/8iCCI1KUhOJbo9TGJTtDa12Us6B70QhLxdy0wU8wKaZR3g5qRkoQCBiiykM
9wkVypbnoDczVsFHGqDGcDRns9qn+NiRZjhWrPskxdg5olblCgRub8JvuTMOM04HaxTHwXxR4dR8
x0J3hD8uxBwbK6VqoaK3kWrZI9C86Yr7p+cwHuE3x8wchhsdjH51PXfh0uss1S6Pjbku0qccyBVN
qoXpwN8OMK3qTQPcpDcZFeF0dyXNewsmETiPx1U4X7BQy7mmCp8JUeQROOdkegYKlFzh3I6ugdkD
XbzOVisvkoSuOwXjcAGlKprOqwmTLtlDJI0F5wBV529h87GeoyE/TNg1dzC1P+bBklD47n0dRxUe
K8IiOtdM/VTsSmepcOKtxkL00mKvBI50JcmdzMc7uPQD82u5qN9GtCpOwgq0sE8WtRC+OXwhQq+J
sgN+QFAU7P8yWwIGbvL3UUb3vBegy3dGL6RC3O+tE7wgwr1xXftIkEqj0uyLfpH6EU1KXoLXxBRh
rzo+Iiss28B+5xKXDwlf3NLRU+XgUKYP0dcxgX9QWNFc/IvSB0qXesjG4g8I97k3iFA86wIOR0KV
CVeqh+Baoj5Sli5lhdJbYApdxPDVLm6YzhL7DfKZkzNOZa9VWQfxn3qeIe1v2yOOdJG+Wk64yetu
j1jfUzIsmzxYt/aIRT1EyKe21fOcZilR+DMkekW3RLw6D1c/mZUjaDZGAaoJyaOF+j2NUPeLEsba
GvRuEX6svfyHMlIj2Zf4NFCA6xGuAZRzZTeQLMmhpSFTwBqe0ohSQjAW3kfk/vhjkChgs+q9Io7O
7vev7L85HxDmJ54kzvjSk1Clu0Uvhw3OAgREttRQTn73obFc0bMcZjBO3MD7q4Sn3zGiR4byrvdH
FyLTOGxvkjPdHt/baTWvazVzqMFdd9gRN9zrrsawqwKx8kr639/wZhLatEvhQHJenELXonBu8AXA
aXfsKTvUKmxem9Z16GhUNYATG5iOJOqj6BT/7OUrYFH8inAR/5t/cfJABI1ArMarmzRz3Xeg3+kj
7UwxYAZg3cxIfAPDV+R6pQ9TfUvCywdd9FhWd/vuHHGrksMSOEqs9+zpzg145PCb7l1yWNYFjlmv
C2aLwAJs05fYWypUxhD9S2GMS6/WNR/co+Ptqik5widmLxou6waMoZswYOqi3e4FqjWoKa3ezd/v
tzf+VZmMXld7UATkmr41HbNHUaJkkp7dVoD0NhtouV6KkF2rb/E+TWabUE2WbMCKACe7A5r3RZeK
VmDJGhAOcPgicaO0hQPUkheyRYupMMCr3vxOsShO6aJbaL9XkQqJ0+tlf+DFT0MnK4QmRoRyfUvS
QImC2rJKvuEf65N9CREM6VyIPy73tRcvI+bUF9gtGLXcZy2QlaG5Us6S0oFrhfS4nMFASoEQbAZx
Owqg6/betXYHvKHXqbw4ADIqsNNug/TzBG0XNo8+2gDAQPwVB9L9b/8YKWVOIHsKWvMHzxpak28A
VniYPMuoryMLBUIWy4rQz62DTjcSja+zJyuOVz7sMe5TT/SnuAFPwp3GpCAEzF22EBVu0AWxs/yE
QZlppCpxRhZBj1uj0xTOzBsJxQwwnH2J7PdcwMwDUPeK/7exlDwCkP2DUp3H2P56Gb5HNGIZPQM/
NJwGIsswZ1mBmq224WDkwbA6ubVqFU9dnQzplPkQMeLVW8hb09bhel9Yi+9qLaeELWEwI6FUsrRa
oJMdpsXxC8JKxozA9DaIWXEjn/Iayd7S0msyu30XrdhyshWdgUARdRLUZ5izYolKL+ts9iaDiFw6
6wCzrhFDa1keixdyAUi0Mk+w+2MQgbVmjckqXcTKFyrxAFF76kafp6PhfytWCI7vrZ764KldE8c/
uEaVMhpSNFK48Kopj8PX+4aPfPiRUMsMFA6zPYfKKjne7p0YjbMoq7v1G/NVIOp3sQ7X4QPN1teq
AEhmH5ZhVV3D0xFwlC+NgN7K16k1+whs3buuo6w3SPxgB61NncS71YBxAr3/b0Pw+RfjaYGQrJFX
ZiJAxOJwkzI61TlXUomBk2MMAwmunfg2GrqtcmM2EULsRqn03tnA/xldaq1jd6WR2fY8cpasFwBb
oP8BRPV51nhgk9BgUD9YtkwdWhXGFzE6/eCma4JEKw6udGPDRBhS1j+28CG1S4qMjLfZuhLyd9dU
C3YbGYtkolbnta/ag8kHb/TmC+bxUoOWRXP9hZ9oKfqY913H+3bvz69F2W6oQgnJM0N5WIMjSfD9
lM2NhqAitrlAhwvUEBzr1VuuREbjZd7S680nvaUrst45gfAl/1TH3O4IZsYb0cBtglMwDiZR8BpN
vykoRo2J43J4w6EYtGCkYcNX6DW1HfYVTFnJERjib7R2pYBNniXFFmPImkY3mjcVslyzi6ld07/i
vphpi8T7uCvVYyo3+Hii9Vgk+tGEp/VF/2VZXV24+uLKcBsxkR84ZFPNhZYAWnOn35HE0zBW1cwS
PNztGZqwzA8Lp4sXpjF7yK7Pm9vHiiuDqLZYeb0szfQTBTgTA9C7LayQp3zcrSFldON7A0koC9Ma
s5E+Dnyft5ZAb+OKBFUJn4de8yh92NEFYdYH4Nrf46f5rWGxU5F56UfUWGXKTXDbgGvQ2CI7Z0Ui
Qf3Va0cVMeP10Tpzcs+PYcPMbmSsMQrT7XpvrcK5FIffscns741TD6ouwJAektoCD2jcu+olmxdH
3F2aaV+MzcbWaJlOfgNdoevEKYYzKkLSaMLBz6y3W/WNBsWFXpBCWri1QVGlLbs5wkFvE3AZdJ+h
e6mgpgtbbS7ONyyc89M7MXjuyCkfIpHo18HQaiDe3FLfXoKfgitX9AuXDxGZ7jyihr/RHLh+MIEg
zj9WZ2Zhv+F2aEqirm+Y9FPm5WzeEeXMB/tB4WcnofzcB8H4praH76glW99aVGKft+N+TgQDcOgt
1nv44HtHuDQ3Yzf3JX0ghU0+O9DwIrz+PY+hqTfspoL7yTxEFKNJNSzr6sKc40iQNoLFWAkDCZ7i
r0qdlhpkEGCzGzpTHgWrRN9G7K3bYZJXiq89NkqFW/sHNgSQDMPi5iuV4TrhmyGRy5/J+khSTMDu
2ke5fbpMguP3+s3J3psIkRhvESlbb1HaHwKbhnUmnslgd9Q3FjK9NFmSN/2GxvXpoT4iAYO9wJXw
0vI/3YjEMzM745lhyMN6s0gLkmF7e640IHRFdsCPmqP4R1TCe44Aw3wAw3ltEVtZrx6Mik5O086n
Fz4pyllcbx9iIteVf64ILmdqr9eMTRlfw78eeU/Hi5n1WFDtpooQbRNT7/pUTWPMBcxETOmnds74
OzMSfcbIlcP1ea3jlLuIQgsjyYIIotOfwN5A+RP9u3hvFSFcJCpd+eNx6sy5IH7Suq2OLpuucVQI
cifnIS83JkdpLvoSN+DznoDxP6g8bOD8WXibl7yd3oIF7Q6S2Odi2pS7eA1fB+OYL0Rb80O6aQXS
QVVvAdXIoMwdpI0UHe5y4JDol6OmQuYN7nDG77IbLWB1UaP4K+FjZmlbeZGRFJGZzm0F82X/Q9kn
xrRPSCDenJ2XHBqDWxR81mbP+FNfn2Noe0iyueJKy98cVHAcjQSWNq5vSRieuRSkrlKOjtYZhvuQ
e8M8aOKMMBOkmQoj7Uqj2pFA43cJy4lJJhnA2ECD4EKdXtF6Fzpf0WJyhVCrts+3H5pacC+7iGIp
WTIEUmYEuTWvrK4PwVOBcjUsM8w/K9q79LD0TfxAGecy9XcGrLe1KquZspyIHOvGTSerNC8HShSU
D2jvTznq4ePgUagANt6D6NAA2A78Rnk7mymE8DnIFCArNXKBP1iQv5lMGbBmFX3wLdBsj0aRtPSd
IjM0QI+XP7VdXS4Ab7i85kkQM97jeMjJ7Xqca8bmmC5sEHFZg1JPfsQ04p4G9OIy5/qOTzqaVJW0
PoXGxPKNMUWOWkb8Iu8xC3/aSus0/b3CHqQYdQNaDZu43jaVY3UC83idG2YARMIZhFpy3eFFNb7s
0vywhqPMHqeei7gKOcXtxOp5NWUlaPUz29wuoFWFu+a1CMiLXec5nw86dub+t9ulI3FLglY9Tgk+
9ukyer/zRtcaD+xWznygVl1lAuxWLbtnyCf0cUV+Ulj7w35diP9d7Nnc8Ltjpbt2SLh+bmoOG9SB
rfP0OTXq8VB8tHbUtdoQiaAQoc03JfOR7kRlTBZrwxW7O2enwHeLnSxhfzQiH/vhjwtQFnF1DCkt
2gOujkgjEEGmowyoUZUtydwA0rH7kM29pPWusHW9uxSWP6RFCaVHcixBV1R4McHZhvzrmUBbQdx8
3QVA+lzqJvyWx4ndXNmzmncAUFO4X0TKk1qYzL7euFE6f8RRXm++E4lziOCbzWG+ELVzAVNanzgq
R9/rsrThJRCZR5dtnG15JfnXDUZKyZaz3pCUqCELfAVoLH1+wqiaJnWxZ0LzeM06ofa5TjhzHC/O
mVwjADwI0brCUoj3djPL8UwkfpRcbCmib8EJ5xfxfwY4ml9NS9lEQ30w/IAFgWS5PY9MY6zL9ZYs
6WoTrWE8rk6lWQMVPBo8EKQPGacjYuVHaFXBOz48OYv9jmht7zyhtNYj7RfQ/E/NiI768dM06wtu
zPxHUDMaSJbo24iQRJins99Ycn07+2N5d8lz9j1v8wvQRliPgr3EltJe1vp5d5laTR6Z6rvY8JMP
sfIMNDBFwuxkDYDYO1emscNQ8yUqpeiSg74fBBUHgXd2479Jpdq1b5oH+/y/++TXbUaN89N+0nMg
SITkLsdZxpQXIcb1dlML/tOpu8QzxmChLJ+j1vdNF0DvFn4VQ0H0+W34PSTWgzhSfSdmaL7fcY1A
DQDK+C+8qeeBguztznDatfexIsNiWyuwaYhP0RX3vWHmQXGdw27RgC5vzmOuzkWBnwSOx/q80S55
DKmubtURgBZhRMVujnkIQYD6ZboNo/qMrGJGeIENU0fQXfySxKfZuSspVlIBeSm3AZ1mQF4KU4hs
7BGpPZ1FPuFK6rtSMqXhCU6bwvU1729pI816t3cLrWBHpkOjAEFDsKqGJdRJzAw1e55PDPOcvIkX
FUg8UhIrikGObhOTKnMZe2prD/8pGd+Trr4mJEszQJSnGZ4oJNfJJalMVqFpclqxdnpNnN7lfn9o
zwd6CzIQULYxeJf/qhdIbAVZyUJBF2NjrbukStRzaPqf0cv4MUW4fUpPljQE7CgRplzzFNAkrd4n
N5S7knUAKoyeTZ/10kmqnHjnj/1cvVv5xYih5pi6Z8/ikSGZK4AjtGiisWDtszD1w0qMgADibbzF
UQUZydsBtBx1NXwh5cDEhjUChXugeoUs8ct0Kjrkn6YlN2QgyM7R6gGuCYZrjjaCOwM8jC6D/NsP
Qz/QG8JKdfHk1gzuniwZkDGgLn2iMwU60TR5/fSayc4qiO5N49gnATTRBvLlqfxQVgkiMgQUZf86
5TWAj3W5etweW+D++0iNFgjI+g+BBpWA8NvuQlJMPGRg+5BXuNEL4hiezBJvEjn/h/wTyCx9mRdM
wGNPpoRqS8IPNqmkQc4zul5J2qICVbJ1tJBKOh1ttCoHL6nIKjxYaBakcb81JPvjThFFsJwipmWT
PQEMzWEWHNBN0NE/MFWv+4GP6c5wF27ObSalJom40voisNw5x7ldjFF9YZxpw/T82I9dwAzgPSFS
ByiLuc4IxOX3PJ6KhdM5+Cw1j+QvtRkXNiv/YLbxtbSITU2yru3ufk3cEZ7JWfunwBLI2ImYk1ZB
is0IKaqavqBJ6N48j33P28llIcYflVkSqlgNRVeo30vQ7Khlpht1cZsdPissdr3aycx3Xb3AfN6i
YZYMHcI/vmvC2/hQHdz3uM+YglbYKoFImKsVSJR+oOYTLXuJYyqaTAHyav808yaZ5ZSvK6mtgZTM
rlU7hEsEwRla7D0AIPl5iCj78GVTGP4IMYy0XCwMN+ZqokRCLVy97mySF099Z6TZa/cu9QfBnkgS
zkcvXPz/lauiC1XM4/Ceg69bX7O7gHRFW7kzjLmyrPX4jUVcVQmtHco6kvCdrx0SIgBBUfvJbIpA
VuTHUCcphLtNsBSBb3bygJsUZFPWC0TUnfyfsA0L9UwosqbL4ZjWDTQvUgYJtttpbnvy8WeRdgPH
yIigigOYcn7pIPthFeRAt0ResnR2bjl5gQwkYKKUXX4y1DHHxu5ZKCzET1pOudRAWmoxkYii1ByZ
1y4R+GMCuTcj/D89b5B1UaPx2yJo5qrO+lNGoYXAoBKwssLOAeQoRj9974NDJMWny2iMFcyUCtpi
FlTYGnhZNKDJ7pYSJ1yUyvJK31M/b7AtgiQPMHh081J8gpcZgqKTVOw3xW48yqxZJfki0h5bZJyl
kmstb36M9m0KD3DOQQvvMFS0J2SHey5D0zv3dWHH8sl3x12W7nw8iAU8MHQvyqHku3NXyvt5A1z2
2ltTx+Do2jBVJeTS56hvB8OQwvolNRMB34F7pkmoSCfuNVoSY0QtycDr51EPBxDAWwTCveQIIAma
lT6y0+/gY9z8RMcN0vIBfVZshpQUJdrA7Ae+x7kWaXghrBCszZNXfZl2/6Ttv5vJFemTyrTaM8qe
mYzHoD4atbSD4JFCAXrvBQVji9yXKVoMN/nNWizcQem0Y5M8twREcU46FuPE6Ql8JCbfmqZ53gBd
dVINUd1WEqN+LgW+t6JGVimZqSnniDiyq3nSxgNVQabbxrOKhcmleBHSf6Ehkh2jM0GxGse5MnxL
ZMyoJgD2FfXW8hhKeKnqkMQa4CwN9oEqo6I0Kr9Nh9IXVo7tn9uV18MrnarpRhaJGo64KMyObd1z
veNuFXSg0NpoOJdym/uuTm2WaA2S9yLQc3sKEkkGJChLyZjce0GAH4j7LvXO954iwbo2tnr9YAPr
WFJ4cFb/HhgrDVZ97ZekEs7Cyo4aUVouxhLYX3rji6hGr6MpXmGUamorGwx49ry9K3UCJHajkhRB
7Vw0RntBBF7Et+IvI7bQNW035VfWi9szgyqjrbbEkIcLrxxModkKTm36jKe6dB0cEJWV+kxIKwpP
dyHITW/HbeQYK0X9eddlTnh0Lg3O5SqCq0ct79FQD40obhl47Ql++aVWHpYbZVxfWId3zsN4EBll
PXwWKDfKTW7fdqP7/lMmapT9UJ9tgDfbIjmm6alNuN29nQKg/pZa1QuEPOPDG4vOHqZ8rzysIHLq
4X6g5Yaa0ussRQBIWAz1zxV6td5nvXAsAexlpFOaqvwGX1plo/Cd3zs2nVYw7pHEvPMdLnCPLsdW
Iczz4nk/7Db7WoLd6DNCFaZTHKkupMUmQJHQASSy27Amj2Iqi8Xet9BsyxTEmqTFaN6pW/oODmQP
YAbi8azA4cppWM4Q6ntzMmE1OPPPn9HzbqT9M14D+UzOmwivrKOIod0DX8hg16MeUHKzoBzwE86r
+QGCFSiCMvlDEou+jbi1vMwAhJcsdEh1XQfCP1tL/sfXD3FvU+f8nXcY3uT+9VjXfUjAa3CMMzal
Tjp1/CFEFhTJZiYP2BA7x7Lhhnt+z+H4lxaawtaJt82piCTLTqBpjo2M9o27eaQVH+tz9J3+qORq
0K4wSEOUIjo49P89aGGxY4cpbTjG4gxgjQFwH076FaggxGRwoZO6lRi0fTQ5k2hBIN9djjyAbYqX
NGy3XIWCampIgtmxbXG2Da08jNgoTJjN9CSZPvT4OQScXM6ks2NOE1LTwpXXnVJ0GcDwDM4YS+ia
+An54kn8HwpZtA85xySwwjlxVa7NJr6dF6rg3gqwTCAaQ1B4WHJG9/qzLygIoyTxrW3z8Betym3e
VKcvu8lOMCK5kgfK1SeZRSPIWre24h/gvEgqRmg5vc0zcRCKAtGWg9wTNYdi2TIwmu13Cg+0fCEA
gjQ/afWqQqQuEjTiXW9/t0G5VzcgEyblU4HZmAfH1DimEDcELl+7w9x5sH63AkbHo3cAL5V1wRCc
Q5powxttW76muiIpyd1JkXVzl/ElP0fNQifd7jHi+3n+59dzQR6AavI1qBnX3pD/hRis7nryy0JY
2X2mLls0BUoAlIOonB06Qz9gUK7r54uoME/dnfS3vhyyrOaee4jRq49trthJ+on10ukmRKvD+5Kq
0lUPHXpJ5dUJ0ynbFn9/izlzkZwlP5eS89SkeQb56GMJmK0q8qJosABniZj6OyFfROAFeTVMd5/x
bHbYXVwAnWZejnulARkKLitdIyuJWDcgGMo+OT186qHRhCZaB1+2ZlNtbtX4Qs39dbAHf2WsQPx0
xjwP5GMg30ROS3l6oBddq47ybxBYudlfDfIpmDwjdBTeylDPTI13ivRNg01djxFY9xIPJntTM7+u
UhsR0iL3l5msK54BjhBf+KNmKiqLiZ2pDblCHzlh/41K0buBskfh6YeXwP+q8AufV2bucUlcrYER
7X1BYVMrhQ9rFAnAbhNhLx8wgIHwBXqE1wzyR1E/Ugb6rf+AW/HM5aXYFKAaVzwi9ftKAAcmHBJu
HUFMK7XlbB0RKFDpGBnrPx/yjXCOShC8wDrea1TTSfyVR/a+wylyKJ9C7Hp3u6J5F7MA+eBgpQbI
/GQKaedzh1MV+QHlU6x28cFuEWljFyDz2ye60MLIFYwnOYAvt6V0HnRalTEKLRENUPtjaM328ZKR
+vLUtV6EbwNldOylTpJJy0v4RngMqxowHWux9qLOTVAsPevDqQJUWqv8zPVv6ER5L1fH6YdJmB+C
pOggoMh9Ua4/wm4EQw0W95+JnTsz5z7H0gPaaEkeWBZ8ll3x9D9aH0TP2Aghi8AukLJthfwt35o1
ytw3BRKSAEefqWUZwHvNuBvVHTLim4k4hMWKKiLuCQS7Iv1eXJUPBw2rIbNCt934ahYpI47jCYTE
8CO2rssvAqG8Xd3zkwmqmLkRu8afRfOfVP8JX8R5erZJq/DEQPT0h4kaUta86rkLNBG8IMpWI8tH
QZ+fDiz2RxOmwCOcA4rmLQkCPIXuDu1us6oSX6LFFD1Mu2OD7Dmr1Pq/wesJZ7iJHgTxt/RWnnGz
Fv2km0hRUrRF33VO1GVW65KEKrdeI7kinw7lsMjTPv3xdllhvhEY/5P17+ht6eKv47y5z+DHuZ6G
MTBwcAJfCzPcLM03jp/dFW+sLgUCxVr4zH6DluCSMSSoVp+vgaEO+tg888M9XNuF+cu9Z4xMfDJf
AwhgRcOZvqWYIpzTykrNlVE0z3Yu/rFl8zj70xTtCXEpBUyq1lObX4PF1myhpUBwNZSTe1KzXz03
lmfoqVGmZFPCBsKf6ajWlMXvIicqRszGSgnh8JqlNbZvjgDmUtpBRR8P3hJouuECEGsfU8BGWxXw
DP1p7ez6PAJ73l38KJx6hZU9LZR3swAj3ySSAn6mi7ls3UCrSFc0SUmavFsoUm34J3jj/nuT0JXL
FqXeqo1W9XJ9ku2kxv+ofD1wsvlcOwMn13YdMCqn+YpvkCl5Hw2gB6MsFHBdTnic3YWmW54h+HR9
I7w6XND8QcsHk0qw/EbwKtG7liFG+yUi36iXtLAWLdmeuXjDb3LkJebdMHsWlHgs/q9pdBskej8T
erkVE88ykk0vupEKNpgfB/6k7AI6VhlPgcysgH6TlAqLh+0Ih2WRFwH9XzQiugkFNwc5x8hAFHyP
7Kl2/SAUmDPzMkfBEMMXe1meVtruHWcU7vccIHHK2XONyJc3YI3+FRquT4evAVSjtNBviQCQ7S5/
CMKivCO4CY5cNGqd6yiwg3CricPHrQlvG3L8DtUNhNnKLlGumpu8wrntbf5zj0Yj+74DT06OQs3p
wsk47ysGEqfvHioXKcQGrd2JnkXYeVdl0xR7nY6peWWBX5OEbw5stzWMNsc9VTmk1uuiroKCCxgt
WKjMDMA2z6CpAPis1+IQrv5s5jCYW2ZWNHjfrQFzBJwhjr89he+jy1QVnk7ap/T7NV7jUNTO3B/u
Lk4n3+bQezSMQtIG0brqTEmGB/bAJbJpL/H23Tzi/e3l/xTB9rrIyBQuYwOIAJzf0pqUiewiCqbr
qhQhDKSmopgk/ym99f12CAzvSwf8Cv0qbSbW5DCIHrDOVHmohiqlUpWoSi/KNErHcxpzRVNt1vCU
CBzu+3efDr/SggYKLH2LfzZ+gfy/XeEULdapuzhix5RlTmn3mb8RqYP4gbMtepio3AbQfDcwpAKg
HckwEn7swjdCXY6zVp3As+gclXtYGT0akuamo+taLA4CdnHw88kkxfHIq4j/lPVSCY5BrBRBHAVm
wBxombD5UDjOvDeRL+FuQzRqW/6raGY2ZGrMS0tu6gC3Xji5kciMDfpYHC72yjF21MCxUhKRJiF0
IJAN1YxkViDX/KgrZxvRewl+Dvl9a0uhsZxo8iw0W6RI840eNs1smd6qHaQY6UnztTxX0GkwqGQB
kjvJfpqq+ncrn03+Z2sIaWYbY1+6rvI0QbomDZSipb+rXEm/opuMOwENq/ToxGi0zG8pFNdd09lz
zSkJOAA7OSHxjimSrQ+ukz/1sSli68aAfdeshw9r4xZaIoVO8y4t3ubQFpxSCfCBhyIkH38y/Eul
TmvZpPKZIkCDHltw+D+1aVtnsbdfek/veZebbg5s64XafOS4J4lD6wII9qcck1mbNWvMKU4O4dd+
bMcSUHCZfGWLPoYyRwvba65GCyqXk73c+QoPk69qumGxbvTG4+ESzc75kSDZoeINVZel4dQJjgFG
x/SxayubCSgpLrSaERTGB5R6VyWC/h1AP5ayo96iconPBd8VFwR0T8At30yq7vId0pP9tOzUqgDn
vaskI2Mearnwz+EE+g9W//BHPdkaBkj5YGHW8Np/DuY+M3tII/JZH+5Tw/S3QdhEK6nbhiFXC7Wy
tg7COuHjfMwizXNtgQ5LgN92iPqRhxGXZhXtgEdl9ELym8GRj8z/7T4hYByo9atvvJDIOrsskzjD
DCO+FacZ2Zr2TYIg+Ec1lf5BgGOPVEJH4/sZAFv5twCfdM3EvtXBifrQZMDq9sLwvoauGhAKu1fX
G3RjPqPRjC4Jb06gsOOZqIPdsmbdHXRAkNCxQyaQwpbWpNv1WGAjv/loVDWkQVNv0IGEbc/M1kxB
adiDQITb+DFG6+rzq57Hub7BnBbevzPr9tw8mI9/Aty1+nyaRk2HP/klgantHS9ygsAXaY5+InbH
HeasKaHn/xmPIbfNggaFhoLztl8QhDuEN7BAKEhu4kwYxHxrrU80Uj2czfZequD0u5xXtD7Idnly
Cl4qQqQaWQJpy46GBFBISb8Z1WpTi349evZPRjuD2JJYNsohj/Yu2o1qR5tSMo069IA3531LRR4R
zpYdGRNq/U5cRR7ZpBVHOj0i9I5ZG6KEE2B6M1+jY1NyuYPL4p2ir5Yquyse5Dwcc+8Mr+T49GWL
1lCFC3LT9EpJV0fnSQ8jYmTxQM/rzoWpFnrfWmvF5jmgkoVJTKJb9RLP0sgNfZVO7e9j5wcbYoMD
rK4Slum7DcI712m14C2z3J9omquKXZq7LyEHHZ9UOQ3TAJ4qnLBiem+kwmQMzdk07CVlYuPAdL4h
0n0IYC8quJlDDyqKOQ/oYVgoiwt5Cg/df5Vno2AW+JTz9qgXOXI59BZgEwGNyYVOb6EOZK9bM3+x
ydvv0KgZDqyTV8TMS/k68mHgbBAiX8YalISZ6pT6pHkvoGbcGJuHutf6cuL6NtPwAS5m0SuG5epW
/JDNiibc6YlfJV20xRaTQVgi+OcIZrzWdOxbKPAT1cX4Yc99Gzj4gJSOyVpsF9Cx8lNCqXQb6DBB
+cDNtRsw8axzhbw4GZDwRdWie9wi2uh3i55q/s+jhRFtHEDyyc6asNo3vySDfZfSgtLb6DRiVOuv
7RLQBqYxVKrZAPVkNbaO4GnXmF8e2C8vhzSPWur8sEhm28GoafMyNjP9GajxgpV9F/Gbp88QCD3W
WX4X1pEEDU6vA8RvTYqcRh4IAdhyCSGPLKKoH8MuWoAiEW9jGK1rDM73wT4KSSuU2s94KyEs/T6M
7P8G/zW6TgqYnDX+bks40/XcAr2poS5H1mRDIKc63beceKhL+bT/ils/74HAc4HD6w0mZ0jcbijR
5BJgz5SVJZgXjOIVT6fYWCoKkCXtPjXKHSUxLKQy0X+wv/Z2/O7zkAcvrgz6TcMXKsYrVP3nKw/7
9yDCc2knWws8srQEc0R8/oCqTF4KEvJjyG2KAJxqNi8/zSoZum8b/Pc4fX4J9yuPYmMvROnmnRcV
+Kb7QUG+yvGKyadTXtpSn2zLRML9PpUKni45/QRj/i/TEt5YYsgcCNyxHU3jcrkKkqCWw+Z/5YMb
J5CJ5k4eZSchF9hxJ4v/wwFwj+z+ej48/YwEwubIqG/yT/YdVXnch8owj27DPsAnWuuuOYom0DrN
sJiXewiVbqP1UUWwntz5BH81rvtw9Hp2c5GE82sRZzABZXI5d+rzmOZq9iXgRepPle8jEg2NO1NF
ZDiKd+/ZQ6yBTf24r5xqC9DC164FwgqGIhG8WqLmtMHX2gBcTMyL7Dprf0Lgq9IjVwty4oilZs8A
oBEL2NPA34+CRqvS6sZlWlFgx0v1PbawT2m+IpBihmWAMEyD55ufCMTEK9pcTZedZJeiBJbSrzB3
LZ7LljzCGP6UJT4DPeN4ChC5noy+9FUt2VapPde+Qshb3HHlT/JVZ2WQwfAhgXIgjEnMF7U7FfE5
5il2joRNcpvaPCjP751+SQVIrWPg9xUkvJs+9HdqXaJeeG56HVR/buzDFy/KHuGCtDXpkdf3t2t/
C/wDS4R4tSCORkxzAHUh4RTKRoIOtOUJcSotLjl9hSOvAr7ZYPRzfJL9spxw6e3Ch2s9qdNL/LN6
IbTwfalSQQPXGg7YvAcCV3XokEjiOgC5rRg97QNdjj3MiMxOlnC4QCy1bBVCYopmGZxvp3KNJEPf
zideqBOsh/GvQHuqGMNjCSdaG4omKXkBC8OqzI1dTyMeu4PIgGtA3hN2hs4YpREBHb3uhJ63pEn1
Li1ob/m65f4+LTw/sSBozGkf2JTTAK0yB86NSW6pl+75XZMqEfR5w3DSnf4mqHd3TyZiSMaXWk9v
5g+rAvRG2a5rSniXc1t1pwqbaeOsqev4YOXuoGPYOm8acQctv+LN+nQnypGy0u0x/BYuFRkD/n90
ed4S9VmNHdi/vAr4qyobn3cFyJG1s/Y8M5xEHWEdUVn5dOI+ppXNrVRoU6L6je7p+RR6+v768ofO
TPGeC7176Oetu0SFPa7w5bWUz3GRsnkcNI9G/OHPE9q5IWmzWPHHUR/5OJa58P8/3ScxGS93BiRi
qG0UVuEjs75bApxlCdc0oSUMXwXcoCyLLRKxO7QhbKrzJ+bU2fm8lV/p7n4S9rdL8TuW2m7Do551
WI2RVLo1c4hRX6rdmz0a4taH25LytVApxnQhNBpN0R9+iAlEIH+p6icbQBfRVc2l/l45WjCj0zJt
fWIG3YX3xSbZIRfYYTjA+o2hLPTF9aMnn1FgbMsguPpigI2tIXuh/C6MW4RUJSZdaDfG62fmyuCE
DcH+i0IeTxGI4QPK79a5Kyda7GeAeqenzirgBC3owDSjyknTriv/zejH5ZQ1p5nPA7pYWSI3m8XH
VzDz871ln4AbVYmbKhJKVnwUeuz8lLVdmICnFjJCikSV/9b/vs300cwqXHFaX7mjo0plYOLE/++k
NQOG3JIkkrGwht+bzEo/2i53h3g8rrgZiCD3sZejA2xraXkfvdaSzGdCbDgZOZVUw98IMBn+H2Yp
1QKBV2uoIYpGMPsCOsLDQyDDBLyRctjtqz612QK9nGdJotPc9DSQullaFo6MdzjCxJt+nufJ3t4O
uRcn10fCGZRwvc4DjbK4tmn21za+7IcKdHBJFyLKsfqnaX/XFd523a3JOArOcR/1MHlssuYEm/1s
Bo5GnhOGjWdab8HaZZuRK9fzFvKrH/WjoMOdf9BGBACSE46akA+TwCI691lp2EGUUdyPrrGn5Pdp
pIUVGdF70MH8y1tc5vYyUl0R+Kk4uc2/RulsW8OPQI16qdgrM4UcDjvtghZtZ5UkLYPL+BKNJ0Im
/2Zo7J/dltzaI35dPUdNJFs2IvVEX7xXi4CUDhru4DLrWLK1f9TqkKRQSbhNSYunHROXHe21lyfQ
qi+29FieuCS5f6Y7cqDp16O69iAPDV1oWK3D00/ayU9f7Qs0xS3Ji8E0oeG0t2TCzPvmXZRO+YMh
3kSayT6sj5mukRi3oDi1XldFGmOj92xpZskepEhShPVAigLWzVdbHXvHb7rjrRB8sRIk+lAe7yOt
vPoWlDMYx+T/C1x75KyQ0cYdi6GfbHbgBh3imIgnIJrBItpnCEVetD9TjrCqRYRpvHCvCoR69pwd
AJKnFD1dD9C4rUUAaWz0gUDcwfHZqi1J3cTCdorGJJUioPg40JJ7sGABEuoeccgKFvjqvCX4TmNc
M0RvG15sU6CIdnOJuxti0nf1wWWQus59NgLmjOwxMmtmY+k8C3PzYnsvcIRa2Fccf3BQ+/2ZcHon
EbfNb+Ql4lBESUbLLjzpzait+IeB/x0HHbmIc4Avgduo5kKZTqRxYNC1kHtVNPVgH7XFKaI3RPKY
yCKcz2bdE75w55g8tGGedSmpGW3w4lm2bbaCzZHGn8Zkcb1+0XmHHLeujlJ7ZyxPcGXp0CVJKRNu
yFniI7iksuruudjABUsH4PSmk0FCCdIWqP/kexeTn/ynlPxTCQnh0NBNrB1D1qtoWeo/ZmfRWF70
PMOsXTVRQ859lHZUnyFiPr98wA1cW567zXXMGSJBe+rWTqG9apG4HQkRdAMh2GeyCUKsHqsQrZRs
upnIaNx1WGJFYImUkrtJ/mx53GX9IWvIBUG6/pggz3P5Yyv/cLwdDlHzN9a+6DlIiXr6W8Rc72rf
w4w9j351qsdNYZHsdO57xx/bz42VrX+mbzg4U6hRbbr9NS8GUGGiRcZdtAUynwMxZ55jWoNc5SRf
x26eYbxHphA79KIbiXhtlRdmWvdqrt+VAKSEKrnYeVSlytQsYzOZlDaXp7ftx6SEwS/om/HFIrFF
iwyjCmHIaYevIyekRN4RCqQaxnTrvCrhuHASOegzHaUcvzsEM0SJrEt7vzA41q6CKP3q2k1DnVKJ
OWUiHej0ziFXwqAN8+sJZhdzUm0QrfE/rveDcWuJjwgQol5Aj+CXn4+LZU4ihtjE3P1XjLNzSr8B
q7VVbpwgKPAs6sOUOxdBpRe+jw3wtSrnT4T16dM5561K1jAvMX6IhcCIvX98X+uHksaZVM2uGwT2
RpiWSPentptA/LwJywB8cDYDkAevgAH4WOztYUCsPRxlainkwhZoG2VzybUliMlej00zipyQLb0Q
xZQmZGPtculYCi98wBMlC+x3mGCtdd4NTwqOIMdBZ2fNvuf6g0rg77GBxSc3np8VcWIQzsG77/2K
Qol9a2/yRH9YbJQ6JNHIAS8W/v747ozNRSNgCCldI7+rQ3ELi5mRO8DEUf8qc4pi49eLkBce8h7b
iWpb7ixKCS1kfLTN08NlYqWcX4P+PHHnTsKVJ9y02+GoOpebgWvAtaWlakVpEEHC3HVG653UIfLK
50eQen94R3hBqS36HcpJxA6+tj7lUXy+2QK2qBXeKsetN7gv0qn7HP0v8Zq6YBkt3BLrNaIHrFFy
4bLx7MZWFA+4IzYjKhB3WvSJQpTc0dTKqkRAcr/+LFu02ds0zBFCgkAMV7MeJqUyeJZiKmDWQ6Nj
63JAU9rUHkCijV6/1u7yO4zTU/rGMArOL5lq4qM0L6yFRWmNHX/BIk+B3NkIi2VNQ7fpTNoNAMGd
3tsxIyVDc0jPZMXL1d7HDL1Kek+a9W26KhSPgguC94BRBgseUyxQh0ADBp8k24E1sE/PSWHyt5yC
XP8XvZUS6pyJ+wS31ORt7nBj+9HF9lO48y/le6LilTXNhTYZTnSWDmfdWIddgzhMuMfFiFDSPT8U
dE3XYnNP6/vap2otzcWx9an8+vF+feYgGqoTgQQRtq0c130mna1dmfF6VGTdGDGF4OpeXrHIM+kM
omRr06jywWMLK4ec6qlqyBagoTm0PzoaeMaGJD/wj2/hq50yZwxYmKykHu5xtwzj+tBrWsMQ2sh2
wnRdTECTyJkOhUJXKQGBtZIaW+vixWULAX7VU4dB9Z7j/TW+Hzav8zXfMDWv0BFUk3bCA25VLPTM
gzFRZYL97BEKRkqDk5g/ZSxjU7T0dg4tBzJg5XLckJvmapuNTUVGKKa/WRUd8UTeoqLPnI1TmKcF
MDRdbtiSgZHFe7dGB+M+5AZrlz6fprYWNh/4CzU7rfF2zllC7oy56RBXesacHkeQoX4sA5ccIMiM
CprDekseeKtDAzL1vjfkkf/4sLu+NXJFg6LJxxTBCARCoTkUf/JxP/OjSrrOGb19vcz8g08RfYHG
iv69P86+eiJODhBQXBVAkGppTTdUyaXcXsQcBwfkY73YBcAILrv3irKCaCXFj6iuxwHe/qGGyKzI
XiluPYNFw8jsUYX6Qlk/JOx671rvZZGHQmBzeQmqMMykojTQjT9kj+7Z1bgebv6esNIM/zqKpOHu
mLHTa1ACXGFKuuz2a6Mi1+D0ps5PtqRKPiuL6u0GUIwWupcA/bAOMrYarHTHDjVXYfAXcjYAwHvm
Ud2Ew8CLbhyoJxAP+7ld4egKTftjJeqMV/8J3l3ztoBg6TkmIfKvCu2xxKZqU4oiwumNpGcMBdlt
jipKz9upYPVUwO4JlMNR4+wB92ZFbrexTtAG+oA3gB4skEF0Fpx7rWnSMve93OriN+Cz6LASMXFK
G2mSHonfOtfQ4srzbLoLvYuvttVZPK6HhJ3Tllex9qEcngOWAMryvEkdLP1NmM2JhJS572VC2SNN
vuIhwJSsyOYMRjYzty4uBDU/VhsoKBUtO42gYUKyehrClr9VcEzbs8hArjrb15gMEUCXm0xuOkKq
JOQij7NZBuYY5wZpx4kP/EDtzUmug/7ZvlXDyG5McYiAqaLetbl7aiq6FiNlbqkiVUrxZvJbc0hj
VRDltq48S98dB7/INKbMxEx13OTjqHL0sMtyYz0UDL9u35QH5qDfX/QSN0Ek/ZTGhSyRU5qIb8tH
+4u3lWN4kdeCQTsSwlCj0aC/4bNZenNP1vlTOct5rDO4LvvZJoKzeoLFmsCop1J5dJ/o986/E7vN
BHvg25+leG9SyksM78nQ5ew3n8iBOZ+hlbZUhJzGyHOfVj1txr88RT+UwWohIDfpz+gIVx9nkHwW
GvEGhZixYq2wQEBxZnz6F9lZtJhtm56vGQD3RucwGcnZgV8A3vIt6tP6jaVZ3am1GQOWq0OcP+aN
Xmowa0iMBykndiKMLH2d/sUbGpb8RDKWV1P1u9iHCicfu23O/6NSMzuTHFrdcCRGPg4d6jlw8raX
c0EFnLUMBie7VO+Xl5H3so3C5epDcH4gh/1xX2/jJYuJWIbk93doyFI5LKYk3c0bzfZwXbvzZDye
3T2d3x0OzWll3euK2E7wVyiuFx5WF8PAmoS6DaUZXYDjZjxJ7IfcJ5TQZ3oenTsuuCbeSab3VP03
1qohQNssSqK23Kn4S0VxRuvXyJOYxdeVMEvlBb8qUBOjS+0tj9GXs7zeoQzFyY5RJ/E9rTQqiTLe
DbHXZhVfOBxHWomJC09f0OdRId2YqaP6eLDBfzY82rBnCKZiUEytT29jTODluBgqVOP3ZduKMEpr
YbH6ocYtR+yX0ylzRrUvMGpYXQICsIm76reKGeunkmZbsbVmB039lRmApWuZ9IMYs9cjBNWPbhAP
bexiwjq9NkADCmn76PXCHWkWqQr8OHczHGgpOhpMJENGlVC7Q74oIDskp7gB71Jt6DL5IG8qbZmD
FbTfYtk3qQvdw+t0rWRz/8GQyrFBGGIgXwA8MP8oT/FVfOJSxXkdouxP82MBN8eqbX7JnXuGShYi
/Ml7aRvxN0Ce4H3zVxS3LeVKanjh4a6Rv9CFMRlztSQqczGnRGPgXhLKaXeWLD65XHcjSWuPxP+R
aZI1UBSYnwWJefkp5lcO43OsSRRmYgXh4CFOP+irk6gWlbJsNO1bBsjnDNYeyJcxGwR+m/bcIfRy
gGGvBASwXdz/42IiVGslIi1hmIxLK/Mv3Mu+yppkSbjfj7hx/CCI0WsowUYJf6BeoKa1jDt2b0sM
ogfOvNqWIsbfyi+5d2bmUqulAVqR+TK84TyawzDbS4XRs1FwbylvNypdQ3bE1A60urWLG8DlhuNM
6xAxtBRDVypQxECJUoTfETGl75OMWpNmT2qp8wG/IqXhX21CYhlhrfVMAbxjTLtQE/CovMz7FWPQ
EX5AQ0Iz5jE9LNtVQ2o0dLsXvLeG4SkDX6RNIzC1dSIc9T2/iepfn4DTYIvNCbSLghIAhrfLXU6S
Vp+5C4RoCL9q5Gt2CPdn4ARD/HMCCH2eS5NMDdz+jTsGk+XrVPROVu/fQfNIzwQrbJABiJBspTRK
sc54bND5I6MhyBr2xEL4Xz8WOnY7N5XSTiWsMPOxD8GLobu42Pckyy6PeqPDV/y0/iWE1Rb7T3CP
UPi3pcBptUJhcp3xEsTDdaOcUUG57EcUk+iiwwjR7ix5qCKbDJhUDum9bEIQtW1tKX3y2Wivexj5
349e7fTNBnzOcu+rCoSEQj0qbIDngPXpdptydep4BJDC6IKusklAqRQ+wtJOZ+iqlou8Vmg+Vp4u
Holo/T3xt1UwehFfYKQUYBEuA7AiGPJH5fI03uVGoc9d9MKyV74HNCfQ2lujkywXgH1qCc/xJ9Ea
w9hlslUGCWMl9qOJl2ZL32BVU8fvWFeoc7zzt9hn2C2bmVJLpnyvt3B3sl6LPSl0yQ7lRO1APVN7
if3htYDGaVQAmPuM8v2mC6qv7XVbn9Ju2UUQBxtLJOjBf/kqZ0PPLdwvZIXw4sqk0LXGHp/BrCMH
Z84d/jGrNe6HbqLMczRz28vnkyH4AiyeH+lo9Kx4zMv4HB+p0DZ7F4BFI6cB+WGeQ9gD+qOVcktN
uxiP5zAElwSmJRC/fHXApUm3vjcfEzfYBWZ1mb1dAzx5hJ8KL5ie915fejb5/53WEHBL9vsqG2qt
b8u09reiB8pPNdtRhmcz77cb7DT+4ILe7yc1UbEH1kd5gWatnins+Cer2BRAn+y/X3aBx3uTo5LO
vKtP6pfJ3pWfIsTptUr9lhL4zO6nZtwrSDDaz826Ue0DxZ1UzaLUvbJfPzDhfAlPEufxCpfhOjV2
798xU2E0JwJyaZR92TrEvM3P0B2DPO3rg6Z1nd7g6GM1HSosEl42YTtlcg9LgIvuFyKverc4is2N
+cUKuzm8R29dLcq6ZycayTOJObpBx/P491kK/GXzf6B6zr66mkQDWWcZPNNBFJTIxRBBqFBxCP30
Z3+QpePFuSB7jOBiMXEgcWS+6lMJOjFYKVrJQfCV1uV+Da8h4cv6ExpBBG8GvoaWfDCbOJJuSJck
iaJhqGAOYKvl2jimEewl4xAc/vaj5SS1nE3e7EA+X359kkjhmdcvzzB4oYuHQ6M6QK2qfJFPEJNo
glPF0DwlwI00/Im1GF95V1V9D272CCSGHH96301sV3DnqajZopgJrN/mOeikRP57t8R385O3sllt
X4dBKakxymbaxnQbn/tex5ggYSvtrske1wiYOFu+a6tC7/8JoC7wdXM789h7L8aOboCe3sh17mZk
LZ9tgBlQCV70KSQFqGw6mI/l2g88DWnYuoIGl9QOpHMWC6VkY1SjrRSV4c3z7rptlfOvjhmkPjcJ
jZKBCxeXdKBAkhq0R8u/uVHLXDDeo7oJ3DKTcyO96LIdfBevidLG819SlhDEESV0ZRj7yNleZ+u5
IUMNIPVGSMNyqaKlmH105kKFOUqA7bTfS+GalhOHJE9QFfLAvHRhnxegO82jF/8OfzkSwsHiQUSQ
M6jYyvT1UTk9/HPiHbPnE8HERS0WZgcnf8+Y35C4GPt3jH8AQlE4uZi/k4R75Q+kkr2HvwzbV7g4
O4LCUm7OzV6IegUsXZEwHRjkkyyLnwhrrEv6cjnGaXlksijYXcE64lW4xI5EhC0dxLhmHeMGmgo4
iF6O78DjgN7gQMqq0WwFMmVRaVHVezQTulmLzEZ4+M5yvMFrTr4mQNKAqIwW0M/k7LlUIsBbt1Dl
k3XsdpRrZGV2A73BW6kj5Ct4dfLpb5PTuPKP9Y6o0AYlCFBAiIL7cucE7BaC6AqZfymo7+SXXpbJ
39pE7sd86YBRHaff8u2pbdTyaUL7qHikCIHnIyjiYmqTOE2BSA5+YEvmU3Nq3DRiwoyczGrJDJ3b
Edq4Waj2YZO1ELab9UgZzjfxomOstLKE5XqldCEEzU3I69bwnUvkTLRnbKJMYMK//1wX+MFnxGAq
YVDdhIjGZMa/vpHweRHqNog7UJ19c0gOohcc9GPTatkZ0jMyY6BJZ+mVjK7H7MlpScXBKSYtRi9X
bMBA9RaovYFW6PBmOujeBTvaUILKst1M4DSoyh282ETVYbSCPkY9inubJ4TM5nLzhw+gdNukeVl3
xWN1OKoZP5uJU3elHloJLzmStpKyt7t0TdFg5ch/USsltrG/wCjryIgGC569zE0xbULo6ruHz58u
khDp+xzuDUWhW0srZXXNiEL6bbW5TBdpME7M+c3z4j8iX+6WmJ/TEQrY56DmkpIRhDDrekMJRvf7
DBcaV5xmesV3TMndIH8DjMXUwl0t9o5QrTG5N6GDWgE0O6VYD+0dtDeLDSQM54eWefUB2lu0hdCt
w08xnrDYSwqQMdHJtXZj0Eoj545CaFscXRglx/JAVwr8xav7LqfKnF9u7C26mY1WgCCORWho6T2r
ZfMW1f4M/5OsDX9sadHUlEpfQJbMS8O8zt5I1pVNRZvEuZeQBRQoYlSNnn+hNNq/GhvIkU6JmmpN
+xZQncuTaQIX6mVXqrgjYjpA7qho8rzbvQ1vMDUcP0Lj939e2Q000ASJAjZnOEuFYME6Plxn4M8x
6kyVkHxLnC/mHGYJv+MmWclfWW7BYlTXU785O7xzPDEh8Z5KfGLZtgBY1A9liS5S+dk/WGYM68nr
0dFCL3A/RrM7Wq7c6aQo3hjW4Ji7Ti0i4Tw58NjFtGkhAYbeXyKzLa0bCVswGbRKsL6XC3N/+ngD
Hlzpei76yHIU26/9SWtLwMLQhTiYNTSqxhptR8TcEbhoORI8EZRyC8hHQqFSDG/yPn+tE1SQ1BPl
id0XksxGjdX/l4SryKDY09UWN7nDQoPu5cA7gxIGYslrOQ8h12MgRaxDEKWZXiR8CoS/CKcG3onx
MTpQi3QBxGQg8g4/tUYtmF7F/sqpSevrTOYzOQFqXCgdBV+uFukWZaUYlJvXHVPtQopJSiAO0MtD
XBmbbTg4+WKOePHbk4YXpIjg1ZA5RTk8+2gMQx1uxTUbbrnnWc2F2nWYjdYatw0CTNNhDuaURJ3+
Q9+VfHzMoqkm7/FYMuEdGQDLTAfhzzncn+X3AxmlSeU7nayMBAEYfGc/PmT7r9W7pqFxiWS4mrk1
ADjdZgKlxfoVPKWIEuz0G6hzQvXPIsy+/i8r+/uwI8HJhRrePifOvgatND3TBWGNZan1mG7kspty
hI4zfNuj8yeFaRK2VV3EY2wJbw8nIrAp5gM0tXpvAAaCwaIwhorYtgVeAqK1qBVqczrs+przZ95B
LSQ3Jnvlhc/II1SO/CBSocH3qiFXgIcUHYYJecrfDAAeWEBL7dHSM+uTC7dHMGre2h9RXQr8SMzn
GzthwwlztLNvFI1KxL0Sj2CszvvMvWmxQzI7B2eN+Kkqfx4BNnaINAQ52Ki6RBTF0cxAmPY84Zzv
mgA1mukgd4ZgSek+m/odvI/KRxofKuMlygXitZQintKbcCmCkgyk0HmiqJIvDkmLIwgot8KMi6Wr
8DVwKh5PRVZ9M7W39NiyXp6Og0o0OgCpB5OaQ08cYJIrApzKECYJgs3qcJFfL6+v0itU/HIQ5wRy
qAbRJsG993OpLlfmnr2ESZdtFGQQh2d+TDWZpaz5mBngLqFJhLpnCqDNBIUp1W3NN1uqWcn9516y
aKqjz1e2wMvKprmhMiKRm/nrHRBFiHcbCcqNKEfSXhvYdHyIKYD3zDroh7qsFJ7ZRqNAmIt564dN
kX3KzINTZkT1fR8c24RSAUsPReah1tJJscBVbqTSfNqol2ym6y/7L2E5zVUY/wE3YXLKBif5rAwX
x1cXVl/Ro6QPDrTlPt4ACUHPgaVG2u3UAWo1/Iu1fbX2rCKnNKPZSXe5SeDoLwLI/CznMPwLO+pZ
aNGef54vkbS9L4LSDBEMs8VvVtpLABwt52cs/ZNHcMBWFQh+9cV2aM8JjZI5vwyPFfHRaBYahCX9
4MCp1F/IBisnvAad69Mr57nu83NI3fXNVuqmMPozWPCKSjrZiE3N4bMs/gC+DoGAQVn1fE7TOPYi
rLiW07ioQge5miSZQvKrRaP/GG9nkBzeniIiQIFw5INnZ9BWobndPdF2SvRMpnTVd76/eJYpMZ4Y
7bPy2pprXD7NkmoNNxolqsxgsgigAOBEVVX9WNCbBFq2bCFZTA3elFldIOmFXjKAwwcbRFMmPzXX
LlzQssSmlcGrRr2fUfxp3I+PqrpTx6lJxoypstbF/Ya5p3y1xlJd4PZFOOku8maVChP/IlWZRPH5
lw5S+YP9T7tymwhWEu7X1xD/6REFsy5uY0+tkWh4gs22APfFf2c9lOA8RGyuPctE0qDMIaWQUO8k
tfLvyer/V0CVwbpKoKdfpwCN/BdHIDF0VlRMgZtDHKThR7Vlg4UmRPwY03Pb0ZYHBTU9iIdX0yVb
PCVJYiXjes97m3TK30TyJApPDpM5ftNaxBGbVusxrZ184I8tDIdZcl0aQpxkHwxyz0E3HFyqWbn5
igK+TVKPGNTCD66n+udtQm8gCvdLMpiK/exQ5s31nRuFuLB/SZBnT++95etRus2RTnsta2sfSoCf
IubWsdbcU5wpU0KfjmvigvSmbP1ll99pldzen1PvnarY8atLXlnQODmEumkJIzUq58f9cf92hB48
ndUJIBzZC2AlFNrrHYnTlxirywwjqu6okZ+mEf+Ve4UnfkZGd4iv01h7YtxqmfaSQpYCqQzifiHH
ogNs6rdTUyspTq2RA2p1l/376xtcNAq/ij1QBervz/bUF7NbfzI1hNxQesBWhT+qD3NpBkMXfUS7
xeJ0ZwEIkU/e1EqJN7H9SvOYP5zWUL39CB2dxeW1QNLYuQWz1v8z4DrKmryPnmWVAcizwipIntlf
ZwvYTjTXN7O4afvZJRQV24w8VieReQfXwxBfO7ZJ8p4rmoRqVwur9lyiLcjvD7hTbAsfzePSJ7dk
p3YQvUXa+UdXIY5SPyWvumdjEMGdz6df+kKgr3MhU6owUXbS/iRh96dt2iUtXIaM0exRfN7v00uk
AyF1OYJ2creI3xbSunk3ZMN5jninrb2mFg0jcD0/zJfiONU3ZLIM1DhlV+UjPXhOGzQB0Q871hbQ
mrt9tBYcku5AGBU2oftMZte/QuGu7pRQNWQ+CHBhQ/LgCiaOJrI5hsrzias9AXp5Hm0od9DXHIb7
5+R1rYx1w3jWx+eQTvJyug4s4hVhjKidKGOrspPpqo7SGuWoBzekqzhPr5Ju3wjl/HLzECspOfVW
vIFz2rTAz3llTYbHjjlY5QZcHfThcl3fWs0tPm2In8XJx26iMoBtUrOBeZ6wZhGeJYE8kKGgFChy
4ecfK8dkcrEq6OywasPgKOArHNH2VhLUcc/0s/FQnzpH6CgWhbGBGZ1T+0scr3wsHnxK4epooYFn
ggNz7UPEHMXcHKdNzGTa/wTHR6WUulBXWUy7mWcTfuPPe8i+OhndmceMmJjMq3pObh0EryKGKmOO
fZvXPfsewLmqMvl1eWjxrfgb5MBjEHnrM/nPvIY4GD3VQoS0w7EvGjj+2GF9jNz+U21srspBgzPZ
mZpXbzXX+SgN6hG7QGUvTz7rlSHc/BAwVW22I6FaKy+8j/Ceob+n5kXd+NRZFEK0U9SoELidKTD5
4htWm3Gg1xGtx+IAQkoGlnc6iDdjzyXxZOBGNOGkDuEYmj49pKUCICJpM/apQK7jfO5msprAQWHi
DyLxFdVHtgscRlLwU7WGbM0YyUer2GHj7vQCWL7MeOUPELx0UPwQhGx5aycRItvNQIGj27DBmkhs
ZiH+IJI4L0gRDRQFVPLSL8FqPUs99zPPTuR2pB/QdpOCB09bBA5Cnp+9FmOmlERbaUY9b40TldSW
Pc51AozdiIEr1c15uwlg6SFcVTJ9jXVJa9wHGJz07oUrRAMauDb1b9C8IzMAVBqM7ddzilnh41/X
fIvEaBSerfKzwnPidMfleHnHp2uxR7Y4sOglCkwMxRQD+Wld/eraRAVjejRDNzFp1hcaBoA+uwF8
QSST2bTj1SPja7D0cVZKvvmw23gKxKseM+whbKmIumJlfMXboNQLJpgVpqqjOKySO3vc+NBb+JBX
mwuaTzy+sd27OV0atyVja6fRxE7R/1/5wTdTw3hqpp3yNkawDsZoNq36fV8Bee4nQTJeZTXPbEc5
1iqPoGMj6IPOOaUArYv5JRPj01vYjY2xAsXWzxZ+UDJtytS5SsteEwKcRRWlJAUgjgq3eytVmuzR
lHXu6WpSQ1Ic5BOp0WwSAhRdh/2yn1zxgyE9ieZIFL+5I45Bf0SGQXKWAbbnrXJp8mtnz7yzXU3k
WJF0VTlfCq2iukwAuR2yTg+kl85pnzzb5zfOqJU+w/oN/YQBDZPdr4oMqPhoyBrGMiwkRSTVy6We
AeshoLUMNjUsKoQhKJKZNt+V2nt2HaCozCIrSDYTw1ZkqqJdctmLS8nJbj6KjZCPkcOQoFVpmLEW
JrqhJgJcItA7wIwmRqmpB1M8tQbZQY1g7faf8wUPDky66q85tjQxxgOMguheaP9P93dhc1AGp8KK
0z3zes0rXbB0l4qEG949Oj6vtUhRp5XGBKx4PpdPTWqbmuXKirbNvl5dpR3OIaSU/ZCGAqNzPr49
aqCbu6Eak3Vyn+5mGB4zGXqCNPB44lNNZnBs4IDTgaOTBXEDeFxxwyjF/QQtcil7YvehRaeyMsva
x8xpSCVIURaae5yDT2OkfHRegZhcTQbLog2o31mFZCqyuPoljZMZM7SFeBXqtmxZvPyVnoLYZvBj
1f8LZkcC7fyx9ut0uHREuRAoJqqTmfEGklGORzStqkjg+PFz8O7vFUxeaXbHt8mILrZaQWWUmIEq
2eKY1cXee9YF3P6rpCrQrTEwAHAOye9aN+WsiiSsf/sRnGWuxVq7NlKRCh60IbUKHG1YE8P/bLbk
VSm7xXnkj9SvRhPWzy+w1WiLoWuqwqhcB3262DTMh3uVWorpK6L4EXQ10yXXDTmRB+8dLvb/PL08
SgV+gI0Z6PET5SBm3QybZqFRmrUA8Qr9wUMm1GhtWJ77LxNEPUImVGRdiDhi6pDpq9rgWk9/sO5b
6q80MAQf5GoibvPpDKVjt5SiEy0FRR3puBXibrrXMT1jjsTJwFL+R5omO/HJJPX7UBKJ7K4LBFlI
8csdWsu/1LLiW2znh+cDnAy/dU8MqHIBYtBXfN0Af7kBB/K/wknEzGCx6YpWpSM5yELH7yzzPkxo
20hw0c5Njhbd/VzOCfQGxoVuyDpvWPiHA4GlBVsH6CP0Wq9XUKnYguYKle5gqYeZUQv5VKdTcIJm
8ZPAzZdVi9eB9HyPN2ajSXcAjWWt6c8cIR+/iDnSnbLCIsco6k7j0RNazQgo5Fy3YvRjBXxR841M
RGHVGDEdheHmDILrX26d92faQRnCFIdWvSBFhyvRsJ0AV0Lss9LDWxwjXFYjiP+HR8W2+36tLXdx
r+qdz6a3ngF+NmrUAymUcsuIYtRjFSesjyDHx/EXgcDd/VbBuGBOQoNXWZ+GZf5MyZY97EXHUYng
59l8pdTXzStOgmUkGi0yA+ZFdAV45JHUPHpUogv/G8bmWzVLy5yOGcPYLDAV0DD62PWb+ocQLgwq
zFxjGU9L7AbO58D9CXH4ch/7OEM4kkMM7+u0d2W6QeHssj8cjodxNM5GxFY8EPKIXAM3fSkvoszn
LbVLbNLhw9vrkabSoa4eyRjTCWDeVC1XuwRPDqb+Csgdb3bSyK0x+2lhPnQizEdOy0TaNgQOLn/a
ZpQNy/mkivx69jhQ0+VNyUwLcw3gxrBSYwev/LeGuKBH6YP8zu/kIUgJnFWM6F69CgyGoFc7FI5q
jJ/5+B2Twh7A287JPLQAg7b1zVYPIS+A2wISVkvKA6+dzTqZ2CGVJnfFwaMzoyZXUWTTu1JzxH8O
5JDYpA/ClKaIAgb12/IsCGc7zoo8074rUt+lmmBDSapja8WmDuYXCMYMgDLXuOs5YlkRKSy+bjpq
qH3wM+HdI2jwb7QJZpOMreC+3Fn9YuZLPtZHuRtoq38FTFQ0320oIfqv86P1puriwvvQoZeZHO+u
+EOW33YrL2+G7sWqQt7/eKQBL6Lkkmh94zrxeazWWHQn2idr8SnJuu/w+mVywA0RyKItjQXf2AiV
qG01nXhlU9i2+Y07CfdSVnVWGQ5OS/I8xs+T4vy0Vp+TjLS46KVFJeiXuEVflI2alyamaLE27L/e
AuoRvW0Nyq8TFR6GxkhrmVKkX1MFgXvg5guymh7OR8YdTq2Z6XrbDIGefPB2qN/TyxZ5UPQ3Ul8i
WQhwdmoo/+3RudXMFOdVIas4NqzQcBoms/yGU6t+64aIyRHSKpjDm0xJqx7HP/HMJXXZp17/xev4
K1P1zRKOJ0gKUhV3Fj1A7sy4aWsXSOeyc2YD82H7vEXFk5oRfLrYkR1BE9cbY0Z+6h/eXo3Awg0c
CiPfRdV3+6tI6E6+AT0XQLwJUm6kVVs+0A7FQf3GRhtHLuCYDXbvN+mwpm/vWGAUgbA9GzE+4Q4q
QouQyGVALNJKdxe4Hf1bPJYLRErpHF23/OpfyiedkjEAkcUmbEJiQd2VCT92ObydPqTF/1Bhe8PE
1+kLFLglfi4d/07B4A5vd+oq9K7On0zJk2iBcmcONz4j5H4aylQ/yv8BQcl83N7FQMbgDCNkdh5O
g+wUPp3cGAV1L/+4CNZVv0FGdhkamnyczIZ3p0VWPdUqhLYNGV/Bi3L2CVl8lU7H5KRUyJQK91FI
cQxnH2tpdB5AJ4xpRkJ+m7HNp8Iq8mr5b1xxDurjYkWH+vhN0pgFlbA3bDc/kZX2hdTaXTIKIyZt
+I6zVhr3ikkg9rXRXGMsf9Nug6moySIP0FuZlkY9XFRN53StW3LXkCJKcp4b8OEzH7QU3p9kVokE
FZhjb2vSCdlbzn7QoZLyxVDaS5lQzgyVvFdO5egsrZR+TVVLs7ogf6NIMqIn9NALVB9fD0O01Ey/
YKTAsx2gbjQGGof8ey2DTKceydNkEuAlwNxH0H7Rcsfr1mCjk2N3Df4mUx+fbcxJSFbjY5dMjgqK
xa5H+nwbqYEzwdE7zWm3HW7LdfZkLRQcvqmm0HRnMEdgf31xlzG/MHrUmx6Wpcw11RYbz2i4rnJc
zsytKYFNOgDtCI0GZ/tZ4fnhw3TDuaj6Taefc4bJj+AK836xNZ+Mzxrywe7/I4DB6T2Zu/5BRhtT
b4RANcofLGW4i6Q96MjQDl3vfzEXRoRBGBdLrQidPMyaVtYR7geJsKVuIB628vzjECVCTZNSe08q
v+/oRJyx6F+FqRG6ROjn1fxpfeMgh9nSOkJPMRbEKEwrjQbkBBCJLX7P18wCbJHWB77LDDRM4pkc
Rkp0MBqz5Xk3uh6zqL5Pt+q96eALUTkqD2AhCrGLkzdDJ8rphoSk0FtJhhRUOmI4g0vZ5NAASSrY
bg4H8abzVqX2wLUw5yGGe2Fz2LSTU9nhkIrzMdOPUqBC+ZJl48kl5+a12AZhR6o1qkM4gpmLCY7q
8r9suIZ0mmE5nYQiNOlGqi8v0c0dZgz3RNkGEfH3QLQt6FzX2AEfL5KBZmG85pxe9YqyJ5THeRbA
NjkxGQBL7mBQPOZSXkWXWqT5N6mI92CtIlJv6BHLY9YamaFv6hdF9SdpabwlwG1kElRyt6osRXrw
OhFedK5kdBM4z0/u0dRilJyt/I0E5RMANtuaWNKzh+uHXXN42AccS92oJOvaZiqNJn4DTVvnYpLO
C1fOMWMWfmQjBOUrmJArnZBgSc2w0K//Dwc533hlfHA/sUs7yrrz7pahOrhsQD28IBWbxwUT11ER
SHSlmaCLxnG0UlyRh3KZJWMMx/kjKUG4aeDU74ZIGviablhmOYtZuZphFd6N+O6jmABtSK1XVgLc
IUyWfBxiRp6qRFpNZKg29953z1uqmyRZkZEPzl4751jqrTsDbYMZJhqXVA+/dMqIvf1Q5FENLSBS
/PmUEvWjHGUX2kOuo7BeSt85oc08Cc0bAl5fT769WuRd2lDUIvLt8Zl0vTMjEtlGc8Hrg1r7CTBT
3UM/CW7S2tYTPqn2hk7H8cLNfJbVwT+UfRDvvwrnLEIGwJwj6+nOm160omgMmbVTSZmAkjPgmPCW
atlgZ8CYNvIph+u30oqx4dqr5cw9oZrJtRBIJ/V38ZqQqF/TjhmHMJfVPW7Yg9mAzaSWUctdrdVx
dtwrqW5BqqPfqTMd7+w2x+G/LBoIAHOnkDM0MM3Hhwv5kfFxL49S2Aqsi90aISKyAFwQxmNJ5JYY
vYqpYKK1OUAwBxMlkgJC98W17igI8PeguDO/AhOMu3OT/aK0MqhS4gPJQsnaLzkxjDaetUpWIPl1
xSWgU8h3uGl/TpkoQr9Q6lrfPCTxKfXDL/L2iuNPpNEZzBZFH4pv3xP+I/tUnJz9yG/di6Ow6ewz
lBusTTDQ4hNrKN+LjfKsFJrxqnlipESQOIkAwRLaacSBQJ3TO4YqO4+KKaqK1TeXx8nr1Ra0XB3/
bCrKvEWsWAkFQf+Uwt9SbzY/t5wCqJGb+leVSuoEMFMBqR6SQlSyx8Y1rMh60V19yhf4SezsT8KG
Es7bNgPYEmtDbhMm3fkeGX53QVkAi29SD3QedgNdMdpkt3fd5FOxNI5RStNwrRz4TguhwJRVPtoy
FLnozV4U5j/puCovrTmY7zF2kflfW/+0iuLT35baGKL5P7mSfSxUSITqNWNMauPFqJ3dTiGjNSSk
6mx5AyBqw1Z+QH1lkl0l8q5y1DbheCxXXWWQppoD90iVrEsPdjOg9hCo49ut+EtpJIo7X6qw9HNJ
I+J165PaH4AZGbH7CEhiDBn1Fz1+sszFI2kl5tpeag42w8+NrMuYnifC6tTdeQIk03hNUsTwbTiz
clX5IfJ4zZ+gADAplydEqAKHvE6EUW7YcHryW0QPxfFPwhhNOjCBimEqFoH39ozcocVAtNQMbJnk
lHZg4yHXU08xh0YfYUjz4tlyojXMKN4Wd1TSzbdIGo2ZgWjqHQFbQ3X+MAbGicwfT4s9wq04M9f8
zdjwZJy0kCDAKrVuSf0kmljPW72Besqs2v7Z2gRBT5POhSAKR/tf4rI9DyGFqg2ZV+EZf33R1w9A
z24iWYjkF16OQXxqQW0qySleg+th9nHJhN0dR9NerBoosSxhh2UZxRoux7Aqgz9tobOjcLAgf5Q5
iX7ZuEiqJLL8wvVyHW8TI4QGjBjQuQo+VEDRl7ofKYWETjU04pDgWjGeKzojzyZKkBM+f4poiunQ
D/1e3z1TwnZLmgg4MXlDSkD96o14p0L+ZzzFGJARW+yVmTXKBe7AB2EQSnhwRJXD1wrLTXrE2ib7
uQR0d8pWaDTF3u6OIJqDmJlEaqEvkajqnjIMhhbjLT+bAZGmeHQHJh9Gr6HBn3M0b8kQNRLKm/dq
TS21Myfyogp1h+dtrsAmXlkbRI1vDt5ojvucMr/rDmrgonGf+BkAJnxrLhJY1rDIyrzOPq1La9Vy
rt/nBn+m1Ooh3qyJC3NNiNs2mMpbHnrkcYaLl3pGN1w8SZ9cZet6QJabqbcdVjqZifSRfFsdRa0B
97s+Ljz8tlBCehWthXNFu1+IPmCB0jz1Yxun9N1YSfDVRSbnSguf7bhwfFK+G668shHxqpOVOar+
9qHxc7Z171bGPbzNe6vShsFrZiM9WcGSbN/HnH3msYimRCJOx83PLVpMbUuuUbu1czQlXjvCR8Xo
JVkiSb6BegP5GzDVAyL9XZykEY31PuC/ZrKB57adewBaYP9ux3ODJt8CTPgov30KJ9q6687QBz6e
QKWKhVrjS3flWh6FyTAI4hthg3PT9ON58CcU77y8TYip/NteQvdMgsLHfqxYUhGazBtF9zSlolsg
6prDhEIJZNnDht30hRwNzvqF9nlGShSQm6aXVpyoROgAVwZRCwkmc+mRuqHI0/3+LcPa5hExH7he
dTpOoue4wb0S5XUrJPn1HzUPUsO/kxKXX+vhKlj0vW/h114UwDDDifpzYFtDmB8zjkHT25Z59m0b
NYt2t9xxdNWXjUkL+gzD4UZYMAyEKUwdYFPsgHi6ETOTosVHaXgzU9cWXxVi4d6zXuiUoaWh7gtb
IMa4SkjWy6Kgk/jOF/zV/GIt37xTKrfgOzIPufzcLlJ+bHVBnzjDcK+LNkO8Pe9FeJyvE9hsX7as
doO7g9DRTn4NSPEJtUpuAKBMqO43xoHFHljmyHNbR7p77X+bsROHj0WCb2B6oFqlUe/i2QwP5V1Z
jKBZvR0CtG8NwaQlnaZihHHiLNhKq97yVU4koFgRofDhX1l/OmWE81oQPV6/CLwGpgSNZknYtwr3
QtbQHcWFwAz+jiiRijO8S2n8uH9FlIz1EVyXStZJGlxG/ziNbV7rAmD8X6FWnPyQVf7OwG+J4s6s
4pf6j2XW7aX4MuGXV6Rdds+jsJutY/YjznB1QO4I6/HW1faWR3NMMNqUhaNPjmGAphLTYdoxTPSk
0/hbCr128HkCW9NtNsgtrOyIeFqOTgCphnfR1V0TrJk3QnWQACQPe4PmixzpSMMfow4hvVSuXmDW
K9Tv7yMg+mTvvX9HnMlYw3jj9Gsp7Qjbe57e6NrR0BKZoojLBQGKuPR6GqWiqqDiHIIJivFqqYLG
Rk7Yz3gTodm1o79HbvkwhOYL5TONT6Q+lPo/2+IeIljqFmd6w7ew4cxh2dTsB+vg5kJUvWpOu9Gn
zf8OGgJGv8gddKvgJzRAmEM4bKSDh0J34vIfAVFilNpZGjmGJ5ezOS9roWj334KV/OPJo6FTfBKO
Mr1x76h46ROFYgpFccK9B37IXKQU5pE3cBxM5jC2rDNQjOJ/DsTV8ytdN6QD7YjMcq/HAFN1z98g
E+o0+yPZCHUMsLoTBiPyH1b5Sq7Shd18OpqKLobO5uhnqDkIjZt2W6J+w1JuZGrFP/81snEkDRpo
o4LNN7ejnKDla2rFCtKhdvAGfO4w0WI2BfsiaPGqyEC+t9klD1hXzIS9VBOViYLuayztbttxTfT/
gysS2fdV897Vece/7+SfAWF7Rm9EwV2Ov1IygkOGgyva3AurKKzCB7HxCw1HW4ytuaCBAcgEukOj
L13ql8KtxkBrjnmFIB2f8I6JG4Fx89fK4Ql37GukLT9hTP+fEZSLgOLhKjV+otw7GW1wZOnaTXfI
BfTF6hhJWmzfZS/XZjmz410nioAVOneyJb0Lv9RnvQ2T/Fuy01pziJDHviB6JsjrL6VeEvaUkBHF
5NWZe7o+0N4G5IC3McCHYDhIC4v1Ug8ZB64R+0auXtxSUwuhY18jJCMYjqUe0o5PhF64WPpc8Er+
ndBzBQeKZ3lyYklGT7rINpcy2RZnMYULjcdDdnBPPXz2fSOVjoJXMUzZTNutZT77DJW71P/EPptF
WR+KBoRiQWeAB1Sgmnmx0w6t8fMLGDssmPZp2tRap0K7oAqFrY+005U4hw3FCsDzmwLc7ZCMAvu+
eoBPcrqwqrtupwaozd93n+YE003EGs5DTIMj4uYRwRZGAzbz1O0stvimk+qcmmtotpFVC+1fY0xk
PGBl/x+Mvd6mJi3vZ/GE3SH55v0bynBIS6tfSPstr33lSp49keBlJOqjf9TY8SAHzvpAnvYFuN3W
shB/K57G6anp5MeIpe4WxPMoXJf2HgJwpAZbh4CaJG2ZkXQ315J5UK7KoXvJqI/8PVakZmCD+c47
hrds3WTF+RG5QxymrWFulAm2EIZm07UlbeFrKfmuATTW3NbYNjfQlYs2HM+8F4ILDy7mwlg9o3B5
SViSEeDgha4pMmF9Eo7noH2r7Y9T40fMfQq0XB6Xf72YpMwi9xiU7AaCbTYccyhcmsIK6RaVYZ2h
IxoIEkm0dAUOTBjtcNl90rFYF9FV1PlM+2L11JwAsAXvZXPAbX8uJglQfNT42aUWHnLQmDa7y3FJ
s9DohR9ziYlIE6yDQbc5mRmTYhgs5M/prI3LkusI27BhMccf0W0irLz+qBALNL6fmkOu+Z4Zj/+g
9TVduDej5YJs8VkFkSUAKmOIIN0uFQoSqShlE5/sS0jXxXLdGGWaUX+rH/vSltdT99zigZ5IJWT4
gi8D/7f3cXZf4E0NASzMA7QQV0Xlxnq7yYKgiwnC1DE+bsaIA9OqhNmWe//FIT9mov/QS2U+onU2
HjHMIbjgzQwzIXTffzsKhPadhptwUBpM71wFbSaprEOegWvcg4xLfsEYVSpxatyTi49F9FPiI30W
PhMjd/3mTG9ep19GHvRbx3nMOVcEqIeOm+UVjUf503BooPA5cLzHZY2+VHRwMpoR76oOXYhmxnKc
mk0eoS0RySWuNiIyMH+GotGoajAj1sRbpYZf4+prQ2jJdLl2uWEI4dLjSqKqcKEkAGOMJmyBVAT2
dgRydNkWYpCyVqWnd8PNFswSzDKhcyDis2wQWD3XZiewWy8No86Nlj/FVYPFrnOH4Q0etiCygAs/
M/J2pZFUyNrRqROMsYQPOQBXQ7+rSkjnAg6p9yoVxj/GlIANPaulDhQ+PnMN4xP+0QljSk6AQ4uU
TOW9FiSbthjkXaozRKKkh60uUrR1cXpeE8+TerEYiAee9MQrf8BKZOAUuQExw7nWiVv/PHqHl0O2
wAqXUndQQslQVXQo4/CPluar5hGfG0MdnKF8BbHju/UHR0Gs/i03G8hn0fP+wzRniix4oZfJ9EH3
YzUst1VZg6jP5ElYovSxWpN6YXSh/7nOS+FkhYgQ/kglmUPaAD831rLYLevy1t/09rKulvOLkiJ/
ir9VQ2dFRd5KrzgQj+YREJaV3T3NPk8rdZQQGeM4Kc+sP0idvizKGLeexiAI2Nz7lsBuP+68cW6x
FGFolCBG57PKgm67NnVwGv7NctgoCJsQuWc49Fq3S2UNLRldDA14n+yaP1od42ieXyz8xPrc3TrO
78sLTCNwDtnr0xvgC9+LZ4S/QVQqEQsHjC9RXczBf7W5KHoXttbveEy0dVm23HII0IlEtk7O0h4x
d9UQ4Z8ATmAzAtX3kuXWENqusO6QctyHMwTMfIYWdZEiE8LOZMC2xX/OzCmuXeuE6r8gFm3M/I7l
EFZ5f7/3tk/+GCQ2lZVGhJ/JJ7bSXAbWvg3onPPRGx2vVwb5bJbk2MK0C8CEGj3naQKCON+699YM
4mNMoUTFdL+8w/5T372pVdZF0U4YxSddVZFspAqSo7a/2u8rqOoWN8Eb9vmy+yDZ11F+kb0nb6C4
CoFLjbQczrjA9lOgBgFGhyRvdvNzyRpD1zLC6drU5gjVOmSmEuen44PJZiXYztA7vvcvKg+y0Ej3
sElyXCxU0B1nnGKRT/t59YfGDYMQJUrubMobnlysZ4/qx5Gys7S0hqWWLRNYyVI7kjxWJNLk2Lfb
d5T7/XI40RAdPxjX/72z1VyWUXQkHl3puE2Mu3HCRt+etsRglFOrcPWs5lynVnW/kRFjNixhygAU
BlUFW70dAxobshUf67uEordrzcvjlERsyt6YqTXAW4KSFY/HtRgK4pg73Lbb2QRh2iYOiOzz7ukO
tSDDBqwxEwr46K0Ed4rjMPb/RURGoHISd+X9gOy5Sr4VuSl946rZX3MRRmysKLHT/9rn0NhvzSoa
weakAseK/E2vqlc1sG/rwQGaKXCVg5vooPv4DbpbAGV9rfNIfrtf1TUPcqlK8EsgFEFe6CkO31iA
TDWUaAwUeKIBVPalQJS6QlCNZm+GsQ8a2nE0E1rXEttKp3tkTRxhsyUnVrntNZlW54MgJzgiwmuq
pX/E3igLFwaWAscyp+v7XIrQivLZLOz/lxTRsUxYcKyKGds6UR9GjHUlPSACW0KrRHwqu/rguqZg
p9a07Tbfh6Ph/GEcxFRS8MJDiifOn4x2NOY9s0sKNBIV40/RVIYOk354Ob+BfhCN+yabHTdJuhny
WnczwuGDwxMKssCCTLoGjeDZ3K+gCzY2zwkAlVL6Czp09xqQG5K4A+c7ij8+Y+5Nu371knB7DTSL
s7LWzUhkvwLyPqeR5AIUXGJ9QIoRu8w6srWDCDQAi1kmxSuRlvQKYZUexO9LTVy43owWGNC33pPJ
TpfarHPir4CP2zmWvLR2Wj0hlJpRVgdgAzMUXG3VT7a7vnEp3QMr+LiNNdB5jYmae87KG+QqZHUw
a3ut9MvliE27zryUUkBKyHT+QdEO+hgZEIdTHfNWXVSMgNlvJdSg6e/pmeHZdrP/zFwF2P6emSHn
tc9BxpxaThgMz+6eOktxmRS8Pm5fFdz5gj8I3AW6z0UezuKrbqrf9ZtbvKFc75bHSr0eScw+0Acr
DFf4uZqWnnseTzYTU8RWl+sSnPG6uIGVWqkAXzhmxYmXCv/XnwnxBSeyuFqiToCVOqDR3/oytmsx
pAFfVYQE/uQt5xKpOxeY6iPdmfL0y9/f5bO7tMV6K4L+MAIUkzc1rh4pMBFK/mgxaH49emXAVPm6
LUPIMIl//mmElRzSnBbl3Lk5a22DwsE5On4J1LIZtptHMfx3vOFlJzuDerlgjvTrpFVFQvx12Ra1
HSjlYoOWkrelqAIPsY1j80LYQtDQKXJ9jMlqoPRaGuJ8Rwvqy4rnNpYj8aKYX4uDYMCrzVp66ol7
VfqATBMc6jJ0YSitQu7mNCSGHkRtRAITGx4QkRjaRczmY0oqfdw/YDsjcJbJDgSBf8uklyDgcRFl
uJYoxh7kx3TxzNxobXer1DI9VFvktlDra1qaahKV/iJHsCHCBmdjIYpdYJQMtdaurxBnv8QdzNlX
pZllFKf1FX3Bj8ctNzhuGwNOR3gQPdhG8hYA53q9o/6wTs8mDZT2EmIytwi52iKsAclv95bbbaws
PSWH6S2gA5TwryTJpoZCnGy7pQOdkOMOy7p152Yu7F01DO+ESF7ZVqSkcnrvEcm6+mZRxDSAS2qD
NJ34h32j/7n4h+11TSSzyZIT2f5UZ72SlVZmwWgAutUpIYc4wo9H0I7MsEbISWVXGgqqCnQa2DN/
peSALgVeNrp4Vg5+imUa3zJzXPThVO55oCpQSQ5wvMz4eWC0Kz+YxFq71qNAGzZ4c3c3Dvvn0HdO
wx3sQdUuM3lU1JrnJUjJ4y2kq1c0+vZsbX3hbD+As/eAH4UHqIvKPv+4J9CcWkKqCFT21Xl43Hg6
JiOpuo5YKJsveoSCF68lkueS9GQd0gNJrlQ6esq874Bdtq02l8HebMZlrzB9Uk5zKBtofmnEt6qr
6R4ACBAPdQA5vQFjKK0Puut8W+JBbm5fVD2gfCiKbxAxDvRJInbN9usKKMRnxkgOSI+VXcedzIAg
bDQZ4NTKNuAF258o90O1T2LGYb5+6c2H945kLBWYomSCGkRLEOLx+sflqJS1EzF9hRCa9g3xZyep
l1ak7J45T1herCYMK2Iyk4JCnLKRv6XX0y42E1eI2xA7E+4sZZ79f6jVLf/qQrr2kA6Fy1S38OvZ
uVWa6atIer+/NEFN/Ou+YqfHhTZFMVK/XLmDGhpCl3DR9+am1nnqOxhYNy5x1gNT2kPkmxLC1ucr
9kVxCEKV9G1OuhoqvrdnUh9naNhn/MMJ6kuNmcFxsioGL8GvXupUtJi7eOElH0yqa+TYA76bKM80
luJiWixEnCoAkL66M6O4qmI1k9dH8i+9rGWoGIPEoUvqXO/zPUDsJdPPOydYkNXjZn5AvTt9+RP3
r4F/rxezzDuKT3ytV51tY1zG+Roo/hrbo96R2vB3U47vvfzLyEnNEhkNSv2g6sZwwA/yyLUznMoy
Xx7rrI41uJr1dsW3PsGzGeI9w+3a9G9x9RQO/yYdDxJvuazn5UEST7V4X0myC/LNrh5AHvoy4/9g
NKjAgfKN/I9e0P3y9ZeC6tTwKBm9Exl5oht1INx9d6UPzPRcwxkdUH3WAkxxaCfZuvyymYd//Ejm
9y7g26PX04+rnIp7BCQpvA8aiNgZ4xPW4oq8YXNIM5tf4MrOE81RTm0Jd6++65ojvTHpjjvqA1vc
SLYoRBnXK25dZxq1Qo/60H6dUzcbfOlP5y4krXDVmTu8puFAuFPedsDz3Eg0NQuFUZ9nQ3R3F/qW
VF9BNc79xTX8kJGyUFW4/zv0cYL20xpJanDBJHyPDwK1qPYIV8/uuj2Jsz7maihPS2K5S7+L7M75
7CjJe3VmAJ7acoVMO3IYHWKDb5DLRWveD29FMxIOFu53JuJLctbH3RX83K8Q6soNpTYLXWU11VO8
rODSVaAlLcsAIH4xNBHot77Ppn8W6IYo9JLzZ38XmWazsePIlGYwAhgWTHB+a1XOyLcxCkLkf+eD
J/DsWi81pURx7o7b252UtE6t0VQEigHRMYad+4+tfvwpgcMfTv02HXdF7Su1sxmIymGaDT1isIiU
tV5hFK84jeFqymqoz5R/ak2olx8V4MNbOXhzDk2ZXMqXkC/eD5Bq4T3c4Ba6RjZqxOw/5dnX2gPt
elD13Hb0hBIasnSm5ozZhZGkpGedUSQR0HA4YKO306xGGJ0NIt79yx7eGq7rtQMT5XqCYcM2BZ8v
uuEdKmOF+l3NcjIjTDTjZB2J+EaPAJaxR7bzbV9ISC/in+c7YWz0eBya2H1k0s4ODoESD397zM4E
hcwagtxT3RvIHJasj9VN+sbQsKd35llhMrlL+HXcxj8w2TfTsgrrNArrdGU3CjvgoFCJQnO/dFYP
rrv0iXAiXsxbDwgpXnml5oYRmUvXaaBQfmKr4PaG/A1tic3ag9lKdam9ItM7ZFlycTbF+V7J8qdd
ZMgHEf55Q2LPK9R8Q09KSk5Rf4RM5mwXDYOLilSXpCavE06HFLFBPQeNeHIUHu29wRAHa2l0ZQIl
SGPP4BZRBkWHWOaflPgWfhYyAMZivJYoMBPrFnQ0zIh7hZW8Vyu0faqv3NTFeBkfnSH5QymVnYvL
bjNxInUuUd3DIJn8XaJZAvcZ+O7CBIMayPi3DjRKzD+YCCbZqVnPb4O1VEx7p8vsA3WdhIYFy91c
8rj/AZ+gK0WTKSiwVt8HlCxiKS+f/XatJfAS1P2EtKNjRK1ixj0ewz+j0GV1F+LfsAJKe5heake3
eo/uN0TMbth5Dos4JlTvQ4cabs2/kzL6qAOqU/RlNxHmkG7fNMdGq8G+/H4SKhuA/q7tUjRlgTSV
Qdxm8Xol+6UL4ORJUbXAA+zSnoXnk9noExx99h7yNJ7T/adqxgpHbB1e+F2XWofmxmF+awKmynoy
XAKsjN0xjHadSKUm1r6I3Egxqo07FzVBrkT5CGF4VvbnUOQkmmmHBitO0IFxOSVrBSgb19Cltk38
jgYj3EarswDQPJ8KcgoayXFqqN26zduNzU+vkOeMRYekjGBWYVsBg2VxNFMmQqf66klwxUDL481G
TgN52YCjKA0N/iHoV+XiCVEX063adc2CfTCiOuQ+u6Sv/YIQhKvkbZCgbWNzSAmxuST3Xm5CuTWP
OF3TXKdXnBmXC6apEoSqvRYuxwYUgBssYyS01lyK8JlcPAkpB1UJEImlHyxwp6vdqDS8+hyz7ank
ra/Tq6j9gGif68/KKNefthXuUPZVt6IZI3v5D0WiXNXPau2YVPG09VAxdR/rHn7uSASa1dvmubzx
YoAhE4+Nhe7aHoL7B0BqPaaT2zajIcNw6QdG4ntmjreeQcSesZ0knaGxnHnKwDuw1OfCmlNKSRR+
DcIaUQx3gAqEER+bGkop0kVD25dCoKt5De/j0sazno9VgNvSTXugwWYu8KfLB8z/VcBzKLe4QjfS
H3laX604nB54FiihckjM+CPkmFKYiumITmlH4xECJrJkg4BDDNgKqsoGEqdLNYuBFkOyRxy4uE2k
eNVOsqAMjG6l3jUJdqu7m2Pftobnv/trEymrM8pO+HAp89C2aRucY7x8MCqVvkvuwVQqe7Qv/Veg
sed0lRtfPb1vzmkfo5kXlvwPcJUjRvYyq4p6iwA9LL6vqi55xjo2YtKSR7qKubdoFZLEAAhwjK0x
04qKc+KXCKTBW7Wa1WOjtcnI0iXCgT3Fezkuy7jG6jbVnla+rbsPGSNL/1zbHYxTTp+RCUjioRRa
36n8P1QQwWD8Y/pMzUimVpUAFZS2OQpC1VTwX7LKcyb76P1lu4XQZtb41JXUwCtuMkPJTwAbCL5W
hlu7aI5N/PXnsQLF7cZ8WwhBSjH9haWrbY2AuW3vFsiuLIbqp3AI29iAlSq0tsj5UtLxdf8Vi+ii
lJCgivaTum8/7HAjuKUYWqz2sLOfbJ82Xfp/fJCFA7bkysR7uLvV17gSn7ZBG3mt0XxN2+NBGvEo
r9cloV6Ay7r3FLtDNsyx868unm/S8u4Ru7oMnHtuR3cdr4FtIqVrwxCZ1p19mbNEtYpC+SkUAA3+
crdhTrBaCBNhDo+tTqwssKrllEHNoGFAQ07giaNHhJmCljNC3LwVMJCWvFuGmj+kNe0ejqjGx9iG
oDPee4k6TsPKSFMWQV92mfAfapjomf+s0XqyhHB7gtAHKdtbU4WBEFzdJ0m2EfPe7XijGFaX/P9c
k8JLiemFQbvQxB/jz/jhugJgF3khtZSwJz1jNOY0Q96+zqAiUCyI2SAdlRAfZBjx1CA29zdzuBG7
/lSlteM6zyMK1zIKkVE4PzEzkkCPiJSOPAEjjurpsqxRcNwGIyyLO+1dUJeJ4Xg8UEJXkfqRsCMf
dB4lhcn1Y5jcazdBD3CDKcnZOBohr7qE1QSHw6x+BtWXoWaSyCiosxjeN256PCTtguxFhlyarP25
3GjI8iTzBPjqNuFzQJeU+JSpNLONXNTdwsK+60XR0/wUy40rMTukLyUYSPIpbqWCbP0AnjFAFyl/
lYhc7ZnABg6LF1lHqHmt0n4+0dKSeE+BI3qeOeHpgJpsj6osOWqf4gnNAxp+PiD73PzCQy9uLQgb
nlJ0Ky1bTgzcIDwudG2DWJfCbHZO6lrdTmHfz/ltHjamAgcMVQYt7bDrrP8/xVzp1pldNubnh8XO
3e+bepq91WEjPdbpIbVBLDWGGU6cAjTGEcDguSBgmoYjkwqLG0bF4kBCiCGrqSYRhZ+1YmoazqWS
ph3Ox03N1ckNQOYN4dlkJxasZs58B+o+xwuORfHcFwRAHyUQx9jkcdcMDyVbcoOG1gDnDZx2o4s9
7CnyZlM7KuyzRDpVmk/TCrfyiAC2ZyFfbtE6IYd+5QLqACUNwIOxn7+SvqirlEz/s1waZSid3mzK
QNZ/Ex5+5pqhjjZvr22w7cfMDTbjBRbZHeLoflWNqiv+RMbltJ5EufX/FQcaaf8hgook/Av+ciPn
SJqdRu14qImhPsTv0HEASukIB1vhQWObQ1VQ7vkspprrhQx7sVB1TBt2GpFhy4oPvxdUpRZI4gp4
YJUNXYGBoIGsZ0ncOK60nj2McbdE0vSmpp+cIDIAcS+39Le2MfBeNLazoFbC6MWb7R0LYPDM3Rbb
I8rzYZFgVIDp/vqgRtYnTKaJQik81pHMQpGSQPjw56/64qedxGQ8jVb50yE4W891stwcd0Ro+DSg
DDTT8ldytdsAwsRoxkefDGU0DkpS3y7FIa4DKAJJzCtQyrK+8GN9F0abjXD+p5pGRyM9VeL8Iu1F
tCPb7HWaeLipedk8QVGs6rRho0kTZX62znVk6hsuimi/UZw8W9iP1DIbwHTAjsBtisEJCy8ft9cA
kNCKQUNGJ9TuvxaxwumosFlzFkUW1fYZ9trDLN83fZCjNuLTEapAk70IsYVIqnPx8QlT6s3Z7jz0
TEjxKZkX6t+4WUJyqXpfe+hbslf33zcYcZHkG+MSKLNGOiYH80NoxA4IYcuEg/hFxWuis4pK4u+1
lUf7OM52bxJNAr9cjZv17JvDKUYgx+TA2kqWsMUkaf05MDqG1Y18m4aqH6OEWXjtpH1DLeGtAz55
iYfsUhLwVyzEwo7xhVpN0oVz7LNTStteU1QSVZbhWs7e/Uwt9hL204npeCYNNkwUwLXUu8wEBG6C
KddotSzJY3sSbmdqVHCA3ACUj4lIBNQl1aP566bT8pgJpmteR59yuQyZDKdB6IOO3XQi6VBIsych
iAxriZcKB+pHS6rtpWR9FlrNS6Zd4aQkfFwlArXNKXIW/aBBD6hnwWLuEFQ8rEkfnBx96WV3cnnh
vQdNIf5t0OoEk/FyP+36apnZ9JDkkHgY64FlLstv+mjTU0lh/34kXOEcSmE8HhtOaZFTB3f2PzxC
8Oa6Cm/ZWCT9ONUXmEpDHBKYVIG/uDcCUIXtpiElqGRMqkGK0ZPjJOe8lPMBPAXCWwFCvJif/b6G
ylIzrSAslVGSDOReZ0J/+XAz/ynm3TZW+BF1Vi4Pv+WtLDXOpFG/9vZWg2ggwunKBReZ9EoigNm1
uEfA2DeKWH5fi8T32NU6uYe632oUgUltj5r1up2ynz9oGEEj8muA0zR7f4XdcTjpHBg8g8XN2FEU
TnIz/EKphcHS9XL/L+rtOmNsiVmjLRYmlSmmZkQz04jnaR3DbrKRbflkG75Jy83LM8LBZlVzTTTp
nk1Xnw0b5drSWuibbrvm6mIykHPTl/mgmoTIwpau4nMH6lom3pLBmS17Q8vB7DSEl4cn/GPHVkoj
5AWLb7vO3bbvzh60vAA3yBNkX5RlCdQ5DfJAITp8Tlzpc/NPUIfFdLy9Hsm6w04ddOpGD2ejo7zh
Fcb5NfCMe7mAa4NhMulpZwwgMThNllbh7Isl2SHeWUaMtb1C400YoKsHa+4/TYDs6siNQ1nI7wtr
7ruJg2O3BYmUPKEYFLLCDMrBxulu0KRZKCrLAZshdxdlK5YjMdv9JP1eScDGC8FLdet9C3aNjup0
7Ytx45MmbCSaquiS/9uQRngDh7m+S6rd7wwVzhQ+kg6P6P+/7GadQNmInom1JuGeLCkehCaPzEPb
d4S86abyJtXJUNblV/7V/I0DBwsFwtC9its4KPB/Gb/ZKHCVqVu89DXs8bGfiM4VQj80cufnxqXS
xfMSIzKiNqc/upuT7Hz0Z3hfgOf890BFo/Ks5bxRYLNcI6zTEPKA7bW7ltem4cIHocLnWl5k/LGG
AO6adS+wQAXUGRTR0kJQWJ/sP1V5PRys12cB6kkVX+3HvWcypQulbFcdJAKGCA+78GP3OPRcR5dV
77lo4cikf4gDKuxDH4mfDA300ORcyAPXCb89wnbJXm/7lzfTnCahLBu9PqKKgyk+F5ZQdt+U5P9q
3ygGm50pdn52yxwWLdcv/rCpb5RmT+SASX7UoTgT2hid/xxo66v51QUNzTIsCWRMmlwfdFx68rWS
1BiW3Gu+rNKfUnfLSEvH+5SceMynS/OktGH8YJujDAWnUCjQ4jiytLZJpeeK9bKFz2dgZqMK7HJz
F1tsvMHBQGU81vNdPaHQC5nlXIvEu+ySQiEWxbBqPiM713I8lTli+kmdjBc1pWAx8V/XWVxJK0R/
6mwsH6CuKS9DTt5aTTzwLeZ7HIoKsZgBJ/yR5dbsU7t++tJoShq/XQvmUQAym8JZQLLKBOdqSbVe
5jJaM3YARENUXxp2yZ0ZUWOEJ76/52/g+SpO/v1HDCQl5AckRGWO6YMHrsxWJ9cL3oGgtcjO7FnE
tWr6aV8B1aScPYr2O0BbsqP9HFpPs0IdoLCJtx3igomCliKaZ8a4j7i0ndDlnHntsHdGkTFQ2Nzw
6g0cEnKVAyctOzSxTO0th+CnuPDfn0ll83ggR3Nf3aDtO+ecndDTVH+HPhUmoEUD5nDOMxoLnZXq
3yKQCQOKWA5OkTtnfJm96Gi2MEp51IPMm3ueoXx/h+smrRVA/6qOWqpc1ykjbM1/lvZBGYsu/JHm
hk/CIuaIaJAOoL8ZRP7cUdmhyVhmmDa1h4kr+EwZcxy3H/qs41Hr+fdRUPkVA2KEQdTzsZKymLa3
dKFrgX4vmzVwjqtG4IIHv+CK4AZgPQZ5AG3Ue4e5Pu45r5RX7BkgLhu6zbyT7dvuZZzSgbOBOHXR
GuaJKqelUooeU25R9QDKexYhaXAKvgT00HYwnXcO3F7vik4gUS6dI+AvWiAKLfxDT1zKbE9C2okb
eLY/Np4NbpOZGRdl9ljGv92kT7kJe5KD+6FzsfZTj2gpzPKBHrQmAgtFlOwJvAW9f1QpEtmlI/sg
h4yB1DJiNiOKRPFYHVfzH6ovFYX7kkh8ew4l9ppzMyGwwBtmg51t2OJiLa8ewAKbNJ2qP9vLSBgJ
Tat50zqrygBfF0lxw5PWbwS+kkGxiQKenV6m1CfCoi81mAo/rCyevqjqkVHdUTDv5YD5me1WISmX
7Rbos7MUnD3dCASY8vAkeVIbMGmo/k1IchjU191xl6QvcWX2GAP0z5Qcsq5FtoliXNnGwz2w4FDu
bb0c+pzPeXfyvPld1sjISyvS2neeUeVK3nlQzf/Jz9gjDXgQs39X0UkcioGxUOlgvfd2HA+sNmmC
TTB6HsB2/0RGA7iakdAwaBV124ul3disz2pGJleN8WHmdsAks2xE2CBgnNrB0gy7iYW1fx8GDZsd
HeNEDwJ9cppW2Cbpr/cqqVI19IFFo83k2VVdvDYm1l0MzclLbxjGIpvYYVjEFHHydR2NOpJWwGB2
ZeSU0SRV/yVXYH2F+VAZSsOPPk08ykNHiaELNSElgHZk4apCFosiKEI5d30Pv+EZjpddw8ldFSty
GCd6moq/mfXiBUfn10k70FISYkamT9EfufJb6XcFtbomNL7br6uXw461uxxowcfBdT1jL8yk5dYL
mKOQmtuGKAwu06nXs5Wzf5qjwRSgq3F1nA4wkLPMsVJ3C20BJL9uU3QkbZyfwVl5NkVNKNuWZaBE
lZR8UJqeIbgAcrP41EDga+2Ubj5Y91xHpdVKHlbaOUFcXWihC4G2SQNH1MK1+xAROdL8BOhO9PEZ
YsS1dVkXbDK5LKtpf0EjXUWOwmAY+NwVNzLJB+AvnoIBvdQTBfKxv+bSmeWNTpEZ3mIQYZtQZohN
C2X9n8dop01e14aRq3oKGu0eKUccnG+xGex04Fjz3iAXJseb9dSeOvv/Ql0GPy4dtx7VdmEsdOlW
frM1gg0zGvCnWMt19A04x22RYtcU9TfMUk1yiAdvtX2DlwHxACv87a7Zlr6Y1CdmI+NggD7SdpVu
cV1//95pskhYgscJl0PCKAplRSZd3AINtrkHEATSkwvRVSa2yd4jus7Q5FNxKwmjSYO2twX9DIQU
/CEiWYyJ6OUa/NweV2AKKsMWzMlEOiffMOm9ih6V/3U7Ae6L8GlAL08ekAdQDp7rG6QOdRuGZweZ
L2ClvfVkv8jAT21OtMZkBcHUagxaJkdVhX30ykKk4p6rQHCkIAagAr1ZZKFJMoq92XVSXy5Mj8oF
luCZM9dSp8DAjJDOlltKJ5/hPkfugicHDs9a9PY3vyjwJ1RSX+G758Na92mU8ZrDijmLM0sMy7qr
fXPwkJMrpwK88vhOLATNYfVLhOxusbNF4oj9bW+rw06dah3UkQEFCpDBQAeHOFWc5shPlGSFDqBx
c4gLetzTCuCJa4Tae5EoFN97PgcQdnj7QXeQ0p9FBcIo/hd5NC9qvSPrHym563b9Et2wjsSOHdyh
VoHmIm0OXRYhryybZgJxfx3PtXdBd0RYdJGGWZkcxxDvGVQYOt6KdQYoWBQl9pPp62zeILfkncNo
BAzge0WZ0ZM1LYwAY+le8wNHTBFpE4jLeXNbru6EKrXGXQnazJmcgERTf7zyUwzQNpnYH7Mjo1oL
j9jswasDJiqBRfIgIahRl9Pfr/It8sp0iWBab9HNUTNhRrbr0M23szqn7yscQD8iK6npCdNTVtND
GNkVxlpGA4nBRFO9wju2BV7roO0uGVovukQcbuEeNbcBdfGCfW8AfuTiQww11Gr1ndysMmRJqrh8
mOKyEmu1CPbM666PUbdkFRwtvbV9idVFVYujWxsxFFNfbBOaEQulstyUkyUE7bTOy7c/7u6101pA
1zuop60MEC3Hl1vXmFydoYMOsvqQvCHKmfcvQ4WwNfU6SmXAMnNhYKJ+yr5oluism29CJDVv4Tzf
fUVa+1OYje/wj289In84nZO7bi+/Kw2FjsWd+ueJtVl3sgiW7D9KvlRJd6ElXyIW007h+v+t9XcN
/S3rBYUIHuLkyZZkSd2wXbdbe6soAxFi9QAe8vFvCcxb8ohxDDVfquv9HEioeitLgbCzpTxAYhLa
CO1r3MM8V7Tp0BSD4LLYTa6NglZzyeZ00FcuBWYFNhMX0foPQ+gDlzfF+L6BNfdF3HkyrPpDZuOt
xAvbqM7wKA2cATTu/2qp7XAGzo2HqmOSPuNlNmL+2ODlS32hDjOpJHZjGdvTIuPwK/yAlm4nUoIT
G7TKNbSymowhleddSWeOCydBb4iGoaGZmGcKOHzjX6QmkSOQv4b/7XCCMoYOT0WdVdZGJkwBDpEj
cNWhDq0V2A/RAvQ/48H2BW0mOPR2/SRE/M+0Q0TngO53Tv0yj3Y/7bqdsc4wWY5wcHFXjulUDeSW
5p78t+NpNwbnliG01CrCqs6l3+5kc1zN8xmDZbovZxdLfuk1iA5Soog+aJm73nG9v8ZVDQunpzA5
3D/D/2dK4RW+Uqd9iF+LMvw9l7kCZPx8t4N+Dh3l0IsM7cflZXbzXdx7IsK3RvsQm+4lJnoXcU7R
EjPtPmt0kFjFYaJpOKbolwJWhwKNTE8X8h9+qzg0q7FA76/mSZpRVtx61hzvgVAmlhCcbHy6Oxll
HRJFtX9L42LrwPkJJ7EYIXRIwIGr0W+sWpNVYuZk6FMeemUQjmRF0HXRxGJBM7vNcKQjtDTKIt1s
IBSxPrlrEpGXJU9okJrBPj9HskPjAbnP9kdRwlFqdzRSzp9/WBWjtVuFv7jALdchs3v5XhJ/i3uT
ODRgTZSF+MgYbziJqKsbHdAxLPX2dPv7YflQXd6zqLyKWrEYxyntDUal3/mEJ8aCYT/wG4zqbhB4
fHkiJ7Y01eg6ywHZ322uFXudQsrHHol6VZLFW6YjhUWYC+SaU5+hPNaWfXTmjm7u3s9jjujcggAo
HZriX8O5PTKu1GmBBa2GsNOuYoEqT4kCjYhm49AWHQDXXs74aZfz5znFugRU4kgeTBxUgq/0Aw4d
kJCmM+J+LTH3DL1lHrB4C0PLET0cSELm/hFFH0ZmhdJCsxpsCggOpyXNdujqffRVBZb3ObBtaniJ
U1GKizhElpKapz7gO4LTP495HQrecTw9b3yjFjO/FGIYW3Z+78FdA50rD6mDq75KSbKFI4Fw9h0b
3Wilh0krEvKZZv9aBV0RU2XTqwxigYQxsHBI96Kr92kM0Xob9eNeZiHbrYegQWDtU0Ko35TO+yoB
yyAM9WXcUNkjtROIMyRe0Km4X4dsXfZJZdNYHvl2sb0YqMAvYAxtT/UeQj519Oufc1da/rRBwHiZ
HY4ZQZZcHirURoX5RS5AQ5mjcqGGk95AyeHLMnOI7qYsE4RxO+iUwjOX/AAtPfXhoIHKyYc9tUP8
n3QPEzK8kxp33FAvOM/9VnNxxWrNjOaH6D0zS3QFQDJxdq9DIQmUhz2t/7vgA5BQSL/n+ZWFK/J6
WPAK21n0yGYw4pDqFnQKBrPILyPjcApYo55aC5u+lDQWTiW4cPciIza3FK2R2Pw5z6ExrdjP4943
mYZCzlA4j5RegFKTkR2Y5Zk5oWy9j/W9dcyOzCRLkxold+wlBwqNPzcMg4UAI1VfAu+pWnk5Vrr2
2RHZQi92N2aJXJIlcdSU7qWwUmZjWCZFzm2SVIy9swq8xLMZPT3FdubtRhW8WYHyw0k9v2hq/I9z
7b1QOe7h+zZpXux12tDDf0TVuqHjUnXM8IDmg4JkO9xNhKGSkxi53LHqulFf4FjyyUc1hnHlHq3N
NEy9MTZhiByQ5iefKrakjWwlc1y4krvM5QCWWlS2sGXPAPKCLS4v4HXI3eiR6leXf8d9p74T5s9B
j/ggyhi3G+PiMPDAHTjUrABVuR7lD7kRDaj41a306X9JJ+4RJ0ym9GZeDSotxkKetvf8kqYYxGNp
Sic31fNPsswGsqHse57eqXoLGIg4/Mx77hW6Hyhb5b4r1TYqPr9HanxzO3RZ6/HoL0detjHdGjIl
+mTbZVrzTiJ6asmRJDxVswcBUxH3ejbdKaY/aroAzJtPwoBMKycuyye0AGVb7e/hCTP8ODeBXKBt
FiheYG5CFaxjggAnz28td71hi64Zg6H5OgB1A3fhVIMYcsns/S65pSHC3cRGJDj+5qicTw8EYRew
VWsdUHoCnuq6Zui4jYn+EnVVitz6mZF/OHTNl3arS5oeKBj96IWY8wToHOf2vekxi3yEpa4BcPqX
j0bRlzWrPzWeOI291srM54j04IXNO5feXJJJQW4t4m2oqEVjNq44CzdiqHzfvFumi6pRNLtFOEY8
hyR4VInCHcrzRXZqnNP5aVpa4vq+/8pgNOfs8Var8ThekFyoQNI3sIwAkNAZ1ftegQO3kyXjT6zy
qFxDIZGtB8q5AmjcKdFRrxVeAD4ErOGcVOkm7tA1doMiscs5B7bRLBuDqLv72f54iQlG/D6Z+7oc
9ydNPnUbGFlcB8g8dPt0JRNEKcC30exl6wtsKUngLxdtSjIzmfWgm4FbCHS7oloqc/SFxJSRTeWd
d+ysR+uZQfbKlVDrZeRltfopuZhRdEVGGINy0C46wYeY5Fw5sU5JPOR0V5If1VK2pB5ne7v/5TZ5
Ha7cQ1DghsEmj8iJ5yorVx6GZxVUwSXbsRk28RSeUJIswNZFv/XFVt0ygQIyWBHrkRjJhTVE7a7b
LcVlIK8V7P3+oc59NyH3pKZJMuBr7hXLBHCywZqwq3nU/32ULLNQ5a5CrSO8Pvf0YbeSXh2y2uit
hRIbibWWDCjtF1aXUVW7VbmVApHyXZQUYBYfDlqCqPyGMgKiD+X15JUt0yQ4jRP/rJ5Yx+E9oPk4
+HeLdi0Qp7J8ImwWaR6qK12ClQu9piYdy14EqucRoF0VBnYZpWnvhD4WC+6SxZKLQ4ZCtrgt4HLM
4CiNPl/w0FlUYPR2D5Yvz5rbpV8txVo/9wmVMH6LaxnSEaSTCDFeeGbNzz7oL5AQn+8pTJZiJGAk
O2+nF0XG25hv3T+MPbMhH4LK4nKIWMho8J876n6Bs9CyfzzyfdVAgV6ZFoc8DPeOlkDpC4c/2u4K
l6me8SpKCNbU8+Rx28lsg8AA/XSanmw3r5SFgilPrtgH5L2rlgFRs7tzNB6QEiVedoKDr5FMaXcM
r4eBJIx3Cywkiyy/EjqIloGWu0DWF38j5ps0NJavSPTtJRl+5cLcBgPoSxkQDwu43yBQSVj8ueIf
hv2qp8LtW4c1K6b23UnGtyO73OF0Zx3qaVyRng9Zo3Wx19/wDgxrmhzO4L19ZdbVFUiSdlBi0+hS
+tgani6tpE7kqhjOiBmhx7TrKMFY7uGiV1Gr8MDHfAu/4YxPo3vuf3a87UhY4NIlw94IxdYEQlPl
uyfFhiKOVuKuNeXkHe9IiPFju0l7YesL5A7YX5xK1reLTy0qM10YXUtZ3gZ95T60Ci7ku24C7Tx2
JBXvXeOM6Srtk2xmi50Ql2L6aXRiZDPWoz6WaWqyZjhqzi1QuSGjTCjR8/KjDpiJWtjVXOwAGzDX
MuvAd5f9LwEhXvmT7as31AVLszaTg2NiaVylGu04qH4A8T10KhPjVcdpKl9X6esDmzg2BlTXMypP
YOm18CnGURGswbs7dT/1eR/gRZR/BeSu4cK3cP/aF6WbTE8vxDBmBIFW58TSZX5TRBYCD+/p7ya+
6KdqL4Bzpahp6x1XXj9Mf8vKpkM3sY+SzOPJT3gBH03fo7Ssu0bvriitAyMdQrrZNbmTL5VSzrfE
jIxjfAJVaGPSuJi3L211hgdgJPzsIlwF20XDH3RvYHxe6zo1nokS85Dpw7xmW8cLWL0nKMnRjQzV
tcPbw6QN0WwAYGPFVJW2OLLjmF9de12UKnRhqwmqnr9bWdHQsxrn9I19I0WkUeSAUNXbxO0D5gzi
PjCHQxyD+kc6AFe00w0OEmqHujRyjJPJnBB5XpkmOPTVQ1Wq0z/GmECBfLzylSiDahKzjWFl6QOZ
yT/PlZ6C6QfFanmSwtDv+fwH2BIfU9rahVkLmLw7vMtnLtqdl+rvk9k0jtQOh4jkFUAKSNKdrT88
iAd7AkXo0SFdYvBcbz5qqtnErN8OD3TBl+7rR0UhIqF3MaAVzWAkAx/b6lytUpq/FoI5fnjwV9Ab
gXOe5rMKDF9v8Z7IPVp5KOva1aYqdexjRdNdDv84RAtigPGZRyQfUUyVF/L36igzvEzIsZaX6EX2
sQB3OMAtQD0j2t7n1sbuHnYSXjSNzLT0o8FwMfJV7NspmXKYi+VpEVM4WiDVnoRweYK9eniP9xPj
FvSceZuPKlQMhAqaGJGsfYvKwY51unCwP+TvQFbv6YmTNB8NhmPTZRv/uBWlUkrkFJna5DCpo3sM
kXjvq4Fn54N1wjr1WTWNhtjR1vZyqZUfdc1x/GqzzA132JO/wL8XDx89Dx9GKirOzvk/CL7MM3uK
btY21N4TtwDjV8tA+Du5MADyBSHvlZZSLAlf255E1ueNQ1THgJQEwRqQAMjRZxwjqiNmxQLL6cVb
zDOC8AA7PFXUiz1zAKvXo4DXwvRyu4GnB4BoRmOzusNWXhTim91d77FcdBAAoVTJm9o1St1y50DL
/UFiiqy917r0SqPYlo3+EU5kr3bxLQM95OoD0hc5Zj+bDEb4gImF43HLiaDZkJNz1fxfUyKPs3e8
yfPQHazzn56IqkJ2idEXfKtKxCKgje8HVlmztIHDkPHJ+xHQPt59KupE7kpbRvIftjSQZN51kkRQ
nzZVBZB+XItgq/K41Ul3bKdcFhfhVhIHv2bIUNr+RJJa+NwuUxIf50+02zmOmXl/81xlxD007tt1
Au73vxgX1sK/8OQpS2SIgKgIa0SZAoTqBddUjrmJboJ/vCBg7qZ+2lzGYPu8M/1BDIQl/9x/GlCm
caGQVz/pF/m8ML0saKUu4K/vex2JlTVDlmLKZMfrOxcmOsotWrBSM/k2LhmeiOg4UPVy6f2UxqJ1
9PdQ+FMuXcYm1akYmOvTSOzWKNeziP2fNHgtEZn5obVPcI/Ey17widEgKInv4WV/zU1pZORWJg6n
2lIpWMVtr8aRI6s+icHNsKkECoXufBWdHTGpYI9eOhK18fMVYK5wOmKrqTcXdVBiruupWkd7Nfjf
siJv+GzUc58r2+dbrJ/Ndj3jDJLCcDpJZZCD226exEw7x1MRYenuRHLocYcRq6JFK1iJFdkenK7C
0dk+zPVqBSOXknFf7fWBIhKWbbCzB7jz7WC8LBtPlMDQDkz5b6BHHnzPPliHxPpqIBOIZIDdVvaL
bRdQgWwbi34paGWkh0T+EWl7urIGsZQ+YUY5n0pOYA9Aa7scoik7Vv/qCPHEvLlUu5tPAFqhoT//
0XbKaPjZJNjJWmzv1GTKHufuxFUX1986FjjHBAJPbIijDSYNqlaGpndtNzP+oAOysmTEd04Dy4ma
gUrGmIooMMHVZAZA4R/lpSUQS05ly0wsnlyMTyPSivyB4oqS1l8mffeWVLaAKxOxi/CEC+AZ4Xdm
FAMQr4YoUfbtV/+lXxUwO+cY9mEP+VrCHCYQLql4n4KpD9r197E9YkqtuaiyB3amIgPNut6JbHLK
sXnffkXMXHg3GUXtDZuhqeKDKrnFjSXEOW9Jyfr6ja/t7Ulq+crk3VR+xnBX9+b/g2pmeTU+1Ps+
/q3YEFIkYXi1r3Bq1aP+CtBTVkhrFAl7aS+ExYJVI4mTPFx3yhloRC6xjmNwyJz4pjHyGTrEfj2e
W1MPkrvJwAQe5SqdMjvUp0EY+J8/pYHhPbFnOvoCGv48t0ImdodXiwZd8Kcyagzwc0IBMEGRLqfB
3C0XorLzUckpjRxmXBRv9sWF6PPDnB/He3Wd+Fdgu5P/H/MimRuVr6NhHB857HXQfRXyEwHztZjz
zicZwDpa989EiwsIaRvN3FB8nRPUkm+3JxSC/b8tNvt6H9B8iseiG3/jdYsvxjOEy59DxJZfH3cW
WfaLJriKGY2d/wSqncv42SFlgrI72fRa1kEUvNvT/d0rH34SbcYVZLH/ByATgvZx/C06RRWmahtx
ZZvTLRa7gvTm7CDboD/33cB0gZ39AGCbmpgUy2TEnqBUkW47Dfc828DcBEPOzFdT9x7m2wDa3BzM
uJcIN/azBrVyGgjaeMyHbQdSQB35+1F71rHiC8XfMzAdRYgabptwBhVCeeFeaf6r8tDnmv+kZerU
m0r6hrz/vaOSNjl+ux2oQ5H61YOLwmTw7tozDhvCzomX4BEZEZQQC5zVyE4ZK2L6HvjeHlujRfHV
Kja+n3R1TSQiqqBv8t+f6MW72kfgXfKQsfZZLIH/u9UjHB4GS0vSm9WxDi+m0wiE2Uy2BBjl904Y
rTh1rpBzgO8x/rlpl3+P4oYspK8h+n5k/KYyRg/5IT1jmMsB704ilY3duFHzZ1XBbThyymrFWa/A
yUIU7fv75QtUhftbg6ZUO4pIB7hNZbU1nAIyIJm5+S4WrgqrMPpk/fESsVITPVokHp8XCOZlU9WN
5jEQt0lwk229XwzJSu49XZlv8fY2SZmIoI9uEKGQ4yqtHQUoRFsYSkuC+VojIYC4fMRQOr/3Qdf+
uYBL8/2Dg0EtilKPus+5/MoeUYxCBRXNVseGbFJPe2gq9UZtWnAB17UxTZvS01GbdS+Is03XH6lA
N9C/n/uIZRUJmCnBNfcq+ME3++71zNpQbmkprSekgVqsXk75QcsJEzQDdUVrzFXDeIBATpeXqP6A
OjUWlze5XPjW1KYhOI90Ip03YXLpd+mCTbSqFpWP3Z7S9mmZRGnIBaz7FkC/gI5Co1DbqlBeS2oT
YdbkEFUoD3Ej2msiR0aVbJDw0YWKgIQn9xJ8rq/3tpsaF5qmlHUA2uWzxgCqtdWlxjDj3ecP3EJc
bzZQaMpdUidF3rmBKuMaaFEk2A2gOkwNFGSerWL2YsgWQHGyL0mLxMWVeBHPHgoX8PT/XCMvJtCm
TJcwgOUqN3IkZDsz+giKgHMbnf+beZLEyocDfXH7vaBHJNJ/Z0tEE1wA48L9J26R4rwzqUf4DdBT
7KxR4XIDkjoLHJ67VOo2UDCwziOMVz+LrtUqZ6jYAMduU9WorPNLtkAr3VsOiWBlnZhrwnOyT6lj
w4j20weTcQvQxhRQRoC1FzZ/eQIVKIDCLsj8MagDqG5Y/dJT7l8WjhEYv5HtEOygp6D4vGjxcZXV
NkHPbm1kJuWuaVfpl+IH8ZhZFRVfzm7gBB8jytw4ULADS3KQR0cwqrGLU7/tW8fKiAh+6Ga7Pslo
3D+BHycZsN7hre9Tszbl9mD2Vk/fOSU47VVJjXNs03oViYOMclN1Mn68Rlb8FGNd6WbS+BNMmwRc
jsNUpi6Es/d8ZWxqHkArXJGzRA9YClho81c6PqhgdEe6sLTQ9LqAWiXxKG993gG4jP4T8rMrfz2h
BFyWd+WwQz4ro6yYsio97Pmg0sshPtqGKJOzRAmIrvV9VSgm8VchckdO6iOHfXMbH6io32/MlOs8
XG10pDR1V3/oILcsFq+o1DbXx/+uFGloi8DoEr3WiN3aqu6ZewJVGlaSpPducxIiyq0+BDpq6QhH
ccUsPSKkYGydkWYp/DgSMBWubzS0ya8nPLaxPOOwX8Ox5pzHbsjoh0ScgI7kxTs+Y1x4PiOa9sBD
3fk/C76boQHtXYHS3o2wv/p7qf8yG6OPPRAugsgHnnzztC8lvmauiyQnu/JbFM8kcTVO6OowUIgB
+EYiwj3RzuE+4B85UehdFYpBWdIVhnRdMvUx4R+X2QNR4NkbQgmTh99dbwAR5W4Vm5U+35Pcf+vd
ah20qSBgrN/RICYC4zSRDWaE8DmxOlmQvn/wEjua1gM7j5UVtktKfyljgER8+mglWEAenEkR7tZD
WNTAVv4HJUvSQZthf82A8S+UBgFwpwTZlYizmiruQHVwob47teIRWpWSeYhDiutlJClnuN1qof7r
sSjeZNWh9lWdKYAxih0yY0L5ZEtnrIJS8GnDO/YTbob9EOr0hn+uklNQ/4QBUSrd7DikXoQb2+U5
d2lrXI+x9v4wdrxcyTvTiQht/ISeUquk/qjpOdNvkPhs3DQjmtIifRYMtmEJgJvLa3LcrV0xg0uf
YuHpnyhGOber735/qfeSCdMFEb2rg6ywgo66a/DxjnyRcbSvu7ud2QwAx5ReQ2awcgnlVp3iOf5o
BAsbySv6aIq36yHviKnDpkkHwlSyfYZQlFJEqVID112Hdd7qyVHFz3bKGChvm6EnbZMpJR2Bn/ZS
CsJGu7X+5JET7v/GHGED6ZSNwKlkqCu6TkxfjKdiu/UFPT9c88H64OwNwOAgoqqfNxoio53ULUcA
fa+e8/B+zAe0+zW4U3/eqckWIwZ4nI0+rvuyo9R3dcZO5UwTSNToEvucs2znFNvThEp8VePgZQNU
JqxGbJ+sN9EOeEyUQ9Ump2zHrIRGWUI1uf8QArWq4X8qW49Wt1Nx6WadHgNSV4lRWLqWkR7Ugp4v
ob36m+OuiSUqDBdjRCBpUqM7SMEx9h1n3PtBxyeR1GQB6OqJPFOfOL3w6Qp+hnbx5YoKW2Bi+m+y
H4s3X+KWZFTKECNir77KN5NQ8mtQTLzw98EYVYMvOOWzA3NpXu/D6h/yCpvdd8Sg0lgbcLKbzx5q
+fnjLJUHIr5W6M2thHv2uragklCKdgdXdpWnxqUV3yTw22wY3D2cXiQik8QSjSZXn3sPhmtZEoIU
RWzBZJ07XpMrDQR5R9mNnAP0P92mJ7qJ5B1mkG3e2Mqc8/ijPZ4sriu77ADCi5BX5CUgG8NSbkES
PQvqTJx/R6BoEffHgj8dPPlbiQtXPGk6AuZSMG00jMr0h9eUO4HHx2SbO0aasOxJpjBu/D6HyuHM
QWnst4CABEsMuFi6rtG3vkdtTh1oZj9khx796RC1mHpuhM38ARRuSLmHtI+hn2UjcsNR+XDlGSYF
n78mKQxiTUWgP+erHjFcup80bF4SmandwFYPPCqhkYi1/xReKkZeqrDD7fJLXVbkk1A5QFWHBIpQ
YdhKEtFU4bOVqvH/XzXLIwj6Jjys7+RF9VjzyCe8mbsRlraeDaUs7+VqJuJ8bPinWVRXhXCTsZe1
yeQTmhl41rl9pGeXOoUmptyTJhxS9dIi8wAZLp1lTbI1ZvAhA8CIToXXNQb3JwHcNDyLhwmwJBbk
dX0iJ49y0NVqAoa20Ox+BV9ZfgqvUEXuGiCM95EGK1zL1V1JhoGFaNYqQ/LobF8dAzfaxrMN9UHy
ajxKGoI0uCDo4qHaOcLoeK9Yd9yEm8ufjDYqkrqq5w7qOxNJZ95WMFUwNHi3hJDfPCHqr6GlJr0/
Z5oOeQZAdfJKvd2ltPxRoUpvQvN2CdSDTn1sT5Y1NxckvrBt9EBzSzQ95sZOynYr74EtudnBAsna
RDHI74npUuhkREBmx+g1YYsv7WDQjuMSLJ7sJv+bSCdkobY/Q0V3+C8e1RB20F+ocH2tx8q3DyHX
K1iC9lrTHpSB8E3L8JPZLvuzQyYwL4hTVBGJGS6hW0R/8Cs8vxJvGD7KbmtP+4umF9F/aaGnTXxN
vQEIOmHFpPLtx5EJUk/EbPo2VzoLNTcpqlMAmUc2gp70tuKEv9/XJ0E3O2/A6vPaN4KYxohYabRa
VlhroYsFp/6/l3k3fiW0pNqMinqMVo/wRxDTN40H0U2ucqEMbvPlW4tCH/gSLpUmxzrk3IJcmDzU
BwIkctY4arsnqJCTFFAMt4puDfC9BtM+nsb5faEqb9sx3cpq+G3ee5JTApLLPKowogMyLOTfFs8L
f+HtGBSLrcd89A6nS/itoctMNhtuddZ5RWJrUhDXdP7Yl4cbC4ssSM/HBPftAUcaEKoSxtGrONYY
lYsJrP5kuRL4nKfYpnpYLGrt+cRN27RR9zdYxN91swB7qbEnANwT3OBXek4cFghysB6HCC2LIU9o
bcnSDRAtd3UvgBQJP4HeE4EZ/e07dfydjmpetQs3T71HCkP8P1NCL972ghALvaqV1hz4I4TzT2ow
T1Nf5nW2VhOfprbquBn5QrBmwHmTvdgT0wu0z7ER0BwnK8CmuZ0ke8YQJGNc4YqZX+QV5+1lzdDU
f7Ws+xa5ciaoEQSmDQPhxfRxer/RTV+ifp2QIXuxdNhctnrg1LopdFHsp3eklrFMVU6gz5HOscwx
xYxGXTlTmAVSOYvXXGCcIuM8Cb5r9N1qCJijZrh44YvBiSk5iMLxYsU0GWSBjV6xrSU8taWFVvON
CAqNxkqLhK7yF2MWY1/10HLiBIq8McFjMPtD//fp416/Sfe3b8IQ4A8L05tDU9AQrpQ6SGbKbAVR
PXNLJR/YCu8UEGz5NAR/HedE0TyKUiOPn4cgNn96AX/sbH2Du6dXWZ2LgOpC4oYqUSJtctBsaScX
YGVjTcA66RLcC5R8kM0fQgIrGz3LfMGFn0+bo4s6mhWz6lVGUX+NwwB+1G2vXr0BcIYbAOhKU2J9
LWEVvbNZktqvjFXx31yYu1PsgRAiytGUDTBGZsLeP7AWDe/GuAC35chFKI6hZaJ/y2wp6VEJ2JmS
SGwLCB9eAAWEYvqt0rojWWMPWdApsZvvzJ1YhDgDldX7mkETEkqwJgF3k921EL33VolNoF5L1YzV
cFcUHQNQD4eMPzd17sihYVYPXnzCVQe0jZHYYmkSqxGO63wU1EL3e8K86XI+fxdcnX0+CXt8/G+t
EPwoTm2Raw4KfVpS/+GHnCoh0IUoWn1RZrfzc44KHHT8mGDmPRDZtYsi2m+AM6BhZEeux8sSr94z
H87isi7QOH0N8e+O+9CTO1etJIsbaFBLwVzl6SB5XKOE5X9Y/Hel5yHgCjjtzoCA678uJ9c+P3mJ
CNf6+fIPkLVVeWfDC77MXsBILhUZL1xNfwBaVfqQsa1sA5G4cDTKiUM8bFmkRbOdLlmYeX2XXJjP
6Ov5q5pRPbvdJcEQqZyfsC0mfsMMN4g6VAB1GGSBUg2SO/X+bmrRQp5b2WAKktM4Ti6+MJRhiA0m
nypZiAoabw3WYyfOpXo7qnyrpYe/hUDn+G1H3pXsrwVwC0WJcObadI8yijgHLIQpGuzq4UicsUoH
0XSqdFiBOYn9AjVglqaiUKp4/rW4vvnVUEmWvDcueY3KVRf2CDu6tKiYh9o+miPPyxWS4llciW/5
ppKoeISe8fQo+flr8LlOOlosnCDIs9YPPvKby+dOCzq0Si8WZZRN8U/mN7/Vg0YI7Ktjx0bJfEEN
IwKHq3tOT8Wci+kzsPDDdWl27JUkUXYddRuL4a4Skb7fCXUm2pfnA4Yfs+fVbt5SIL4eKmyllJXH
a8PCp7oJGPn74xsAl9Yrd7045Sx6EN1lrLZjE45vOyCYqGUN2jD1pgbnJdeo0ZwxoLNboh56frH6
oW65/9hZxVrSONoB0gVoEA8BADq2vncG9v/xrjrvkScV7fjpXNfnoGTqE6YLl8hYmmxHPvg3Tqnc
LCN5ahQldGl4DB97tP4ENmvXgpLuEXRyPxoZDBPWysiCmXKoXpNqfk4j/R4rAnhf+HyJCHlJ3qfR
IiJWQWltd4anlFTLoFpZj1Tai8PBq7bhsVjIuTTXvARzqNzVA1C7Bilx/sh2eB8rT+HOR1oGZvbh
qCEEwR+kMGrNnNJZjcRofBLVFgjLuLEEoJGePdtdeo+9WK/rc9MKXZwOmMOg9ps2bjT9vnD/aEgL
XtqQlg5RWDXftCgT04/RNehQXykzLh4hW/TfaMiM4od0+x7Og+QUex2oiu6Ka2V2QFDIDMus/Dud
hPX4XeQ17RX3agI2K5ra9adzygRTQ699ypRnbqLRWxkZIKlK+/LfBIzz9smLShiNWlLrPw9BKn1t
cae+pXgB8chb2ZH7epaOsygOy28mVE0SZWTpEqDHnePPzNGBV/qNRj8vBVJmG2kOejk+s1dGRed1
+C9i036iKLfe8JkTG/NnDr4BCI3YW3BAR2w+kCtLaYIVIrUml/H0Ht8ThPFrGXi9HGRviSDfplwX
8lzuml3ky+j53PjR/CeoyJgSLBOfFIbR5+ux8tHX6vROvadllh0xg3KhpuMvkRREsrUVyE/0xxfV
yIEjFsA5qnjEVb/9mvqpdfqM2xzpgRnK9BGG6DlwAatT3HoOWSGpOq/8jzCEfKnV09CMRydzuxRZ
+iO+buF46Z2y4tkJLpTHjTEHKEZ3jhqsYWfLaUTIaH5YhZHnM/LjHgZWKNqyXTfwgeTooKVuuVdC
/TZVdft+gSXBqAQi8JyBItwY5fTvCjkZHtXV9Lg5Vnk9vmklpKZT+wCMc/Hn99BRuYL5xy424+7Y
+syl9AnCLCY9k1qra08prF6L/MXo6+BIyXHuRV36M6gF41zmNkSRMDryVhswuaryqzVEJW30zdgj
/Mjk1f/Dd9k+PSHk6iPKTQY2HUVfOEkgKsf/+GHATEZSljKMoyanftr48QvzLrh3lvd4nuxoTdqF
Tx6fq1c9L3F5gdmqRRfeWeO/ZiCZUHgVmmTAIsVLm1EC2c4efQtid+Rub2dA6v+0cwAxlFylU48U
I7kZOBoKfFklAoMKR6+048yQmqDGzMYGviQ3gMLzVOJk0G1T2GkUi14prAN7dYIDsuMIXS1x2zZP
sq039wxBo2zhCt7zqOVJv7LBICxuVcNRlhh0T2+Cj4UbTEveIDSyblR57uBIlhjpAkPua1Ap78hZ
N0dvQA9CLl0c9uZWi/zecW8boOl/NQdy4QS8uhgbAqckED+haoJthSYGabGlD2vEKDlztYI877gt
+XPSbPd9bRgsZtOf1lzgduTPPd3UUpN1h1aLC72mHKUho2JdNzd3tYy5GI9jOd25SNTxJ0zja23+
Dzwgk2FPp3Nn0yaOzU9DN+AONZ/4mRTrx+FkZto0FfvhyDBcZPOqVSJpd8bpeHc64rEDpiogees3
IkCh+wG853PXqV3eoQvePgnipORe+sfzTfhG9hQYD5BCWBety0tOY6hw995ElkTgrH1cuY/XKdul
uav3gMkRsKXRf4ASlA18QYatD8pNvybbt2pyLSGfX+lDp6qpo9st8+NQcy2YgX5s5z+nWUtQyGgu
qhNa+f9C7ZzBNgAhcJ+mhondpe2vbXW32eaSkZa0BlMUbTlLo2cePo7tMQxIeCyIPXlAm5IsEvc2
spEY/LLcEPgYgcuKrNSqpvavhEd3FtJGTKQ5qL/c+tn+rFfkvQ5RQpY+SGaAlQtOET0HaoTuw8Iz
QctMVH8bB/2NstlhiJ4VrpUg/tHghuzEXomvgj8BfgQYqEXMqx5VNg5D7RFayO9eoyku0NTROijH
crFlxsHHQNvaZXhOj7JtPuHZNS1/1cRClAHHa5QdlAdqPgCs73gA8ZZeIDk9jDkLq1csdZPLf06y
KBHKlQk/UdWXGO9SENCRvL25QGkkTXfibNyRGZuuALSFKiq1sy9wpvlsjTmKbtVXf0M2Y79M2WR1
14X/PHuzTb5cPiuMtBdN4p1//HGy/IBEjR72pOgdzW3jjgUizQ2yZ+ZRA4YBaYRlzb5nXV1MxJmX
puW7FGmoRKxe2OfrwyaHo+qP+5/UHY5uVoZKStpombliZp5Jbq+tp24eAM2cvNfbgyA8RtnGfkI7
drN/iMZ/j+TTEfbKMr+abLIeX4yZpx00xleVmD/mQV5WTdn49ULT/aZLx1DLE9hVCy/YoPsHjead
eeLvkZswJ02ObTlttTejQX0UJ1MU3ah0g/I0l3RBH0jcTdUhuM16WtT6zOUannvnVCSUC44os+YO
86KJ/P4f0QPnYcwOApKAJDPpnhjXDNN+MWkRMFsqEKqpCjpXqmnkfWzCzU2iApxyI58zvuWJo7Yi
x4a2PFi9MEHRp0sI2DWS4V+NQgMfh6RisFy31atnzE1B+y6KJ05ZBvmutpn/sZEhPuK9ssvh5+TL
oqbjtEsBMavNB5DZyTmYWNFmu2WTjngnPTr5DYoeX6wH2YP8Hq/+qI6irgtCnMdT07kV5d1RUCiE
yhWbib45Y4E5Pi7QKhR6E+EsJ7E25H/SV5LoNKAl8esBCKGMYklKiboUhR1YE19gP2AkLGX120y9
GSIO1EN0C3iefvc2w3qIjO0Wp6XdSa/NV2inZVtY2jnl8GNGNJIcYGqTgqdEhl5AqEnEk3aajh+l
gtxQltR8kKS04zjqN7Im+KwHRnd5vDrQG/6cLnQ3vhsPEsVRgTpUq/eEr0jRcF7jS6cQ2WUw/kFv
WyMEFOpzzNkYMc+/o+NatS69yLHWEb/ClXGNfGE8F8x2fZ0yrwr2kL2NkvYvDsClo82++6TsGbcT
2pOfs4uun1Z7FAuo/jBziv+qc2GyKH9MbcDiOIcZUmXU9mwnXUKJI9n0PNuli0OX5QeHIugSQ4Fd
sWIGvgl4FoZrilJGTu8DxBheLHd2dIjpcVEa4bzdc0FqNUaGuxM46TaWHwpoMwdgLLphwva/6rNQ
S87y7qBrSWkpmZqBMRk6n6g5REjEmscytXEM6JneiCT8HS0wMY5paZtyeh2T3HwrEbG5P50IDJOk
QdIpunUr01aUzVHuhIzUod0unmtolTnNl1e5ulylg2+jS4jpshmJr8vAUHc9/KN7R5yR8MjZkJfi
9CW+h9+GDfd+84tFQG93LwIwupELNmDY2DCbWJINKXnu1P1wOrD0AKbdGXlg4lH1s4NtfjPZiD9O
OCZIQJ6KaekrIyUwH4DhyRSqqYABK4ITiqWYEXOzNwOPGN2wdOcm5khpatnZi8AXvrzN6S2nyrhw
0nxbWRF19uVr/dZdt+YDaIyyLnju352fwf20kWFWxENKUFKHM+R8t55g4ihaS4DftqsyaWsBTND8
cvHWKEDBZqaqTG8lLynyALA6j03daBFB8g+NM6lG7LEKIxrMucyHcgd2+qw+w2NlysGn1SVwP0Pc
CTeuHSAuUKhIAdwvvTyz/eKKewgqEz/d8x3d642q9uvhprE8BDntjNmiZoRIdq7vY1UPpdvkcYg+
coXA/KbCMjD/bKxT0E6a0P9JC3KaULUbE/AlG2OII4BjmWvbs4UE5r7Ya8CjWgekYJqbbNM3Oqbu
+04hpVD/cofJxMocOfs8D5VflGicvJ5WM1JOYvxgxuhZCTBXAS2dK8eukqwCLzAzLa7bo4coRc9+
tyliVn/dGwVFBlBYTTjFWTcyciWxEm9z9SbUmHtmDR3VLqBVKFU1Ock9Yv2QdwvCZpzAZOTFHwX8
lnNBAY6xlc2X/uHP5XAJNBER2+Z2NPtn3cX4pb7MlWBL3Rq794+sucEekMLl0CkxVSqW2oQncq+w
GKLn3uBAjMCb0Z98tb3ns/8xhXds83AAq5lMoQIQJXGnqlDS70J19fLuu6lNX3dKVSs7F4LrZJ76
b/wj33li4WgblI0UeZ7RMm6yiaW/xNtIXAG8w+XqFzgm0CIcOLH6A8CWnGQQ42wdn52QnMAztPBH
SOwOLqZE4yUjlH/qzVQ7yzMCvtVgHX9jiFhMrK7o3MFngIR5MbCv+kzsU3vYpr0xiIzD3fCt5Sl1
QxoVe1t7WZyZ05+f1DtQDcSpJuaZSwLkx5rxJ7zzWzuVmjMN2hxD7J4Fdm41KJmW9PZhojL7u1yx
S6CYCA/tDbpl0Ki9bkgiRwAWPpD4v6QifnlPoLtU7KonqzaWOQpUofL9Y8U0Ti+7rOWvMIjKk3zA
Gvr7bwlR0xbgKuESR7Hng8UBKivvp6XjKkQpYMe78Fo//b3gO7r/E1WJUIlNGMg4bAyv3uxd7oid
byPmQ2gzI0o+oqINXrV/sMODNYms0EIVCQF85F/bOHKtztqht8jJ0iWx3o/SX7c0kDFEYo7eOmhh
TD5ZoVfmtT/dDTCroaD3cc6m8X/84pgLamsQexBMw7CFbcJrCBmnz8lxX9TRDC9JKtBOrsrHtfmi
TXerqbfQE4lKEjA8IriPCRU6ZnwHSIZoQyqmaybYalj0CheOl1EkHifynKy5qWo7BP51/7i4833u
hHKqTEGAVcdOI6KwRo4tj5WVI3ewjdf7hwXQN9u0uU11foBOFbsxvzUe1bUnPCuQ/Mb6DdkdIk9H
SI+tIYyaDrgWSeqBTV0s2RCwFchAJUXokRB0H06QON1gEKH+suIXvHzFPhSO2HhjQtT9sMMnrQT2
h7mlS1uDoK5DxE9BbAv40PbWvZXALcVw/1OWKVNo/xJoZUgps9pKbIBpdnUWli4byjEbKAA14wXr
ZN3+uj3iJFH/tvbq6fZwQvpCSU3CY5J5528d/i/2IkCuMKG3ay7uoJ1tn5Dl1S+8umvghR2armJd
nAaqRpHOspsBTvpP8j2PfbN5Xw1BDfbUex8fZ723WjfJHwVkNTYcljIQak5duxEGY3GrdjB9CRaQ
nyosbiH2z0uwbbUTtJozBL/c8jUR00M1eLafatTjTu9AGGMH98lDNwxEZCmMMBydGkaJQ7nVsLE/
eiMnXIWMECnewIxEbUTqLuaFY0gYWLT+jgcVYFrKwjZFBt0RWGtXdRi9jPWpSJcLIlsBZbitgDid
p+xukP2+UcuZ/MZLopBebvrn9Vv02XJFm6emyv8fPnt8g4QnyIuCwKCqDxHJOy8XRxBzm0b5iOd4
pn1Smvb0Fc7VBmhiF4+/rm9hu2vRmsRYrGEVeH7pL7S/MfzTUxQ4Xx2YfAgAymtHTrVJZmL83YMn
BzxmiMGFT3PXFs3d3yZmvl8llzZSylrzZ+TqzyK5AJjQrZog4SeSeFKA7zMLH2d3mPUVvk2Rb7ba
57ZmpVTB2GK9MzggloGjvOP7Kx/0EIB1ftFz/rWe8IdEV2vxqJS0zNqRrnglQbrSwCa7V2JPIri5
UiXqgY3jvakY2RVSP9rQzAc2ELHwKIHz6troDB8ATsaKfeL87ePX9nP1158M/SU9geBM4fdJZTEj
Mrh+XqCI0GAzFeLTa9XVusCrTjYBMWpRd7keeT73L3BY7ZGQbsy6WQnvFPQ1IegGlzkqribAzonm
+KhKlOlpSGEQKoAp19Rmt1HXXm7o7xSAJwYnq0sxWO3pbxzKpyH4v/Ea9/jOmqkv56PadhjcenNM
V18Hlt/nnlwqhAmqhsNWIefIAqgOPHJGwE8/+la/yr0zUMhC0ZJ5MMCwjZI93sZsDTtxVTObr4D6
/AKg/ECZn2hCmzKzJzZP2zQyylz0Pc7UVAujQDITPlgL9QsgaSHyyb8/IHgbcE3Rmne038MPboPR
TbPJv7M1pixdyt+ez1pz8pCcbrQ6ccJr0YUaIqkRgK0Uy8Ltv5aDPJTJHiJqnh+V0/WMVVvRoJ7w
g+xek2ZAVI30SpkvHVN7r6V9hrn6kwStetx5yfoEI1y7cp8GteGvrMVyEL232p54qKQncc010Zwq
lCVmhJZpyIRnSdLkaxI8F15Mrue5HlsTwhGPKYL+HpLPKrjd8jcZnYM+9Gl9XmXfWkjpxkaS+fdE
PuLzq8ymMNgsR560jXwL7WT2k4snJ9A5LEbOF3HAYTJW1JzqU2mxB8v984jRd6rK8iCPvy1qPGiZ
lYF+54ZuF3zOLNUcPIDsYAEWNeF34u66/d2F/hxH4g27hSMB2mPg3gKmsPsnxeDDmTXsdRzNa/ka
ZIkoymOwVuJJPfrOYrx1GoYb5GCecZFZnKC2yNizZv1s1ZjmJgxRMjg+M1FIz/NkRf2sKj0ukb22
0dMRGrQgvVLaGnhPWZuDy20Z9rBVrvx2/AcPFpXU1nee01M2Ce6zu8j/zNGq85Az4w4EPRJO9Ik3
SBIZ4A9AIj0ukf99DpaooMWiw0fU+AQE47Qh1dnJvIfUxph5Qh8VaAJFfOfmNvvTOHWCuFzkYJAw
p4k4QoVIbpChchXz14bXM0dF9dmZ1H6wAXiMWMCFtDjS7Y1L20htRTa3rmB0yUf2xXXhEbibcmHr
QgN+HDL8vWhvplh2eE133QwlmstLSilGUaAfN+xzgUjFR8cJNn5VKBl4aQHRZIMNRLakCDtb2OZH
gXp9geEZ9vKIdXW0qobgZ7Gk0hqZJGv8cqxlbgBRRbTvxFZ4UwNZVOzl9+l/3XKRtg3gvfv2QC/j
A+IdseShwMfx1bOUPnuujey6zXNYpViS8Awj5H9PgW3NqQ4qhuGuHZCExYkN5WIUwAQSCpEj8Bbj
iS6qAQrlb+pp9UNE/HUzOYpkjwinch5I7QSBTybtS+dmQHuXeprURRtHrL0EGPzH5mJFt1jkt6c3
lWqja23kFWzJXDsaC3bIQYaMb3npMAvBzMyXAJUX7e/POwpURCaVVucqcmNUNN1cP3N4CdLiwhBo
RLXiywM3yLfOR6MlRZI+zokmkXUGjQvzClj7DsYY/2EODKNhRiT1a6vQzqDbI/KNZsvBliuRfb9l
/8dKlQTpSL7kmTZWN3D0dSHsE9Fx9zhS+J+SEKFIx7lQHkSlkmqq9z98GnCdDcjEJBV7DuidhXIf
KKrFYRMqleJBav92Tr2pndITIlMIK7NOyXAssjtX0bPtOsna/zukf+jX1NZM2oHaXsnCPZy3j8ip
27HYpGShVLpZAGh3i2oAdR0Y52n2MeWpdvsUI+nTslqShuv04stMrjGjUX8gFErhq3QIXfIim0B0
6gektsEYgaPyPGGIwx6YiZVOdJ/Hs08Syocp1YUw9UF2Y0TtF+LMQxTlQkjtCtXFMWa/w5fmv2mK
5EnE0sjVWeBq8a61+2I2igknuudKSCCet+Xiq48S2L7sGBbUuR3+v45n6QwBhIN6v1IladxeqC19
beUADbBDlxx/jj63gOpD9HrIZdpzFETod2kQ78x7fHzpS3NAlnGHLLcUD9LXlKoAMR3aWHmirJ+R
nFlnUQ0jGzbdohdVMkGGpJQDYsC5fbzVW09EVwRRNQRnsFjnoNBF5badT4oAP1cU8zhf9/6ymbBr
rYl49cp6+JQEiTLAGiqhwkl7w4zB6J+hRLMcA0WF8bn0rnFjGFfWhU29AVZuUDjzszaGMu0wInfw
f10vsav0P9bbw7H6NCyogvJIQ72xA89p5CrP7h+s1qEj+AMS8weCfZdXYGA8FH53DoVIf5eAo2/p
tJxclYyG3S1lpNB0TPWbvOC4r2/aRKjhvdWIUm9kbCDD7MtEuLczqcjTLWrXowraZSo6i5keLkrc
PEVtHRTpLz/qt7jXQFacdCXXKYtJkAXGPGt6ri21cdxNx3UoM95TAxBFndBdKlwRNQ4KZw7fyIOj
pQpNKrVmc9BUzFylJZM2ljDEQ1TQLueLirooLitfplYH3AmuwfAHk1lCFd0H1JnJqZU/J/4oy08D
tG3M0YYOJ2jOJmOro4wWCt0rMqEwa3VKm/HpKKB2y4DcjR5sz3/rHV0xNzpxtJOABULIwtQcN4eS
dbxc+OR6VWNeSvorTLj1rH3LsmhUO0uJZbl9EaB+5LVaAPxF4fjylXOFj+G075yhu5Zu/+VyBj9y
wr3eJ5/wMFAfEu+eGmxJunKQlSi2kwy7/oRsHWmX2qKu3CAZCwNDsla/FgjEesIH7wuOOmLCJCF6
8/dE3tA4Nig0z3ykFlVA/xYm7AY+P1GJ3K/47ZpauGKxWVPbF/jFz1wjNRTqSV82D/l5hmYaMkdd
DvW8mkreGuQtkYTuKxcz9JQufctUGorrIyYBQvb97u9+y0xNuTQyVHe5xNWqefAe0qaD6LP1G2G8
fCOcE9OYZLWwB49UBO/Fww8I4T2vma0pSNkqJs5n6bo7pgqU9zWFS6nTwiJDRSI+VGsTiy1BhSpG
koR+R0OaZHUwP64+IxVvmQftiQerAKPK3kfGGSLnmk7zeiU96ZslTzWVZqg+0pMZtZCyplWs6Gn6
vjVfKRNvRDrfqtOM+qABAdzDhBLPz26/4fOA5y9KE90SOJiTJiBZ2oTFy2aST+yzf+TPx/Zty8+l
oq0lAEN9WjXYJ4Tr0yxwX1Bkf00a2JpK1TEELKj78Wf/kbbtbhNMhHfNTQaZXMPaWXdb2XYo3sTQ
WLzp7NKO6cpNsnQhCpVIn0Z/xuJvgGYN/cbT3g1oHOD7Pjg8fT3YXYX6mRv8LQ2xqFwcScg01WEG
Cg6Vc6uZFxZMjkZZA4xgYBXToiQaNIHGVIyPo9u1LUjm9Ds30JjgHRbDDkgHtFXWCgkxwQfHaeSp
/eRyn36D20vgcUUcQFdzZayXWe7AjOArEaqEdf1jwOYI8ZPTAQtwybCjjKjtvhApyW4OqwYdVfeI
Il2NqcyaYSRtqbFyXIm92/Upr4mkfbpG2wEv2saRr+67UDTRN2J69sIOOlsfKxET1kibni0VJqyy
N1IG16PExmFqolYZ8SLWTq1CytyYYKDe5UeYkgsV9mMqNlg8anW0uUUbhAFTaF+YTixVHf63eGWM
8c7IkRXMvczPqG2DJ03bCpQ7WfWaRYh/4zcJEyYY9WHuW5UtOIaFTb/kpLPk3Yox7zYgkDmdodno
MuvviAXX72sxiIkjPt75nnqJGjRn4JhqjqOkNf5eqXYjAqXg5cBFDewd+h1VLvJAkRy0cNHBzkpO
LKW6H0AibuTv1YZFau4X5ZflBd76QWNU+VnWetKENRnGCw1BE5cLGDBsG7onETi+3j6E6VajuG3Y
d1RAyDGT4Vj3BPtGjLLgBba//HXbq/Qp6Rryj/2O15hEC7rKy7Sg9Tk7p+qnb4CwfxDeyhRtnL0c
ncYlWwBtZBj9dplHkY1JL9CF7inUuPSpZHTS03OMa2lpZbwRzDzBwuBmhfw4x4ZAaTUFdSR8gFyR
rTtellanNJRRJiVZc6OwcMRSK1YJl5l5tx4LI+eaGTUwRumQ+ASKjO8zfCenQNagoqpFFCs8whh6
LTiriM0Laid6O3NwMXwyV1zTMvY0L7x17jgBPsPJF0p62WpP8GwaYLnM18Rx8H8hYJ2D0mv/WP9j
OV00y7VvRGW/aNvnVEJ5xDkquAp4jKMyogrPfpKyXQVFHmibvOx8kbMRLXiNRC2vzdUgYbDaeUFB
obJ6UO7HBCPUpkHyYfyTs60x5Tb58zy1ACjXecAYZU3XSfp0E6uiSmw7DGvZ6iwc6bvtf221CHtr
z47OT2ub+gLjpfE5Qv9zoImQAb+7QxAw3WT7l+2nYy5sspaDkEhLuG3oKFIFlseM0V+ERUCmC7/J
FMzRoWLmQ4sqFPENSf7VUEROpyoL5cULLEPv+IMnU/+W7AmiPvIQobbJ+xN5ZvH2MNmvg0w+rL5P
XzEaNUKIpY5QhjCGB4lUkx/0u7hcd4oHgVo8IFRbiLjDjPsAQN6PGXdiw5t8s6Exe4+xceZh4AaM
LSy3gDHGH3hbAeTJiLHzXuOy7HIxpncY7MjlSOxIpud/5JGUGIvzwO3VulRU4CS6tWOi3HXLwgnb
k4+EQLpwZOvvwZjyNgyzj/+mcIh51SGtUdjUBP+rFXVRsQ/6CMmUmKV9rMvoGrsNCtZdp8h4pt/R
jKeLBDBdIi3os9kS3PdlE6UNREMe2Bn5ieEIsEMpmA3iYjUYIP8DL423l+2WB5onIzJt9P8T5jcx
YCiBiCMp+X+gHGA0dx6eBW8R9FLshniTwXziSjCFFqDQWbK2wKORTClKleqmGAcBAH7lK+f3zVPo
rjKMPzae/ugy3KgCycre7tLEjho9zmlB2fl8jPNXcdGDluK+rIkZfmDKPCSMn6pn8MoAD5Odb8pP
4niwg27Xj6inz5/bni4np1MuXBbiIbVZq6effh8oZmEXa563F08DOBennM28hy1B8ui3YdAtnQvN
h1dBDLVhVGcP4R+QqKH03SPagGvMhcdLzpeNNmDbLGCu8xym/RaZ2YEzbFBn/adtRjsqTTBhCcQS
buMl7jQpGddfXZ64f0Q/cigPxvrYBFmLgTXNbs1ayE4AoqtqjW6kR6hE8N1g77UfVW9TJMNSwmIY
YA79/lzyRLrNHBvUQZSHSCcHPZORJKyyxhZFgN3PoytzVEqYEBzN7eKW/T409KHy2WNTudo4VaSL
5JHAB02o5te/3oSpU9a5lJrycT0rt9Fd8VJzpY/P5JEXPbmw9j02EmWxGND86ASDtf/h96VuHMfk
UjxTOzI2gJAVlMsrvb4Cxx/KXzrVEtRNze2c49iE4o7k7m9wF/ycvKbQMpc2J8bnbwN+IJNf78Us
bsA0H+4BfZymvp0RVohhwPg6K6fm74MFwt1C39PBPhSL0xglTKRTrZQNjmsKxCO7yyK5no1EJgz2
0C3GSj41tkR6jk/IhkPzShgKJOjR2C32amxl+wbG/i9XRgK1kzjEQPP3M7c0Jd2RamqdQ+raWokr
GpRcJWQBym558Z95Ub4oH1AYoryNY7tQ/X0TItynRWej8mXFqfp55Ulwkd9zGzQWsMGK/9jTbJ8P
QJn9quT6w2H9Xs0VBw8Pq3B+6CYgKni8Va6vFjRH3bJwWL5mWOlThg8iwPvB9bAXGHyTHw63gqDX
Zuhv7l1My8JFitdpfi/yMbgBM31VVpZz4frpdgsW2M7eELVZgwjzBBNxP8wXMUQbyoyXMKPjuSzw
EgB18vI+eIeY5JxOSgNZKFiTlIxhdxytsprssfViGZFQIId5qOwDn3YjGQydWSmzmKSOHCbKtr28
pO5Sc9NdrumGVYZFtroK+euwE6+lALFuAqrL2dMhoWqJycZq0StEk9uEFT5vATk811Znrv/IPZxp
wui8cdLq1WioFKiANILTorI7ir9ISmHicRznVYJUkOuhMpUFOvbqWPlDb/5aKklFgtf/xPvkHTc+
Ymlj94CsM2ApgNJPm/44OVMuJdk3nHEmYjNx13ozYGLgIBoZKpWFX/CrH3xAHj3TtbsAABMRkT+Q
clHuh+CTmrHI1KFwrD2si1toGku7HdW1flV0VfpmpKAqMFu9z0+eZZLQ4UP6IG4V4lI6R2b9oal/
hDBGhDMmWbQRHyp0D/Ltqvxp/pLYPdkr+n05GbBTOzcuZ1qpPgMueSWWNpLS4vitW+S9Tec8OgJC
vXaqVjKUPBGf/FNifzTb7VEC41u6c5FyJAzDuzSYMy9Bo9JRdcSuzlFLMTVjajn6VaNiFv7Mnu94
FgAsgjtWgqRecfpLcgMvhuFpN1XhW47Fqb+e4zNgIIWYzbFDw8lAm8xoTr6voOWitVI7npG2DFDl
Rq3qg/DIFIQE1kAupyIVZg6vGxk+ypDvYwqgvPId019TAf79SIm6DNw52hisQ4x8efj50Ibp0zY8
OuWzkmYqehSHbbipDWoqZEak8JLZDqVz2nx0vcd1UcgDSy0YYFYJxWYLxq78FNMY2t3Tjv3eCfH/
gDX5Dxbtu2ey095eDEVgawgzvg0QQsrhoYR6NvDUOrqrrAv2ou4AG83mchvSKZRXXb9RM3ayEISV
SD96G8LKqNuRC47ahpd6+wlQfFNnY+BDCr3OeS7o9SHZ1Y/Dd8hSp8Ad0znxNzJfw5JrqyCz/gs8
e6J1fqRaRKQ/p9wvqq3lYK3S34pkenF3luJSm6/y0xM73GohM4zsJzaCNBfUcFOBe2O8qJAFiEWp
u1HGL3Zi69Ca8Gn9U+32yOetrNzQYNcxkPD+kN7Wi6pWYZJnH5g4Pwp7vQXGcxJKX9ZcEpj73ZB1
cKyL/MjDCHNzBKdp7iLfYyS/EyEBiX1oNmvF4O2CTWKRJQ+B37OftwQP0C1sqSAPzXadrQaw4IdB
IFUf1rvi+7ZzhP/payuyDWsEd4b0C0+Z/63SLQgJd4STx9jgYzs2bLj+SSZ7ztOxR1S1KGRB1yTH
a8ADIPh4OktKzHQbVKxHZmNZSzhPgGhX8e6cBz/vWhb7hm4l4OsduKQ5BzS1LDw/FXCK2ZVyOl9w
3iQsuJbrzR7bM97zZ59A7PtxpJM04DH4Fd3a6/phTpRlqjDBDA8ds9Q8rtgQvS32DkI70gNG90my
/T+7LDJ7kx98NOz7tOjt5ReJ3aUoT1XqpJJDaFGuk0lIu9yAA1pDW/tTduPBUh9xvpyw9w6IV8Ve
olh3cgBgeQuylmcEvkS3r44ly73Aq9MMbxqLBb320RDNcKxk9rOJV+phzmjcSnxUBQbf5QPnYC+U
PT5tTZ6Uili/lXI7xSpfBOU1cZZAvwshY+Cw2WhAZlU6YfU0KdZgbML/uAlvFTgt87sQzoz2Qg2S
GAWu52Cppqs8OyDC2RnHYogu+hfK35Szwa6j5XuMHaEISQThqm0v4R6V5WPmgQgZUvXatPeAzlzp
1GxCjM/FNmsTTOWs4RdDXKijF1iXvAvGawYsDFTHntp8JUHDHrPAKsMeUc9JksxL7xrMK7Kpf0OQ
PHCEUImS9LhAyIWAf7yoh2l3c9AsxScd7a7XNv3+dIZwZD/6eI+HJ56gbizpPSK+zPXvLl3OnbbP
k4e17u0HntslLqGNu3ypGh8zpibzv2Cbaub28XzlN/QoVTovFdpQamqgVNCNyisl0aZvvV3GwowU
dwndzFSJikSiuUJwBzoMXnU7DyOGePEJriO8LGYK33MtnmXrpy7PMT7Ld6iS23gq3Q2stO8y0Jvp
BQ8SCv1i45GlWApmPhYZq9D7SLcSHSVLKcfJNrRTJSIrCcqDn3m3kCx6ajmsOO2pJL3UOQPYF1rL
hyZCoBAaHfQ/jwpMSTve/8Lm/dlzrtSN+x5DxRhVdBZ9qNk4vhQ4WJksG3wwiz/1hy3az6+moPVO
CrCCYpRhAK6NWTa+YxDM6jbuMkRg5ge/VOuJ9V+Thyzcssjm9MZokRiDonQCqktyIUiB8AlPmRgh
3sEeXEn42hBWMnGDxxUKG8wCGAli7v8e+1KNWq5zjkXsV9CdnfZXwLo2aNBcF2ljtQdhsBjmLIUk
AOxvml4LasQt+rkUEWLMOZAtAitI5XYEFM+Ks9hdKfLPhR31AgTVbgb1FCl6gDguZoFT5iT5qlCV
otaNPTj5ZMT8SQVKBMME2boVLrvh8IlI2/K8jCbBeWWXiomkk53f5rveGG3dVYLjr3YYNjwgDuBC
nF1Qe19zQIvNAeOpxyqimtp08c6oYBWBmbxoL3Zsgt1eF7vAYkFvN7LomcewOqZD0SOtuLn/r7ds
NYJ7y81qNC1KrNhNMn7/g65z60JO2SkyKnI4JTvNs0i6iIYoRSihbbPUfSNVSiD+CUpdG/XPwhCH
6tsmXqgYft2pWx8GPJRRffyWLi4+3LBqqpLz3eGVnkvXuPubZQ4Uv5xSpwkrwDh94I23yhwS1PcN
7BUuJNzFo4eICCa85Zj143/oeggX/xjwIlzD0ovYWyUTLN3A2pFo8Ls8oPeNXiXwnH/kaTvLCbEw
ryZlnGmbx6HbnnIANeZWMNHM4H/GPO8S4Uo1iEHpFZh7Pl0jL8CUIZqIlwkfGAxuS7e91VWHyoaF
JNsmmw1jwM1m3FMQMGDllvkQXu55mudL6wVSKopsvyAMbEh8yf7ZGZU6P8CUT+C1+fdxWB9mi8+P
08oyEyGWcXLwcLyP0kLR1QbhvQfP09tk36g8hYQbKWDkaWCLzwwbiqa06xV5J0Um/xg7cBgqP/af
8dlTAdtmX84hjGbub9qxOeA83RjanUFgbPvXNEde6tXmRq/Kukd0Zcjo3GDUorF+nQMER1XrYe3t
M2nfbd57nFhSFtGNy6dOy3e9459WSifhP9YPhvHYv28KLYGTdAxCAoO7Nm5+9RP5mpTkrzyJuDlH
7ZLY0rejYLVkPrx/YNQ+qWzCuOIcvc4Qvvkn4Y7vrCOgbiZNMQWXc+t9BlZ1F18fb6uaeXykFc4E
Q6sTLv89tMC5MsEMmYwZ4GXBQFW3IzhezOWgqYUExgXE2lrAsoXjkm19kLtKO/QvdfUZI/KKLwgF
2ui6oIGhkng8OZp1/xCUrhq5qHGk+yb+FTcMg6++WNMm9WwxpoF9oQpDH87LufXaHDaLeKMzkA/I
a4V2JXQHDg8eH744CrgKrgPE4GmzA3t5Bz92pINDB6m7bttRswUiMrqVUkFn6vnzN5nd1szIam4e
cpJxZMf4bGUubMbHiGlMG0fGqWREipGim/sHxg08b7itHf/daOv6+BEvN5rCXmDhGBRKey7HtNfM
fS/6oriCcxnJO3vo6GewYxsK01cIxnMwLZv/h3x4sIGSCOSYGfeqJdX2HzqRgivdaCkcl1EYhDZN
Ew1wjdlxfiMYCNiQcpa/euVncFcASqCh8dFS9o8S1LGq7WyPnVzmyUuJML/xowTKKqHSEjsHNyy0
U2V3SZN9wSeHMxAIwBy2mJeoE47b9e5Vi2fYxMdPtlQzO50MOKFko6/sl6b3ZWyYXUbqmcWIRHbv
TKDViMIsyrgdA3/UdOgwx5v9ZyUsMXEabuxrja1zLrOmDjDkq5N1+jzL4xuhHXIS4RzFNuC9ZymT
BOJTN3SvZz3X0vgKdsAqeCBes7Z1iN0ZExtmgwRQgUjEnxiOXXC1Wm1KXZXavOSXEnsiNqdubHm+
QCad0lt/PEqNRn2B3GS5geOj1YRze1RsArFNpopl1/7uXy4z1+F+viGTAdXOsP3hrGL4EpHomOFd
wIAdTp1nPTbtKGzBE/65sZS4yudkXxObTX6zDdbLAGhH25fIIuvjxMGANNKv+Xn+46a/35hd88Xy
hPs6EOc6LYySpKyJnfTcfNUyu1P60bh6YGJq/YqQfrrADSviL3V6VtHHMVImOWql6/heqanNX8Dp
DMUfz+Dog59lOH8q0fY2Zel32y293G+2m3govVtopKFLWM2XGrCNz3nfKWa1XQ88qOEcl20OvuwL
qFdKAizDJivK1EYFH1CRNfi6OKiEcbbpxVaNr/UyQ9dSRXO66ra9PlAO5bYdcHU5Fra2G0kNTK1i
IVzvPlbCvsERhhgxSuoejVX0pR6TKFZ/dF53BiYDFyPn2WD686zgz+aUzb3oEJZ36nsjy11ATtky
6P719xVufhbPm9vWC5SX6vmdr/HFT8zR0SgnbtAo2OTxnaHyabtYlk9NGiAZ2sBC9rpUng0GB5PU
CWaUb1nDpRtrgKyZsMWqT233bn7WvYVXWa9BUMEP4uw48uPrhqIFOZArfGMyCA/50HoSAazIPkBm
arHdEKEQqei+QzwRWA3XDkahUneH6MP7d01F/FITUe7wlwboRoj+hjgdp2gUQ+Hxu1yVbHh2ATTy
sNmYK0KzuRSeliUnhceRpEYU76sMtXstsG1UBeWWMqlXxOxiso8zaphW9i3yPKxE0IYptqo7Fuf+
MFJhQJR0F+99Nt8JQmVy5+MfrQxNXaVtYdWM4m/++Cbi3wtKrs31LCTUv93iz7cWGN863RzjKFp+
xAI2K2FQA2y3IEEk4r+5Q9hGdDoT0KP/5B1OKqcnpQSFw27zP7ujp5xtQ6C0XgPZ8VtEriZMMT5W
I44sVDW+iKCvrQLSieA3v513QeB5S7GGbuNpAM+dtugmx/+kxHKRAFFpM7tWCGgZS8ICU1a/60ri
tX3wIBywJWl4kjx7K4+JAiHG+tDlZ0Df9H31gmVTULxvq9+xwzV7LAb0imdLbV6s8j9nMppXPiv2
ehMG0EGH0vBq4GhkGVMMiqonFF+aKMbf2ZLKr1pYRP+cpKU0MSJYgsQ1DEybgFBRypR6vu4CnFvV
FhIm/GT8KZobuELtsLi1mS9PI2kB1Wyo9up6J66bHX2a7eXf7FE9gWvGPoR70mz280IYsFUfHmZE
g4qIxveC5qHNcuw9XHel6I1W+gsnlU+qtsCATpYKv/HO25kw0akFOEYYouEPp5FqkBV+/W5ldz9F
s2CgnX7wGuz67L3Vj8U2j/aDHkm3WQaX8MnkVBb8wf5EgHydIeeQfFHyYA35eDcdSK8JHU6O+GRe
aaLqWM+0UuTPYa4PdGXSHDCxFBLCDmrKuHQAf/mtMwGjZfpi4t82s9VVIOMiFBwL5X5qkwhm3h6k
mLjXD+sWzRsNGpSySFrVQDTJpguWHOnL5fW7Ee1SijDwJbOOO+Un+s+7mHkAnuxoDeXxV9DR1HfG
d1IAoAd6GSbmU8dnfaIV7eUJ9LBCTEUvykYkTqlpZRCwXBbmMwYnZejWAWl2XFfE5E9DAw1YAG2B
lK5RJl8EPcCUpOTTqBLktp0w9opMCLwxklx/okMggBkoY8DFMRSqFtUyKVyeK8WHJ7cCskaP9U+W
I0oB3Tsl6FBuc213ua6TcCJ7kAlGvI28ZFGTnqdiqPObcJDXTta2fQUBIGwggZRduoU1yfh6/IoJ
mFzYQEPp6mNYVfuZ08ZuxYETOKJSB9E4VqNKJqDwzImrbSQ9HK1odQeuS79QTTwi1SIHNLM0/otf
lg4l0cEGIJLWLJ2SlnqOKlIgk27syL2hAN5Vo4YL940c9yOtVFR0lHs1tYkEVI8t5xw1e0qX0UFr
Du5+2KpM78PyTOqum7zyfKP6+D1bBJl1EKRbreRzoVoSnip6GZsdcV/no+JP+XnbKHln8NitnLXH
G53Vc4FL8imGlLwxrzk/8eLjgt2xDpZzqtannNG7eA0v6UxPbFmrhjDa8xuDar24awOhUPKRrz3s
+LTR8NhhNakt+YETIq6qXJgIsYC0HMl29P9YJEz2v+UGpt+UCDe6nC5jXPQE67RFGp0sqjCd8Qku
YGgwq55maLS4JD7STPc6jvXXabx32u1tW9RWRWz8Gi+eNFqTlxkHV1fUW4zsQJ4dvNfTtDFP45P8
bCdhv7OVldudpgNj3b7cDJkt47WalYpK6RrhX+eUgplLVJwvUPOKnmMrO3Mf8UHoLrCvB51O1nw+
B0S18S42i1liziYAunAz01QmTf1se4nwVkQtY/jkV0exFYUr+mRUFcKK6Bw713RdYrKIt6LK0KKk
7aDA64aZFApACGaMvX5/uXGZsWK9OQBGdIDjJV/amFM1hpZbjq6LQ0jXVy3Uwmzi0UOYs9FaoOAp
HNgryZxrMRz5+/1B2Pkva1V3lCPb6zf7TLH3CNsKLg40SgS3XUnD12lMEVrFuCLf2pixXUoMRsMa
4Dlu+mAdvRSlsHCRfr7Hmksgx65Xb3BrDK6jkAjzplgsJkz7vQYlyYeSbETNMvTlHEIgaV++lxFp
Hc5pDNqo7qmMrH1Ej4txLZ69tkmFoiHxQpwKONL/QBGr9ZKgL3GuzgkrWjzhiLMAxTMEUG8zNwc7
9I3f+mAHzis5Lvf7Y0ZMFbqE83nZLE9JTG1M9fjbRns6TlHQLtgSBalou6rz7OtHLy2nzhGdQj2j
jn9XMTpnYFtt8YvuX1Ahg74A/ovdRYfdpjxzh7awKHPv0FD1G/yvA7xOgfxu9UfDUEU8klBjUNWC
opp0XzvXzMjeqJf99LvAMrRTQLr3fltm2rQtAOJS6djlfJqml6keXQoAFiY3ZXTkDPOb/sS0xVrv
yEpI3CWJ5M9C5bTviSrvmAYmYri8/sIM7xCSLXb59V02MnMFpfeseh4iRppOmJHZe9SG1kB+oa/A
54LDjQLLEpcG827efRC5JLg4gq5kt/VXktbnWiTotqyMtyU/dhmy99eiRIkduu45vGA6ugqakDZb
2HGDXml/382frBI6vl8SGx7Qv3NQQluF99HgJYp+aBe5B/qeb8Qx1z/hJf2FARxM1EfZiAkQ3J4U
x4wN2sidYmAFDmZNu8DcEPatSV/Dq0W08BSKCtyuLlE0RxY03c/AKhGGhWmyEq46U0KZrVFR429t
Dse48WxEGPqfgQZfpHOd8qR6w4Ts3K1u2+hScUG/dlxiosgX5Qx+8tBN+OqtgcxJyQylwKCLXTHn
y0PalKD/HedN9ZB0WbD5358uNZwPAVuWGko40VDF04UzzxoruYBWaTUcfHwgWf7kC2p6zLc8dJ4m
jQHrSF5l3ibiWakikCiqWNKHtOIeQdAjHwVv7Ra/Z0GWnCcTD4QO8SQCByYZmzALPc6LfZc/Xj/h
TDnobUv7PoZOeciGbyLMSkQNDZGE1g0byOZ+jUtk1tK1xecyZNbQtthsXVQHrQTsc3F+Qwg6ClIe
Cuvac2nMgODh1Wenrdi0fJpfnACMe45MJSS4ScXIDKoubGzz2oj0ZjNkETFSQqBSrvEGCsHn8tBl
SI2rHelR7cen5sir7S5L+MA5QfOQM8vaBFbj39l+8Q79ir964/0PpbscV2LZr/u1OiM08UnD91V+
4Sz3DQrkCs6rxizwN66WvIWm3ey0rzMlPMlmMpvpuMLscazK2TVW6btBBuuILr51wxMwmqrXEY7h
qMW3QcN2n3qisUux7SqkQGHSVUmaonhihOqMKhjRcnmdwNwDgqeGe8GwXa1hmM09+aUYDxnnkywr
+Gx7jvMG6ti7QhSkDQAKpfsdLRnkNNBMD58cFWMHmWdx1UAuG1N/E6pTpqS0fuZfNvg67u3yc5ki
zJp+U2UmZdlxb4s2zogg1/FRYHmiLEqPoChY+jJwv4TZ1udyYDVixYyMQbeepsNbFf3b2LI8C+hw
+okEQ2Lltbxl85Vd5JZKWbPJvO2OX4hwFdWfJtGqa12Lr3LTzydfANl53aJ3gSmoj8Tf+Bf/P8FM
Jez5Emi0I9Cu8jrm4iq+wSMUiKD8AVFvQKEfHpsPJYjHdly7DpqCzKtjr83W3eQqDk1QomPtc8VV
zawm93f+dG6cTAsjyNFFdPnJ9bDsPgMHRu2bEN6/vLYViMz18CWkqrB+EYk8uOkJEicbPyiZ5uQM
QH2Kcf1neINOrlPrTutFaJOserujhGjhpgeapo8oskWGx7BwngpsuvurteZ1iKUQOJV+GNZGtdeR
Ur73MEOYs/U+QiEuBR0F4+Yo0Q9RG/RY54k+YHW3S0aU/xvA1tTpfp59LDZtQEgXnu2FURwZYPli
Arc1EL4UPW3I4VLuq9+xrg31UWKayIrKzQ5GVAi7LZ71hg7btz0XFDfrElCdOhfDEcwjFvwtCUM8
SZG9VjS1KwQi7T3DwPhE3NDsWzzEWE6UNAAyDOsG+4G0+Qxp9EZ9FcnyHKDpJJmU7/7vn2vz3+j5
u29k386rf8X6qMoiXwx9hiLHaZ1QaAg7Slx1DZYrxowv69Ix69prkSnCjMoZgCnFS6jJsPxVZIKU
SFzqULZozdyG5tR8gmahUFYgfdy43mLHweGb8XNvd2c/FcdaHU0bZjld023KeDusRl3Sqx666yfl
PqAGqBHJPXayAcykAQAf5BJ2PD8XPukmoDfLwC/sl/f5QcxpeOd9TVZrDbX62VQmKy+L+J0GNFg3
/JsCs4sVti4mr8Zg7CuwYscPhV+ef8TP0YJgeTiec3eElYq5t8PCJIWzzEGZ5Y8R7wDb8eZMqmkS
aWMRs+nDLb0OA2GYC5VzGllKVFNw5epVvaReiFLfNmiJ5MliVYcaT3h+FwktY9hEwfXTSTLJY+Kv
VhYqvBpXzKDAWz5a2N1hW4+Qs4yliRSkZM3gCQn5F8D6filsOorGWeL2ws2UDwd7AHm8pZ62BpXi
6s7l2VAId0JqQemkvmbQV2ckUPUnh0yahJc0lTlB/Q445+ixS2FEkAS9XTtxE4ZT4qLgRE6NIJJh
upG98diYC7TDoceBTfplf+5tCoSXpyXu2Wz0+vLG1iQ7zrBURsPDaOnNCPB7Ee5gBF1VfJY33ur2
d7AlIsZwzfBiDBA/JVHAew9Lp7U+L+IsKfZjE/yNjeeDyv8RL6Ax2n8C3L5AGYDPBnousy5sGzIa
wMT4M+PoF/nWl1Kd6aPzaAgXBD7UEaRO5Us2Rx1iqe+WdSMbZITSh0BbStKTXCv/MJi9zRVJw0Ro
oh7NwNFIGr/HEOrhUQMAJ2Ml+alxU+UN5DAcJ+WvHoPOfh/woMqNxeqp6smAQHoMTSRKtEatGXhp
hPO/lLDkf+gvVPG9gvcKUGEMYrrsyHk986mjMx7ur0Cnh+33qd+rGzjuq8swaCvOu0RnFiVmToHt
YB8oNIDZTxpeskf8EE2ByjEqgJoxkkTMOMUCdJX0MyeeAfUYVm3OjNyXvwPYUiCjGB0xPotrZa5C
SAyLy7ZvzaohkR6REeSLARG/rfpXObyaOzK5rQJVPZ8zbtQnUqPrAHb/m+u7gCCLBoY7KA7iICUn
qZJTNm62j0CjWsGDqfGeM4JIoHaYlGXHNznu1Ns/ywmMIaJMH2G4oulBH7k/s6tbPHF/8lQa/nVs
dDuyB6sOs4uxRNuU2V9thC/c1igAZJoSv/zWIfq2kWFTgjbZPe60iLnhzA3CyB9yFjFafw0C5yif
6pX/oUmUyW3CLs7N5N8TiQz6pqmHaZL4cK8I3TGq6V6IQ8jaKvR2ERK3dms255RGUG/mPuGfPZvk
Ow+sQR6qT//nOeXt2AVf7cvDimGbIAsyuVRtKzHBaEtVRX9rRns5+zJ4VuEd9Tq6ppWYEITD3Fbv
51agvdVPSCm3zlXZ1YJurzosc2UyDs7WkxwGjGyyW5U6X51+mTz8HVqEoDmIUdHDbQtm3Ybonow/
kY34VvZLa/4cxG+hdmeV/K7duJCF4WellU9NIsd2Nq3euAgOTdnDItUsnVxV6+wd1hZ0Ul1/I5bh
NILUL7QKlZdkvzXtql1ddsI1czTWYRh697sLd7GYmON4NavAo2yrB3wLucvaBEsnx5XOMJ1xKgVO
3tUxK5hSk75SZZZvmjfLLp6jcBk4VUInpqLyQM9vZX/N8K9CP7RApTknXEQEygkeAlbbidwjrYFu
fBmMlHr5ELzv4UudzEZ7J1DxooAbyWgKJ3zXeX5b3/ssUy0RlV80cq4a3L43hR1Cs3nET6Bbzpvu
xbty/4oopLQPU81it+JDgOAQ+DidhPSh33J43khkuE0c/By6zCyz/5XYILSN7i4KOH+cyEhceitJ
mTGVpup1Ha0ym8coyLGb8+uf6AktnKmSk6kt7v4OcKe4IV/R3Xqal5F/3iItJoNj3ZtAO6HBM4D8
hh7RGxGzEPx6gYog0zRB3mb6NzRQo85v/FmVKxxswWuZtWL9Ko3f9PFnjNk37SzpnqEM7U7AsyBj
ikaDRHZBlkqY0mJAOJFmGkW2NKvLP1nZyMaTYVKNvk/px3KLu+tTkOWwj3Er5Q+QYTrqE0zFvfDG
3nRdv7zqRTIQCy+9M2/uWdFmj1vkr1cJEVHkGFXKrDZnDCH8uYLu8bUrMPsp7OOH9tsEsw73L9FN
1NrSTiWVoT34O5Dy42zHUx1oBdTedOdbyH9nyusMkwWlsdnJlyUVaCQkkSgcIj80XjtEYmAsRzsO
awysejxRZ4bgUhC2sB2vVjksWhgrzi6BnmWTi2AN/7cxbYGc9w/C14JVh1m8YOZwjZFzZHf6KZZB
+u0KqGH5SQGehHuOZX9YpEuooH61UkSLYu3CyzhqNDdfua2OBWzocHhaHHtO0iWfZjsUugoSM8n5
1pj/iyd2ofLciuhueXiXhERWFCIyVCRYEUTJusPrzxPlJK6MoEMKpRPQOF1oe7p7t+GEWH0c+koi
jkqJqKTZDjQvgL53lrrdV9sgSOVMcTj34ElG/L7sLO5Tu33epDCIR+583wUtWyJHFEipZMrR60pB
Q7vi2imZRS1QS+4p+XMl7tDwzEvHdYMphlu2ecGAAkMJqXBrGVh9FrOW4TZkf3rvVruEi+Br0oYD
UedTzMEyXRvxoKlESjlntCkNdvXI7Vfj9i6DHWUp2r1+9auDZosCZ3DEdm/mzpNjyALFLpuqd65c
69ZoQX3wwTggN1qjAvj4PWE1dsfRYGuDKzqYJ42Zjjr/xD++PHAVxFj9eCJLjNLA8zq/hUnh07is
YBzwI9gA0v8eFv7OGPC9rKIvjoR+C0K8Jiu7uiCaRx5fqQYTJOqnAEnf84b1N0cDyKdggxrmIq3e
QRSMbZ1Uiu03iPz7lvkIr6PAx9qJDJTdn3QL0Q7UTJiqfMPi56EhQ1GFSlyANljLKPq26Ctrt2+8
t/kdef6HznaL0qJ8mVnThVAY/KzeesdgUbDho8Vt3DRhWMVR8cqqNQWFRWeUi+7zSP3zdkhudwhv
WlDjM2Bj2jCdjgfHQK5LyKKrBHE12p1FpkR5GHhpPGtdVpev9yTOtF5W+8XjHh7ZgXSyraOJhlZq
gNH2Ka/mPweUTidd5IxQZ3O51FR/esBjufocA+YqUCgBpI7ri2jwXOEcg5rRbYxYMAPZqDuC32/E
F15kd2uuJAONdwbXsfOXST70ftzIzFi0JfFlJfndPVq/p3pe5CqL42lnijJ0IDxtBPVBe38EZM1e
C6VeINOshhcnA9CiOV3PVDL6sgyce2UJ7yjKNOktqDe/8TCfiwl9Dd93dzmEZWIHKaiVvnTIL5kp
FFMkKxNqThdLpNgFIFphgU5XOyYakttiBFliJdoVUau6o5Dp8qjktfDc9YvIPqSFSDB2dz4M/ad/
wwcErOyNO6/MfkRvFutzjMhTs1nFjjDk+NKISusgfOTfBxOWQdpGXFljs5iEhj/O1Ik1Ai8GUYub
5Fw0sKYNBzmZjuM3TuePUMuh0ImlPXpzz+22T8SdBLAabpA4MgpNajctSAhmd7PUp5cH5VpBD/Ca
w/PkbLpcgyQOcvODOyD0UnJ71JJIbIY288Qi1lWMiKSc2Zl2rLcsklFb7aTm9dan5Q3I/p9xRjtb
mqoTFfmnoONIsEl6LEmNi3FhPt6F7yPzjR2m+cwQLRkOx27snZKE4zki47I41wVi5/z8P1ex1fyL
PyRNe9JeSWtt++bfzWL2KG+U5qsf4Sz/ljyeJYPyaw2RgRvjtudqb5yR2iYqp4+VpjGHxApdlyuj
6lXw5r0uB9UmC6Xhx7DbstpPUBJ0G6eqvWuVFAyPKU97skcxOjvON7Lmcktxo2MgIUAJtBGgq9sm
8Bp5p4SxE+ES4Sl5ig4BoSADF1K5d0Wif/BxEF6NgacKafBh6laKo+mWvibHyqKBWDZtQ3Pcd8Ms
A9q1BxzYiO9fEq7daMESyjgswMbuNCEpKIxtG25N3a2IZtVIDk+AXEtC1f1GRHcJMS8/e0hxvWfg
1HIg/GN95H2MJUgYMeLOYvt3ROVNmJPBdjo2yl8zCKhdZqMru+fox3YPu45+N/zo49Q3yHWOouhM
hT9Ep5C2DegdLKZ5ZXRcNqQ1iKr4absG9ODeYovYkb1ttkypNBr8oAh8YyJAxRAD8My8HPv0fy/S
Ks3JOaw6cw0TA3PSL7Dxj2CU/nNju/a/oW13otT7fpk1XHca+H58qceNrbzs7kI0LrWLc6GxJ8DQ
YeNLVzPCftx5n//mQOwwoLWaGAGVAiNAuQeARl+dS4IxAgRePzVtMsJ5jp6jQwSPV1lr/JshuSJm
jH1QqrPQne8e4rgWh2e5WGzFbDU1EkuhfDP7cRSc5+Q1hoapdu7JVtGhcXl7KAG+RrqM3al7NciZ
pVR6TueOJk+K7A1vxKosomNdPUDyEb49ELLNl/7zMN876qin+zjZrdL/iFME+Z5CEF8kJ/872l9J
pb3lLMwpbqTi8qXuxDwp8pNFPjl8ziFYMqtP1jHv5BQ5H3mxXx+rLotFQiK9e+6OGQk5wtmfUNsP
GhQP5VyvkImu2aA7HG69fepPHkxQSWCLx4GnbPgpJJaCaLYKDO+zwGL4Zutyzzt32+gTxFHiDh+I
g2GkSoGceIeN3zzbAMz6VUrF+g03FLVqYw5tlz7eiVHFxVBs74RfmLehkbn5cCz0XXGyAWqvl+CN
lLeat6tcJg3KY2OAVxEhmeV+Hv2eg7kR5qOKSGwiLNvBN9Ljm/lYXArUP0xem9QYOBbNL5VEuGwn
ImPD1D1vbVAVgrwsmOyImyC7MWSwya8S9/LllizACN/Qk5s21di7cumvnpEnZW1Ts3iCfgYfBhrB
6xvpKCiBZv531f8u2+OPfedbouGSVwdCBRMqfCWX2AYvFlHfriLQ8DBQGus/CXX3i36rj+sefObF
DeLquQLp0lQ/zTZS5jaeQ4KZLSoNcpeOd8mfPK4trVLaFeMANVX0gKHaU8zm4456s/l/FHgkdTid
4zt+sYBe843939SzOXr2pfCfG8VAv0pcsi2X9ZjnVxF7gf0NP6+/YLCSTkXJVjx21iMzCPponWZQ
cjyCoVt/FmPQpibPWm88P+8l2fnSvqphZyk7xT56VQESAHoqE7DAuGUTlEh171RJw4nd/3I0HfRY
7E0JyRMdRfHCtnAGCkbgC1343hAHEq0iGNFpWYt7zRjl05DNOZPEyK7AG8V8kx5z/cC++UbZaIH0
U3T5pvDkYKVrLztH1t1yXg0g4IIorhcxjJm7Td1zC2zpGzI2FNuocWDB70wyhx0Cy375ACYf5Fho
+RXMxcgn/Jvh4f8ql5zU5L1HTCjuQGi7G7OA7VGLncjt+ut8ltaLrQQRCJTa6BrYr5OXgIw8glJB
b4Ke/g97UrfyClux+O3svvF7Jlm2m0fY8+58qZVNFaFG9Q8WF2BLxtKntyht2FdOgDyvYWdIUcLf
9xzL5wsVTGsiXlKV9JW20XgQOVrdiVk2ccP+UkLAXQz16Ar6dT5VrtcyjSOJwCXrGkmzt+/03hvC
iZVs0se37Y273dIqFBbCjm+A+Er8LcFG/XUugWn7+Uq0CKM0OlPUncQGQtsMuTsbga3pyNF6sPBI
dtSbymN8NnMPC0NoAoHJPTV0mTtbbIRpm/Ymx9btxK2kx2bhRlwtNDOJOhR5V1MqNWjhocj0TyOF
5M7xFYHU7XwciYxAefZLMwFKK/nCWetDWePg6tr4ct0SZ0npUvHOljZ7AsX/aXr48Yz8eoDl+2Gs
7DaMxw2lDMt+ep0zwYrgl+xREm5tLusqgx2zFKr4RZVGsrbqhik1dGsin+Axd5Z2LuqVE2fgZadH
6a4kSv+EEzLWhOy5bRi7jGY0IOIxxVrB4dUjRqUcxbJwYWk1DHqbh4aJ6TbBmGgxmUCkb/2SUXgx
f4ihSatgxcYay2nGog3zXwIj8zBmPOuha8nmkLWiYObBdgXFW25n/sIlZUHtre9vDIGgEjgyL6UO
kyeuSDB+bCGQV1PWNF//AiFJDlFpJ99SS/6qFk3x3SuZSmSBi67EKkMa6aYDRvnZlRilppeTSPeg
cLGJIWuxw5t8wzDwxBpO3OF/iTS14p+xjViSnjlTOreOetJdUhHqQjsU/J/rj1k3NQAw0td53Pqb
mWes4ZX8zGNAURnKbIqUHz19wMSrkHmsNXqBXQoK3sTpqg5dwbUMvntgH3ZLS1VtdZPilVCBdBDP
moG8puiJna4GZbHybV2Iyv6q/JFumHiblG8GSqPDalJZ7s0C8rSv7/wgKEbBWMp7n40tRmZ8bHXe
s6hqvAy4/p97vVg9sWSnvNcVOhaX3O4Neiz6V6DjTsR8uLb/q1f+X80qMuI9uK8Y9JUEdZLQNIa9
Kw0JznXKLBYsD6MKaIWrOM22YI6SxgTjJF7kA/EBkyDH8aIlEW1yPGr1gES7NR7RopmojqfBxxwa
H8v8jQoPcguX0/OeYDvuZEEKjRXGsm/jfaPlKrqCxBHDafsNAxAb6spn4AF6S7G0kxJ/sQ0OvT1S
E5aF5QZI93mPiZU324a9ExXWqmQFzjm+4LEJfUSS04jOyRcAHR6o4aKcMtS9qYHKLyE+GOBHY/rX
0xmnKBZ9tjjErK3fy1ePETVYwDJGLru4YoI7UDLhE+D14xe4Z+z+tU7nYSS27eGB1DiGLVJVHigd
OdqIrbL6Fu9rokiXAHDqgDiqBuQ6kaswcQ1hQa8R4iRvvu/VWkb+C/PotKgL/rt/Uy81ywYI1nq9
Su8PFAMH3Kr2H0kd3fzfxugp8q8HeQ+kiDKsiNbB/TN6kzfEs5Xl0Zur65RdHOC2/3J+auxduWwo
/mi3lANviy+0XkRI7FTwn8wndSWKp4ysqMVlM/UtPszGBrxBW1tEz/jlCYTuB5tXQ0RDhWyU87XY
wRX/0bnaUr+VN2JcGRwkqUvJnxetMOezvPQMvF6KvIp16CzR19QW1Xr//FrN5S/mcIgy50XoqX08
5n94bNJDVzN8DwYyVA7IJign4MBSpxJ1yFmgFRlIECplkgQR3Cnq/93TAB42PaaJ95esHZhGGiYJ
lkqtBXy6P1pRiEoUCcJWgLpKaq14ejQBC090fZJWA5TUFxexPnJk1t/R0pmReQ8QSlY/rp3QRSXT
mxfEuuiecbcpbKtbEGoWuWK3sWaypCO7aJHdfwc+aILqouqz3gUZxjZpzvd5xUJ71Px0HZwSzYVQ
HKhp01pyBodNXs3gk1M0fv0zTqt4QZFjUF8GA9teORVdU6NbFnIwc4kllKnojhCGpH1G2gs0R4bt
g6uYHsv4gycOpMvG6JW314RgoZDQnRzijxWGzisMVZvRXGf7ka7yZHskThEk51g2BzT72eh2gXH2
42Seo+5mNpTPTqsIq+maxjIHJXoNnhB6bh/G0m5AV11pfn82LUQ5nBmk18wpVwK3EGbSqj+9MT3Y
Z3UHaGTbEgBGokYAksFQSW0jWdqaE/RWW/kZjqNYfMyNPGQGH9adM1EeHj1HJwqW9cKNZzKVCF5h
jM8YpN0/ham1WFIiNId+ZDJBuTgMF/tNm+o2cFG2fIksWKgB+/HtDl9HLl2ZglCMfc7s1Yw/zEd7
L3DsGOwZrnMEFq7/nElej3sD6qdVzhxAgbdsvbLJf6O5xL4FCqw8digiM6k3qYDxRdxI6AO6maJH
Gi84udPt3Br65GRpT+Q10ngI9MhXFFuSnjuj3FD+Wx1jNpmvu/NP2HyFi7nXUN7uRDHi3x1HTnSn
lfkKP9glprQjBa0XEya9nCQ9qFMVi3EvGG4ov8491Evdne0tjwegC6piTxgF+18bmMpUDCTdIe5G
KF5QcrxG3McR4jCugUe/xmpvKCPPLprjI6uNw9lxXCPxIA7oA0zSFSMYup/ymXEZew2+mqdbUWRe
UgENQWR3ftu54z0LWGe2+S9Iu1jkOEUCRbRgDjVUHa9n8W69WR+PqlOo6oqoKSTjB8O8X6qWf5DE
Q6ejeXQePNK2NPaMbOQ9yo7WmCKcS0dPT3DdUfc8fiUZmBvDhNahwJHnJ4uSyA9nVOKsAKLhQrvz
R/2pZjWnYQyre6tiNcWjSJYSS/MxxfltaosgR7CUdgCmYI3b30B+msV9Ms0L+GCMLWI26Gqt1H4L
vDKgzhzBQxAQ+WrbXCq1ZiAwetF054homrubHbrVm1X5CR42W6KKEu/RXxH2AQ48AzeJPFhYG+lf
baQ5LBPU+5Dep7hDghSfVsLgDYc4A5Q4mFuXE7PwDdqh+cxFGZ0m3fdx2OrOV6Y6jJXKbWkbNvSk
i6NWY6QcMbzvHkS1wmz2E0tD0tGk3cB/JD46+Y3tpENmprTR78PZbmGu1Bo++8cEh79yYU7UtcSv
wqBBoVbdO1AcstsalGeHF1vkepVSkX0YIStLBFQeQ5l9yn9DeH0bIp7f6aSymA7yLhMORJikTn89
1xM+UhDQWD452Jv8dJFXbfwkYMezA5CAQFxRjmjFC7iskHnZgFFcZPJZFGsizZ56V5Va0VwHQ4HC
F24MfOBiBeGQZFErgx92lGQR+AJWOiNJUN6qpmU0F6WJE+ul12vEbsxMdmykGCSi7dZa+q7q0oFX
BiRHSONvMd/HhVV7x8eXpvuAuNU5+Pb3wafTWI0sLDawvvRr6XdCmBvvN3pcq+QxiXS4Zlj8bawe
d3CM221Srh7M+tJzFG1AwxblwT3idJG7HwhBCvDbBlS/EH6NQriqQ7w8sBS+QxyswC+67aHsTwka
NuAPGtV69SmE/QBuw8GoiWUaR8/6aDBVrNrX9mO8ZxjPBKhCYSLV46dJiPFdz0Vjs0NlspFharM6
L2KiP31NgAbEpv+SYQVgOzeQaOvk0gTe2DyMM6SgHjCl0k/Cx2dYngkFiNcNem/0sypG0iflPXIW
oTpY3ktoJStiVLSG4PGoM2670I3iEO9SW4CYEZKnuz2SO6jr97syy5RfhcDL9lhLAtRjLsFVUKp5
SsMBrSSUsXz9jotHmtzjtrRR36LUEew2enSKNEBR8i5O5G6vqDckxw67D/TcYJwJi/spR/k45P3D
eu9MClTmCmboPIZuVotH6I7UlwQZVhGRq3mF1x/MKysPUGMjHsxTICD1lLerkyyIsPlG07xNqptg
E2pBwk+173L8eOagCwRPfq434AOjwXJ0DyfE7OH2NhZ6cvChBNkKxIRD9djo+F4U7i4jNglfVart
yQySzm5WMCLb5HQ5tLsthBO4iW0r5+7bAydFm7kavEb9K4tO4nccW0NAQYpPMdA+DNS5CbL+H5Vb
gqaExGYphaaMojruXkIgHAnXAc2Z/kCA7dms/KJwHSvoLAMsGbFahIxVnr7J/uwT/gagO+sfS5en
xI6DS/6BZ7JQb5trdEt1faHwc6ziQiPdlXnrHtZsD/hlEgiEBBVre+maoTVBx/2+dQva1WGNZVWb
G7+0hUNC+JCs9DD9p/2nC2tyURHnFwY+ZwI694ipfQCv94e04nF0ZzRT48aWHmRYVEEG8HI54TE9
XicDhDI49PaAsDU09IfAN7mfvj8eltpQgyZn85L5nSDjWZJIPntJx2ODqDsBm6dh4ZIu+qLMvkaF
c60hczi16fUus+TPWnDfBfP61TB+OIhzohhFzQpMkltUFO3ZtvEC2NvqHa7Qqa4wpzk3tj/viS/r
HuVK8y1V1QCW1apyIl/pia/yW9lBASUN3pROoUmXebQYIXyOeXGBhgFW5oKiTPmLPSAbAeonyEyD
Iu8xi8ZI3uZCenr6ZpaR/zIMu9y95yebY1z+GQrTRrX5VduT0JoeDKFTORaSgUXc8Q15QE9QZADD
SMJc4XLZkaBgchB0KyCv1+FWlgFhmPmmwXhh+ZwuCV3VCQzlZhjVNoF90WR5RTDEM51/d0PR0Jl4
aTrrEux2lX7JPtNxKpZHCogKnrrhG6FwQSSxjHj/y4/9cdZF8EFBZQ03utAzbQQL4PtKtdLnG0UG
7PVHbaDbGjncCUS8J8hzKU/f3A7kH7DFujoZwYX2T09fG/PRsIumJC9G0CHNH9RHYEX1h3bNZWpP
qMFlMpmx2IWu8e8AXevC0Ohs5iSbhYv3ZuD+XIpx26A6oL4z6OtKhn2hKEJMC3tHexaiX2r//niM
yaC47gX5Ryoa1C7Bu/xmvKNbMLJunPeihDVh5LEi5Kne4tR7AI3DCmBQ2DxvBNq4C8ai3L4vg34/
eojko3PE5B7uZwachGyFRr0jAuZ8ztBNDR7PJoLApsp5qxk1yYux2v1Kd6+KEtaVySwWz+kCmeco
obvCoWQicqkAMsK9lBOtj9m8sftytsCuTFT7aIY79K/NUDb/wZSmGkJf/pHRIO5eVlv5cmtyAgws
4JBY5tHLpO0cQBlVLjWRTXxf1dUX17abCWlNCI/EdJc0kjuaimOPKeIdMyOH786kLc6L/v+2Z0Vd
gEN46QBLjLI8Fofdf6BE/gDpdRbnlGsZ4qJDgfGq2SuM5BHLl+fEYIFT/vpHKevuQvUDkO/YDz/I
RAsV7GhrbmuVrVP1GsxgHm6M6XOLRaE8q8W0/+56Q2Fb1bOjQKKvTZVEO6xeLGsGJ7jSZjYOql4z
JmcW/Y7+U95nfvgo8qJS3mjk79QLwqdW2zX+sYw9JnAPUJxaO4Wfqcqlb/u1rr0sGiMC9Bo7oAih
TLU8ryNUkj31oiNUFkLQh2Sgx7FD6JorYiAfXwxJ2fCPY4pp+NcgWXfrORSyxJsX3+2BByjhe8l1
22uUCya/Oz1plIyXU78iHUpCcXFNFoGEqFGChJSG4S8i61tnXYqJYRXPx11vb2fssfrWYFB/ZUEB
iFVq69Ep8e77P7YSyfaTMtOozjCPYKfMTn3B9v+WWsm1CfPpJnf0A3JClJBH7Bj6eYKQ8pX6mApl
qk9f6wY9lvj3ARA1IUmhKaIOxY4GIJJ8X7Noe8fld3FdPayNFWNMMbnjqLeCgVSYXo4PpaJA1xVR
lzvQ+NE7Nyvku7SvxNE7QXT7SAo0AbViZ5OSCwVczV2/FAHr8TtYCI00zeUpWkCM6hbA4CCLkSgN
KkQzrK38ex5kL7Bj51yrbDiQFsvhlk18JaPt1Am0D9sEhRYUgRHESw58Sfii2eEsFR9YjeI5IZdf
XjPPjx/l0TxjyL+MB8ePCUX8bw0CDG9y7b672oBp3r4ETVX3lMLv85lxnGJ2rx62N7O7JCC6355Y
kTaDrF0K+I41NLThpEPaSNatFLij/Lbz8sXORU+DDFWUEjsMEFmY3f5x/fnEpoIk7LjIxGYj/YSQ
QS6FmlyQzG8P3ehQapB98gYUfSzo+iSaI5B/iqsSGGtawJUAZOgi031CGmEChW8os5YIJDq+p62H
/FTA04D8r/agqDkgwqbSnAMXY7hytzCJQ4yA/z0boGZnpuFv7R3dSTar+1LdLxj1NvLZ9Od1N3TN
F2dfEow6c3A7eS7jIsOxWSiRw2HOeETvFCtgLuA6ZCvdz/TLXxeTE1aN3EtmSYH80w9cb9HJq/PX
0AeLNj02+xGe7CVVmlnNZk7c4vlBV6QGeaKR969VS/b4RRWdaUJsSr1rjd8VoF3lOQ6prr8X2MwI
8PJZNO4zJN0kyJmfgBcqWbacV7PxrypF9OGgf0+f/0eYnqKXIGJNcmTsyScJJqPjGJHVFGxnuFX0
XBlzXWQGl0RuEYaew80jp+aFgr5o+LrOYeZGpUsK6tPz+R6Y8IPx1QwjiuYRQXX5mlG8GbYyvaN0
gWEqIOfJ9DKAmeOCosEdbplht8Ogv1ll/TsbyL73OSzrVVNSjKlpWbklqUwsuN5ayzL9VTFlRiVk
ZOJhzrGWx8ooDhKZif3wyBPlSpycmeNzmo86uTSiBMcjQsfZ8UGzLsCq+1fcfwDcjlO6rFawwjBP
3mR8biONa53aOD0nbk8Rh6gnBuKZNVo0FFBarKP+G3l9q9iEVFN72CKsWHpyJJ8r8AuczE5KXB+h
FbW0VF6C6RzhZfN+SvkgscoDQhp0psPJR4wtVjRVu/XkbiWVUl3pWc+u/5GIzuCszgBsSxZJR6Nu
99RtQmkolazpoGqqUZOSkpUfq0mZXO4nvExM7KUXKe+dpQvzo6TH2yXYq2vo+56rGESiKjumZ3Ol
z76XXgt+gzLFyAnQKfh2ewtpt6Up12r0bot29kSZ2hOxluTY2jrTUGOv0IALx0yaWcAuMP3PwP2J
IZgdRlf2RpyoeiRlxiNIYsyEMwFf63bbC0uc/Scg/H5fZ1SUDQ0Bnu9YaBNNEKya74+Q1A3YvlIo
pbKwZS0hY5SSzmzoYDE6VR0PZ7HETccfc1q8/fEOi1r1Caa59gVq3fRbf/H3i5LYBwRVHKq1QAwg
tT+7iuRm9tjVfRseCIadrUfnt7aZeFUQBrOdrNO24kyxVf3xAaUccEgtHrAekSKfgLNMGj5HLjwy
60M8IBkPmHsWen/1hN3NqeFi6H2/L55tW+fPMFk2YKf9eYXLiGN4n7RnFmVgGir/z3/5Zex0f0gV
Sd5oK4TIcKHxU1lMzhHvGNA1iNQiAtKmUkQDLGmLnZkqht3uLXdMh7+M0H757PExvACweg41RQuL
6ORKXhETzozzxKNQNxlJIqHreqePnonn6upGbjLyDR6REicAeQjgJR9UcLx5Yl7TzWwtcCIdplU6
niuk8qoreDo/1rBY1QpPK5NvUuWT1Ja2L1UQGguqK7HDPHiWaMk0CJpyDzkB0YbI8Gr6NMDVqGJT
P3adNjy0TKvG+2dAmifRAxEJrCw6XxTTc8n19MhF8lIkBuwAInfTWu6NuWiuDQJi1kV6GIzyy30S
yQpenKBy0ddgr2TRHGz3pqsTsi8n++DucDqb9MT0tvy04D+6rF4QBkP6FEjOrnH7z5Fu2wljNMFb
JLdowGQI3U9j+mwZ7qyXbqCHUt3SZ/AvbUlGU4kIxkBfiP3OM+O8BuartPR4wwA24u1gpXWT5exO
GfkDoetHdZSf4wQWUbURaHZ8SdI4skQAn8iMjVFvimhWO57bCBZXmE7g16JWUjXC/cxSmZ49v0zG
+7Dbv6AaxnKa1Y8nqR2VRcUADtHJfYYpg0s2Fa/dJv+lKajy75Z6hdrdyoa1rLnkstJ4iq6uuTNQ
jE6LEBY1u1MagfZ5Um9qopbCeESaAXNFAPfxA63gHa5VTwUVctNqiRYQdSWdyStiKr30J6XScW/e
UnYfBPZdDBsbchi5QTqac7gcxQqjHmySJBGscP5tWz4qKRPGupejJuRVIegHZLomSbzb4xHCCJNQ
hIvXLB3Sk9MJg2yo7hqJy/9UoMMmfKyORJTkUtRf+0E9QMDzvfMJHF6tAluRyhP6qcwsA8lAjQ/k
sn2Hxeq+jAUpAUvEyl+6vSwahDNrlT15zScxJf6mhBb/MX63jbGjVJQIieWNwcDi/CtD07RATWIz
1C9q2XmXVd9tKVBtHJA9A30Cb5mahIVMht0PkKrNEFutK/GO+n5RtGCQ/BN6/pG2uWoYBDc3xJUK
WMZEbeM+dqmwBwM14WnoO9mMMLg6Ya3Euj7dQsSx0llun/zFqpKa5RQlpZ6dX3kXtpeUJ9ydA8/n
hvjulvaIARMU4RERaj+hh2bNHAtNiCg/dV9zYJPCT4G5scqSp2/Rnhtd7fN4bfHP67ts6mW0Tcyy
LGKjMMdu7YfhnogB7kOydP0yz72yNouxuOVY7tmPFZt7kOu4vF2cLaEoB6EXqbVj5nCwVSftmkSq
5ubaz/tJBLTxQDqNirob74qAEOGCExNzAAV6vnUwEhyCL5hqMhzAkzEXqvkFT/RsVIfZCdr5J5O8
ef6Q9kU2bJ0TJJJw/ArHYe1CHcFIfPliPHxw8vF2q+tbdVeTG6cXKYLDltGpABNmpj9rCpg4HSFs
2uJk+atUr1MnDMVkgaxHW4ajwvO4hlCIAykjUHtuczk7QgE3nzt+PT0A9OBAy4zjb6gx5tNcVAyD
0wLypm+bIkaX4aJ1vLmfV4uMU2C6FpT/Hn9IIHZ6VHhAOS/F+5+3U+Yw7kbpBo240ndbsVG4ddCS
RrmO8f4tTHizuUMUTYSFALq5kAywNBaThGpdXpM8TNlXnGUJODTFxA7V57aLoBTMSpnUFUA9wIij
UOWNNYom5LMsu3X+StV2d9ckzt0308bMhNctyYUSkz6CPBfDBmSzzt4qMX9h4nFAIkzwJLF2kSpd
TNJTyH7tdP+HUNrKaaS2F2Tfw+JB7wBKzyp5BVWMrFYKTQOHgEVGrvE5aTiQ/QcjcRc97uxr3awF
EpI1BIeft2J/XIXZLR2YvGGndqeSEwa9mt4Ctb0c7VLS4uUfR4iNibyF5liWSmg3RiAMlHgr2VEZ
J/MeMWFGey0nBktTC5i07sZDmSG3FmvCpW1dOl5q3SiD/4MMSpYDA9dNgPLAJpzF11V9Cq0gB5uR
K52LoDZK4G8ziAYevenFDeqQow39PmLJMCqp7CJSXZJvELeMCbj0BCcEAwv3eJOXPODAGLVQIyzA
QnxtfFIIPkxT8r14mIucfNomAyyW7rpnt1aQ7FrOgLK/ty0o42j5mMd+CcIgdmFXhA1i3wrmMcjW
N2/n8Nuss+AOO4ilASu/Y+oV4MPoxjEFpvCBnO+0K0sM6ep2krTLethc9aWc/tgiQIMFyUdSFEHD
Ss9NdslsGQTinxrGP+M2gkxwpljtq47ss4dDN1ZPav/DdSBeQoWxUWhASrzLImb5gxDPvoikbAhu
nj7gJEprd2O7o5OBN7Ex7tOdw0BxT1Xl3wlJU7vuTaMFI2D8DTFM0B4AlFRcV05zfnECXu/QXMtB
PZGJmuj9ZTstKj0KaE4U5LjqwziaAkxPMbUP7nOWaqE28DOimCRz+irH0BFnq5sT7alYWUJWXWXP
mpf8qCJrGo/9hLMFULvhjTmotNdC8B3m5u9iC+N/qviWD4nQeaatGM+HH1qnG79i0hFUW6cf1RA1
7WauRgYkwIwnoqIay1vHeRyZfLvoXnZq17f0QTYZrsIdoWxg7UZ6hKmYzaOFtN9StpCYqwuoJ80i
Foq5c1+16F7n1DMTLX3lBTBCyF/DekwnIjh0TN3W8s0+QBlpSSF0iPS5ZUZdIKOKJh33pwZDBhxN
eEzNYMzWTopkySTlCHmE+RkW74f0ikBTyzk2HVCsk6XmRdbqjHBbDQp8QNpWhbCPA3/CklXMl4B6
SwEAiFxzFrmHQn+eZqz6trBat/eNn99GsST8HAmlPKiAPL8m03M/Nr8T29FAXC/kc+nOAvPenn8B
b/0h48WbwBH9M5whKIvtI4f5NDMFl1XfpkQIaLyl66idaDlQZ6dRnb5vhohagH9gR9WHn1lvvvtS
Jg0ILP9bs3HCGtywfYzdwcOjWBljDRYRPJbNL+gzA8eeDIpb8hw7ltJQPn3ZN/0+7jN1FBXhpFaC
DqCoL89ZG5o3+tDiHdAbj1PERmaFNbG9Rvbn5ZBhpRgQw/RWuR7HlfqKY4tfcV0lTR0cU6rP7pmx
L9TbOtc2RYM+WAxgXtPWKtG1hvQcpI6OqYXhidWE5jd+qnCnA5kZq6LyZx0ShIcL25Q/5XR5Q4Df
5z+dZ6Tl+eJE9Q+kZdpU6ReGfczGMkNVG5c+Zt2i/4JJXuJ4bnZJ/uh49PAw9KyYsvCg52kxDzL8
QGTlwaLiM022mNCdJGSIQHHzLhJK4U0x4OzaFKK+OmHGBxpB9Xq6pGk1mUTMs3r42apvQbPvLdcC
GkOoll9xijBoplAFPYddP/FXcxpwDNMoWYvIf3sMFLkh99q05S114/4Arc0ME3MNbUgBp1S91i1x
3GN+f9EFxHILLbh1WbEDtw8DyhZjExlZX1NbaA0A0F7XW+J1dPyC6Iqxjy3PQ4sMeZXgoqX9N3sQ
Nst7uGeZWHGCAVs52ND4od4hun25zptaklwz+4gB8l+Ye5ySsJEETjVkrjEIUCFFMNwHgNHekkJQ
/gWTxszinMZUv1dZom7sCCzwrCxCsU9tU3xsW8sWnijrw7xvu3v4/+cmt6t5dhsZDQddaNn1UsbH
waIbQlhkTsVTfTb64FWoDTB9RAYfk5VOwwhb/WJ7LzS7XKL3KL7pdkRlcd0jWPlO0dwuqqz7waL7
jLFWQHgE0Zp5E9XPOUp4uIUdpQzjU+SlvtMZiapxyu5pmuREZWBUyMo9LKpXRlqcYxbuIPJqJcGT
acPn04Q98QVg7TczpgHeCZe5h8V+4/Ai9zPkmXIIn92MejAQKSrUSbnOJRfpqETM/FUMBmGJnHwh
LUGdgdiWNnQKFJgoNTxnRlO2iLUqvhtwTeV4IGXqqEzHWIkbuFOFlSg8g7f1jG4JGNl7GGTzibLM
4pk81R0fvWu5mi6WVPKfianswlxQaZbcvi87BZngi/3SBg5hUm6Lfdtj0tRMLV1zmXSF/DnGaWM4
lsMrNnGGlM/hDQwEXqgChXBRhDREvJ57wA7ttSnZk4GRMEfRjV3JzCrG1kbucHomtVQYk6tKial5
zXPKBlBYK9dwfwLczKH13AExTVUz/Rv0p+KyptthL0JiV/iV0IzfuZ+14chXRc/4xGv4x81n1gP8
EM3qQzw5hrVCnyBDAuYmbUbkzMUVtMoOymeXuKMA13YyItj34TIwAb6tg+DjW9hxJcZIk/LpxXmn
O9vqkx9gkY/7d8YfK7yztd707/JpHQnYD0sSY/juMRU0vohEIGIrwwRwXVJ7WaUhFNXDg7u352rh
oVQc3BnGOuJKjMed/WhlrqX27cVEwyIpOPi8+IgLNYBSc0p7igCfYow9oAnIb1Hp5mSGaVBCrLu4
zI4KtXCReLqz4NVNRhFg1GdlDGpFFwGDcnhjuDOQ25s/PlWqFjtQwfx6gKy8d2HPKlEOEwtj3Dsm
etm2+7gVufI6EYGuI0kYnuJReaoXJFPE3prH9Vwv4wSMPRGzfp9py1brbPIOqF4HO6V0CNg8JKWa
mwI5yYWgzjz4JgmHxmqD5QaMV/UInpr9e8APYNUmYd4bF3FGCVkg9FEGM5FL/OpYBwdnKe/3rv6R
6APzdIEcMqD/IZZSjD1NMmg1W8DS15c9Nr2ZOFc8NHi79FgI5ofDbZ33/7QwFrGveb6rj/dJ4x5n
fDc9HOtWRb0wwmrt2UxIdtlV8NyI0W9aZqciU9qGcvtBxeb6v1kCP/lEhXiHz36D1Teu2B5yZx9t
ESeSniskf9pYcSbVpiyiNCMfiRd3qb0fb2fuWtbmCJKHkMARHqvsXis9uUkn1952hqA/hel8p/SY
oyYfUPBy9j1Fqz7AqicV2Ts4Ld3G0ZqrCJvJxcxWFL7KlDVb4vnKT66NIUTYuyepT799xSygYAGy
/q0wSmQrpIYA9P5fGK2UU+QrwwipIvkhM4n0/trCTYgUt3hjqd3/Q++ef80JztOndC759AhMqmbs
A8akbX0lGCj9V2ZtnUad4TtcOOBiwCis5EhUOvMRggMHhvpltfWObqQiYLQc7yQdYFCEAize6nro
2DiyhoawQgjlCsdnI3zlxPx/EY88IRoKNrWVYRaYKYKFECyU4QQz4h3zVbgpokaBa+UtpDuLB8Iy
eR6+3ye3YiFBTk8mXGNLOa2A3c4xfXXS2N5Qr5klz6wPVpxyw/qZoX+Zz+X20gmN/l2E/maXUBAc
s3M1m+phqmlV6vdCh36w/OLJYsOquyIzXnGOwLBIS0ReiAjz+qqNFR3ggXrnbR2Vn9yy1558rosX
bVJd95NxE7PcAHvk495j/Iw4VjwA1bcz+QW/5/q67CI4xONksXzeZOH4M3tXy2V0FVXJd5rR+ktS
zowXGX3qdRQbCF+MIngjkvxWBXtaydeiZ2JtZ8FfTRw5ToC3rVCQmvEENzNb1JspoBTQ7s66AgzB
6RIdfrUnYp+kDqDm6DWYGfeZpdWNi9/ze94jZA9bB7wpKvVtZnPADaxYIaKg/FEbtxLUxIaBdlKL
eycK88wIBZ/q0Mtvk9bExVZwLYtikOXO0cWM7KA1zLFK6QM6IcxWaNUitHnj5DMWWgI6m1OJHB1e
FrckUJ4M1DR/i1V4l20vJ5vHpLjWR+HCP6B2GZLZt3n/glpqg5hqMeeilOG0TggjxW3Z3hnmYP1U
RbWWTW21YTZLcHJO4uBHVqzi1a66ea/jOe0TfrpLmzb/MWOxwId8OBiz/6xxzHAWeIlPVfS457hs
ghSbKmkP1ngWhdnW3rfHAqAOA38tBHulvH2UnQzIoSzU3k/FhDfokZJwbBRnQR5wd50IQnezD5Ut
4l8V578I2mJUgdanDXWZB7qRsg629XySbjmGUUxB13b0RQbKBbyeqBxrOkntX3cs36NV52/bClFD
fFWe9BbCg6mPd8JX9ztDBHu46P9LI1GlIFScDlAN/JvK649hmeLaepRk7rkKKCrJOi2YoGRD4qXV
L4kio6FI2E55T9jLo1FGu2oVAfmp/t7IEfvmjhIBPBSLVYfIL4RA0kWL8mb8834QCaBn+0b9kqFh
50olRy/nYVSF37c3mjrVOMUWl+D/38V7rzFJekq8VhWG1WY5r1M3ZT53qdEy5CS0D7sGzRygpKOd
wZz91mJeeAH5G13mipdgCXH6Ho2fPwHydIb/L7RvDE7rFIhSzkszzMwmR1DS54mfiDViPQvg6sLa
o6eXtesihKzs5fJg0S/ZeZOtp9W2owx4w4HORvkff+w/s0aeVGVR46a33StR4VuOm/SMxN0BjU4C
p3/NeQO0A50slkZN8O4l1LRGmrMP+R3T1e93BnuxOfGa340Lf30DS99+bfDsVwmPMPeCtg/hEMQT
x8kMYc+B2JuPgx+ipheDeAwHfoloc8jVCPnmKcU7CwXXpVd40TMZONZnxSkHY21ocpnpD6QUH0yc
xbUmjTxzWZRpWkdGT0WdYJdd+RZPT01qUHaMyuiVEuAWGQ8UzHON495HW1fjTDISUbfuPG3bVA7D
DB6RiLRbOBKrFILn6ox6ZsUDXdUDkwE8kaBJ6rPUxULO0VpvVp96YOP3whG0r+cw/YlvWuho1dpg
k+Lv6lhdqDLk7moQM9oXFLGiHylTpI3+iyi7Vki1ucIcABAGZDYL7Qg1UR+zoKkcn99AwFhQVZ9E
CDFJq6UwouZ+RQaWj6T/k1OnmvDqubE35fwLMfVMkPMv2h7e7NOgLJd7lPE9elwFDS/t8+L6QRd4
8725uNp6QXqtmnOkgYRU0O9Q2SB7v+CDOIjB1/GFfvfjz92iL3KT4xPrQBL5w6Lzyc6WRHOGtz+8
KLbQKj+L1335M4BJk+qKeHMVQKCYcteCcH1Ov/tMB6F7R3MQNxI1BzNJxkAzSRKrwkviQ4iPFiFt
Z8oVg9KzCkFuOu7VpZHg6IsH4iVkbINZSp8LjaXJOkHak1NyAgGdwXH/+PLmBWEaDzUQ5LU4CV9B
rOpocr5ZYD1Fna5y9ZhqVURJ3sX97DRafKA+/9ZfHx0FOxbawQwEgUw/GbC5W/5czHQPiLWAk9to
uotmZWT7rH37CqvHbijrtAmKjGehz5uHq2y0mFRkHe+CDogXYKU2L0xyCVcmQRpiIAAJ+3vbxVZ5
0Nw93GSwq7XAxdAHvg4zlQoinJuMEV/dot9XOX7taFoLhQObzfDOrP5K8pezOsYZNgEkf8u0Q6zH
ZIhHMxp462JNjdkqso9pV3VhBi60upSRVu1QcHUafxqSQnEba3zhOl/A98B5tHPBh9yO/Kuhb9us
yehqXyAls2XHwymDxof/i4AvXgb512M3tWGEbiGAFf4ZIcchL5vH6nITzi+v/ip57cnQwu8JnbzR
c+ETq9DlKsjGwaasHoIswbZUed/v1JArPRpcEF1SeBLMUmFM85NY8atB8HNARrpgxUu4oFizgGzq
WvCtyLbRjcFzHVsoHK+85ckl1JMeFSLEddGrj4Za2NB7xsY45efFa+3CueOom5whasMcfo1/A9aG
dgmGryQX/GGCth2e4iuSioqcNNtxqUY83hDAsZVcFWMDaSh4qKlXngSl9AVz7kyn83Z2tMTc0r0d
pNbScrI2JB7t6X/TVnf4Mm9dyFA57TeKwg2jRQ7+KTJt84QInO1dss+1F74aPJkZvyJ78WCpv2ii
CR90tsRIXs+7IVbqdXty/PRpvtvawlxse01JI/PgOEPwFxyUuV4uN2Wd7hS90DJgBCtoBziJ5Cdh
sdMFOPgTU5HBxmqWoKyzebIm/4Jr163dHmcDmPURED2R3nWhP0cbinTfQpr0Xv2NX6CtWxO31ZSs
j5TJACpTUUMSYD3BMNb2cfn3LHKVkBSAVxLz91jBH+gSHF6xZEzwAiQbfPS6BzCeU/cdO/a+KuOd
sBMc6nG7ZLFOMCtn6a009gpykqnQXbwxmdjlpQbPpjNlEp/db89zEy5H/sr9JxtSh2VOAIeRM+29
ZNxE2rWsZbMyQbygETXB7XzVmpTpcT8hvmukIlJKujr4h/mgKYW+BKEYKLbpasH/2IJxapZn/nsx
zvcXFOtvnVk9WP8O9aePDhTqcMPIBzSEiaxJZIwEoKpN96k0Nf8M6OwjNyGHo26rRG/EX5+EYhYl
O1HBP/RMaFWr+TrlEBgPsIqIQr8CExVNUi9YbwjX1VR6L8f3NjHYBXQaBH4xH+VXjq415L/lI4C4
K/yOjnCyoygEzZk8t2E5kyeLdv1v0RY1LDSJP8+16rFcgAiN1kBWS4qI4XkTY+CRZHpkorsMbRPv
wr6zdtFIuKy8DoijK/56t/vMqg3DR7FKLmCHxfk7wNTC4k/GWObEb+5SO2FMcR5IFt8SkIZ5LR4l
Zl+wf/Efrcx64551lwbxVD6ir6oysZArwbeW8eOlCPIQ6SvNzUgdTsurqhGTL6JP6Dq5zLOn3S3M
WUoTxqXCnA7QQcDC3LZvkEGKMzTMWyGLsPHCD+CK9lNlVHikgYzjmwL8bSml7gkY6IrgooC1K7eH
+ngiLjW4NtLH7Zr1Kbvq8OG2Uw6sTSpPXc/FLgrQkZgxSbRRbkGGifP+JMu4MJoBHy+6qInPqUkd
J3tFJzNsrREFKSAGnyKlBq0FY3YFkGt1NEC77ZcVKW3fU/FEuh1gP/arPP3QuctK6ISkatKMrqto
XFkqhT7MfFKk+/vIilcEF8wME/M1uyJPet4v4TqnQ6N5Siozh6qwWYfqbsWbRGIqEVQAYCDW1qFz
omlIIomKvPctouivPBSJQoMDNP3IM13328NDAUqW/tuhTj+gf6S1gtAHbn/6z8XwDdSYgHjjHyiW
v9/r5kLUlp83p4duZyiUf67I6wwRRKuvFcg1VOvyRwuJ/OEq66IADEmR9l8jLAX9rpdoENRjKF2W
iEfHF6HxdHMrYQsjINwtPQKmkFdyTXvqBXiuHn8nQow1Y3ZMMR9cHAMrUYnJhwvH32rB9U6TyBU+
sYnhXpmxDMpQfdS2LsMC2OafuTW0WAtlk0wkS7xcYRzCjbZoWKbIOaH8R2rv5qH7CDuArRQtQk33
aamvGIVCHx1D1HpTE30tGJOKWAvsi1QoWRpU8sSOT2nO0pePlNEAzxMruKEIrv+NOZsHU/AELRVJ
i2VkQjaNy6zandGTuY0eRrbQSIJFGcFEdBQOAL10A7/IeyirvpRtjWUFsrLusWuG1W0oxxXqgf1g
0eiS+KgwOMdlQoAQAULaOPIj7n5YjoySuklo9T3p2E+0V3eEw7J7fkl846U5l+Z6yIJN0dhyE9vp
EQxsqgd04PLJBKwEPTJwyKr9h/AQduSGoSMk4c3QjbJadHSlvufpj/MeDsP87NRxhzzTxGmnsn2y
FHpfezYh4NWc380puG7TaCwGw1R6jI8Y3BfjUqRx4HjCyC2gc0YbqYLuMhtwjqyNG9KZUg5X+5Kl
yZg7cobhZ0TRaP8rPxXYwNSzuXcAXbDUCL0+vFcSrT/CY14NEyEITPDJIabMoQ/LNilxBSz3Bago
H6ZPIN1GyLceDnfBo3ggVcr+fHCmd7R/rq44Ih3L1UUx4ufkSct3Ddit8Nab7cbD9N/dkQqPwlRY
ViGzkh7H4CTljEfWM4S8CayRlhpin2XB6beY5HMT/I41uCx8tnaDsj3y28OlPIWeNgak6bV4rjQi
RuhUk2wnM4ECP0oe9AFqioU94Q9MQtWtXPSpxYsUM2kGUYHgRXYEKhJU+ZzFPIzsQJc8blWgGOid
91JykMP99KCFGnQ2B2K8T6r5eP4m0uz8u/8BeiznJY4zHVCAYiGatRITwWxH5owXCVmoL2lkX7tO
Xv6xBGMMl4GpkofRdgW2siqPBGCrr7abry4MfWjRtKHXVOI2SLfcNPhle7pQoxrEZxv+0H5qmwzz
HvhLhY3Wtuft7d0BAMtDo9cSz+VEKpe2QYan3MD5R7jqfbRf03ahs4+XmSpLNDTmo9XoGh6XDHO1
cFSoyAhhWdQ4WJ7ITlTilGQ8ar698yN6n314K44xgo9XffKbWaK1ihOwHn5lIo6HyNvag9W0yrxJ
nI/qOrU24OdgfwSosJF1d1HMFIbgS0vh675nvMJ9POw43jdnCye7DnTmzEUoBbR7nCTufA1xQ2LO
M48bnF0rmvMXtahuxukg3QMGcdqV3S9U1CgdN2FnjbzNQwoHMuPiD+kXCC25+i04MpaCSG0hrPUa
piclORl1PMZ9rdOqfUCpXvAgdX8X94tjLczXOUvocsFnt/PtCVq2Otxd+b9owYKOmkpNPuoRXnFc
DCg+yUrJQzIh7IZpWJP1us/YO8h0LUstanpRBcimPANwz2xjm9WTpGpSMtbfOAx3tQlI1/CYNIOH
wIO39ql0Nm9bySLgSkABvJwGDZbd2RFlxlhvyogzcDHyYFIZSEmo05G1AsXO/lqdw7twmnDE7lU4
sys/MGJJK8JzJ67pknWAYD21pM8doTBJUV90HTbWzqiut4LAAAlPvRcvj7TbS+4y9mz+W4V94Q53
9zfOLowbCH+uLeth/01GsrRV4w38N9DkuoNfNWaJi03cjAl4BRPJ+IWwV4WEEp2DeHy/DJwiROG6
/mc6nOesuy8C1VnDNXKwoWeQlk9JKiE0jYw1JH+iq3ly8u9R9zMBsnFy4xzlIulXfx8diezEyZV5
aDUTf9eSvbw9jJbBns5fl5irnMcPy3AIbqV6R3BjLJsO2h5n9FvP4+gTgpNm0k2oJVb1rG2w+RQP
lH8DuQ4JMscdvclGqK3x7RL/DY3HCZN73g+jVHTf88R4k6R8d0tZgp5Jh3uQ3kqsE6hoc/L4H2gr
ARG646dxcaX1UkU002GAXIyvP3lTXlvPR0gY66FFreUmzp0gFGlSGPBcme9mCxLXWUXuGeg7w48R
wQb781ilSopKCP9gFf5+NKi1hJgjA9Gk+3FcokwUhYaaMPiqJu0uLEyIHPGsefNOOQuez1ndJy5E
0uoxidpdnU6yIpuAGIWFeGlwjxAcWdFu7XJ0ayXRl63bb04sTLvmHBS9eDb9ZF7JgU4s+V9+DxHy
h3ym1L41bge0q1u8WodBlCPPhGmX58eEeGOnUZ7ape40eMVv+dFmXgJ+Pa/ZVG1MadzAKrB10VZx
IMcRVWGKmJDK6w9CMnuEinQp7q9Qt3KrVddA4KExxKV67sVlyFlf5w8jLCHAMWcBQ1Lcm2A/zkKC
xNAljATT51SQlw2q8JL793lNT0zt0TCO1EPUag2q8nMNeGX0R5duAghjwhHmfwjFjfXVnmbhvVlp
nhfvUa6qHjUgLoFbSPZoI3vkiNX6mqzqbBQ25WFaAyeEk6iII6uxO4NaFQX/Vwfo+ZlTxIKBj4b2
iYGD0VnV1IcmiVqQuI+C5drDSLeqaxkLH8F72PQZFW8HK/9BoZ9IKv3AOmR/fmwpZv7pgejd7Eip
IwVPYGzYxtvbWtTy0plwnht0F5YGp57VP2OG7gLg9MqKDCm0hc9PNHVlzU2MGWuVeRUx2K7H6EU/
QDSXC8SvUbe2OzxPrHKmhses62Z1XzAQJKj3BqHLMDV1W+saG9tNa4FsRB/fjljPhcyV5uN3DEli
MA2oP6UmZcfzfcmQq61b1qAG+Bj/+twigE67HslHusnR1Qn5wrX8QoKCoZ0J3rDlF1d1FNSnfZst
0AKMRmnL70uMp0GjTUPgG1UqizQdXMQNl7tlMH9e2IAxYuiTd+PrynAPzzU/Qg5soR37kyY4yxkO
P1kJVMn7FoqUNup3WQJhMgbdFtAQ7AHnMzQP/5Ogb7QEJ5RGMM8VwBzoHf9UuH8e6xiUgnuXLAy+
9z4F6L94/ZCtevn/7YwYq9a67wMQQkyPkOxfdgqtRmN0PTwsr5u/gbk7WXmmhNEhWa97BICjEgPu
7lzR/i5XL7w/mfsl0MkTYgZs5x9z3wcT4rTk9AC435zohX/pFzyHIuUx+zyDtSa8gICn/0NT74I3
3wYd1RuKpYkwqEYnkHu99GM57yL9IVORGwA7alMJ3f6/mzAz+8foHx6aPZXjqCbvYo9qoKEtjexv
Go+aSUJI2sXo6nadKejYyxCXKPpxevh+PkLV9x2u5PMTNwnjJ9EkDvB6WA6FV3WQm2pzV+ZuG8Hn
jqea309pPrcI4P4moyYc7m9HT7A9DUQ44NxKLsUtenx9nsH2WXfxv+T/HsjcEO2a3YWp0fnGdGaK
JF3bic5XsarsmOu5PO6tlrqxFSy0Uo0b3hyEXSUvqMpTTIENJUZEysf4HXwV/HlbwEZ3/21+ikDs
8odr0Y/WUeRdCqXUGpEoyIhkly22NciTQ01JL3BM1YPu+ZmPVXGi6tN3M4iSCjfeF+aL84mp3l06
oHQGbZ09A8+INB6uKyz6PjxXSfGfGBMPxwwXQPnm0VEjHTp90cOh1EPICM/4wmOicr7QUqx7rqBX
M5eS5IZruHqd1StwQ2fAlJrcpA2UVPiGikoQwurcW5wO7jhXmBtC21GPSeScL53veqELCA+hbWG/
4oQR9cP3gx/OvTEEgeV0sJs+LWocRQgvn0C1Gg9JR3dJvmzEfMlYOEZy5AWqAXAdBXQ4RffBvMTc
wDSZEqMQeAIo6JX05xxNWurhrRgOCmEFwkQ0x/0FvXCnkneJdKcvjcQ37bEMLUPyIhJtUuQqd+dp
swkpUIJ2TYY3MaRwuTwKzaU2J62XMwzZ0oUL/tF7ceJcYfxYjD8I/fPoXwPshBAHxt9VZ5VbOTvH
sy3OwHqSsi2XKNM8lrXgPWf0H8vtxs8E3DwT9yHBHlSree6AjVsZlQkYQJb6YDDO2lyPihNiH1OU
olc4rsDTVDr9vGFevK7Z3/r3xGV0mMqNGjURrjTt7PMbBgBl59qzr9E45CrV5mR3cC126503vWbU
1AOMZWenitr9a0ssgTVuqzdF+7mPBfsxNz2AbuGrzZa/vxBLUrheCRAEnGKeHPw3wRA6R/jI1sZh
rUTT80DUKpHsnea6MMHH7Vhax6e6CfDMerDp5fmipBUQ+OLgIHw5Fpg3w/+fwyasyRxmWYI6NfSO
abvKuDTzMzcELs1VLIxAh63ehFen/cvIZ1Z9uJYOUETnfd1XhI1d1nQ/WPaHug9DdvjAxqpHKcWQ
PSIxlFSrMsksgMM23mEf1LH2YNM9nIF7ixzcWYIASbkmK3hk4puhHt8U1jlDwnTuKtmYMmoqFPjD
TbRZ0UOhEtZvoub/dUhbge2wecmUup1rb9nKcuPcccQK/1aEOwA3mUKAxO9Fd7RyRx5CQLt2rMnP
9TTfbpC2opi2jC7aeGtHzPI5saRIBs0TOitM2soGV4hmSwowglnlvhdXgHauoM7aDqQiyROYLEEP
SM427r58thdAwUmINEHZKTnCpuO3hoXcyoe04ChuApG8UZuiqhVuRMvoY4nBg71Gie7DgVvJjgpV
e6E4HG8V1j9Oxfjodwj/pIYYPe1o6mYDn2SbgiDb89jmkLI3KBUV+deeteUYzkrZk5xjiA20uOKi
wLKAsykEKu/ZlsGWZfhWLiKCHi/1jkRR73yve5Z3wpphHskLYYzDRddN2dt7RefSwtzNUqisU2CY
gbt40vJ/Kc6zGzDoiSMCjIcHMITXtM/Xzwxo0TIOTjt3RWGY2iRWKXB1i/tjbQzgLJ8i3ingrZMZ
QgjmEeqqlryQLo7m3qzGcFK6Bfnls9P2p4Kge5UFIt7bvYhoA9tI6lBQBKY+VQxjKBZOcz2beGiT
izlbLXo+F5k71YICh2WIy31fSZ8DPPOyL7NH5NWuvvLEBlL1CjAypWZaoMkuw19RVWHRccPSRRTE
mcmiU+0RUQNENEuuDQuh5I9i5ZFWWmD5eH+a4nBmrOAbbEhklwQJZkhR9bbSGqmBYX4XvpezvwRm
sDvt+KDPBcCF5pwypR3vw5H1HvW4VrqCy9Cqf/b3JWy3yq2mIWAD5VN01MwvhHc33CKjE+BfzXhT
vr18dfzt5aqNFL7FlsyqFuLb+UO0PF8ML4sN6gDMbCRTS+GYjUD+7VdT2n9fxE7pXHkNojrkh44f
x6yMzQmPs8g7U6E3Nfc9us6qdT541k6fAMzdybtDSQKYS64ZUETULqzpjbanv5VI7bWIsBIFK6/H
Y4Q/gCKQF4njr2aquY2irPVAcxW0F4PvPsvhJYFUctgOJ+C2DvOi8e2MnN3uORmVpeFfp2JgWIrh
r3vol7nugCU7bqM9SVF/VKJZ8ms/jfaD7zd5G4k65esPYesZPyCExBiotNY2GXQ6d3xy5QDyNn7l
05vJ4HzTebH0n6euQ4N2JS9w4ztOXfT5D9jQ1dgmCZ9tdLVtuocxwxiyIIcI3gOwh9GFRTVYwtFu
WgJHEk2znPV6EbzKTwDLoxfort5suirTNdQ3c/ZcRKxj5lZ4xPiBqedoXXCwuQNvhXolIkDg9r8l
oXwhoKLjDvqhXh9Q1dzlUZMiee3Rq0AyR5lzwx1PWhm5amsW8gdb9Z+ABe8guttnzjG5ELvCjdA9
05ubrlwssqCFMH9P/glkP1JiwZSsI8H0oOj0JlzZh+xwjdb6ZL9r/IOns72uqttSe3yt4+PAe04q
o5F3ngEkY/ifh61FJCzKzhdJFoHiU+zx3eqzNeDpFkCs2nN1QXPYIlGjoU7XhddQK1Su49uj6bph
u8+HzAIGcMrlMpHryQLoCkfJW39QkFS2gdLGXw+0zqbfFMZm8YtXTbTXTTe6pv84fxWcuyJ4qOi9
Y0C6rw9M948A3bDpBk3bzkc1sorjympvNtiTIa55zIA1/ksQMR/r+Y169Wfa8afPYizWRq5r1ADD
ZPcC50sDO8AilAi48O+bs9qVXPKIZjzJseZSQnR3eYaVFADSALxu8Lp/sN2lc7NPgJFSmUFXJ5Qb
fWZAU6znqFwkHtA9iFiiZpRuHEgE+GjusgJJ0wLZSD0Awusf2kF80QFIWbJZGZ7Z2Q/Xo6rzJ8Nb
wwr1kZCrdNlva2v50IHsPZQpC6M2NZ/PbWOW2PbV9ZjlrJGb4ea9HClpgHw5WJ9WiqEoCDBjfkiN
jDIQZ+9uZgO8o9hDddMt47EUQ0uyrazd4ZKIp/fa2YDEq0pXBXZb4b0txC+M8yHZY086hdkIDeb7
IqDCM3x82nwrMMx59L8y8E4z6KxM03ubpOkfY8VR8kLsean1vC/1vP5nww2OVzsCN1iNbEJkMG3K
u9Cq5j1abp2caIqzrsTyuS1/dZik6xQE7HNkag9vL/rGGuSrBpEzSxZGuWGGrJ1WxZ349HoHNYXn
MLxLM/4Ya4NAKqH6LhDXw5jFFLn6vplnE/A4BloFSEiN7JrJHFcBtP4SZwAlnUtYU0KdpjFqolFn
zlrOPQa2mQUX0pVKJeGUVjoaKhMdvJX8e8v5SdjIfuQEXNRSeGto3T5PT1f8/2VG6D0K7ytws7a1
7CCbb6fhLKIW3l5t/4MTMJ2ohdGt6Z837B8yFTMvfPfk57XBkOGxlgTG+zvSi6zCPEl6HvOz6Jgr
OaLplKpBEsVNzsRgooWhnhlLF070SnJHlXurfShbud8VOFyW+tn5Xl0PhRVyB44RP2Hb6PBIP59X
RsXCq2Pqq0Wk/QljTN6+eHLvcigEzPZt690uDzdg0kA0NLv4bMwMXdymMdYG7KSBlf8konJxfO1j
7WCQDesfGV+1FkMIy2GKxl4hyQTdAW5AG64tV58S6KF9Gs8FdbcL3TmTUXRkswbVh7Ixj3OEnlYI
lSqHETACXEU0YCIpiCzmLqzpi+INM9xVuyU03jkO8BKysnLVOwRFglDe/VQ1keDHKlZ2giUu05MU
F6wqOnofnPBflpd4gcMtACpF0YozunXRW1IarnAGR/dSg4tLlUBcKKz9jzLIzm96wKtzTduhDsxp
OUOyEwNGZ/oBpgypojbUEvjuf3PQZPX9oV8jXA3yfVTvWYTUKGYd3WKFXNND9q/RCXEKJ7croZdL
qiAiRGGFTvemUCnntrAGF6u0aOCCqE2X+mxdcyJsRhR7REnKGZ5SUFNIQd5PXnecSS4++OBiKUQx
DEdA/0slsvTaH25Ct9EIK5kz3jhfKYxEQb1sU8rTWW2TrxU4nE4klaPIA3tXPDV4rjMWQvoBUoaq
L353lT3XtbndmpXA8r4ZQ13A217xOZ7bgnPAQAh1yvgUMQKHODoMi2fxHXCWggLlY5T9v6+gRYXZ
vxkN5GWA60HrsoyzyVvjI6PPI04tNBK766yr0yAHrYNNR0r1dV5F4+4Bmjqc3T4IXt+bjzsnp0pG
0HO5yZANviI/mhjY+pI+LHP5YiNwbOyqm/HCk+3sintXvGZ8wm897po+XFgZNYp9FnIs0OuCQsdJ
8MhxFsi6m4eshJy7KGK5v6sPV63oosg8OqqJxS9DPk4Q8jJHORT7Ds4bGeLOP+khrHE0c8+TIT9h
oJ56IP7V+s9oX6KhSSEfvb3zn6+Ju/31u/NUC5rmp6F47wOmPmBIxbpuQV5cMnhtXSMBObFaUOUv
Bv8JyyMXBArZ/JRkMWMqMK8uikxwLm7ISkeUi02bjRrlLtLyPgbJ1bLHywqBKfBaUKCDt/UGg218
xXcLWXRxyP8yC+He/5hVeAhcEd07w5vxmD3LGiExDDuSgCCVMfvw0r5y7PvZ2/g/D4iWBWRe7EHH
Uc2CBsq5p0v3C+tS6xMNWjoS5OlfscMBAqiZsSYpCsoe52tLal/1I0chtDvjOkQRIMW0HW5//Trf
z3L2EAO24h7l0diyg4OiuNS5RlIete8NaJLPuSObu+vQ+VDr9hZ+4eAn6P3uy3CXX/HNDnU9jdq4
lneB0qPKhbGUHRKjWOK6x8F+Ag8+4YEVx2wdeGEVuB46A/5zN8yxFdCukxVaaIVI54rSIIa5EI9d
fmAdupIdNEwKf16r9UA88yq3zVxsn2fw8I2aMfTwZFyYDumGFOvVCHzoe1wCapTjx/0aG2MGr1Ts
trhBmrmlk+m2+Mv4m4Lm+geGWVFd0ZZE3X+zc0e6GswvcGu6mRT/O97rdbw+2XvLleRli5/82hmP
+M588QhWRsIrUZZfpBg803PCiDiL9xV52NkUYMhtkOH71o87yKi7GazQXMth3gSP35lwsqzpatJc
9ayMHvXBv2uSui371UkKHBtqsjuGhgo8ruk5EKyAlTTOqQ4nh9ZkZKa5ZHx/6O1qiWklEJJuX9eU
sMzD/xJB4EjV/vjfxfBelwBsl1bIWsqBxi+Ji1UFunc79cEUb5gXpAcIaEYy0TqbmYCQUPH6a81A
J8ufGWYyW5la9C0CzhM1Xn7Uc/2SNd/zFHq2BkXYhAT7ZY/k7PoFcs4WIVWrzkIFP8Xym7JyT88K
D/1o8c8TAN9cYUis3kGMoLRxMDQF41mCqUvb9iLl+n83Kai1hhEU6BMSV35pDk8VnO/05Mir2H1/
D0HCxEnkQO23PIQH+GGLTUgYnh4rrZs3lkivHcEd576BvX86glXVRrqn10ZVybGwQUzsa8aIbxPX
PVMXoR6AkbR6iMHhpqJ9kQnroqoNmfZiQwsKWRX/KOh9j+/l46QmJR/b17SN1cCIvIQssU5w6RSK
ChiAbF1w76uGSeEVL7d7WQSa6YxpbXlgl5OePo5MFFgA1oahQxYL9WwZgrvedHeF+e+XeMIDKcu+
arj85MCPehGg61wFd1j7CnTkncIc4rzF/YEEyO3vC1OofdH7qV6V6iv/B1Vb2kRF8bV8ZXGvzeCV
jl+V7UR8jXwpDae76u/Nj44DeWM61bU/GgCzsZryTqLFQaMtsWjQ31kUsD6Kz9AyDzmE5fE9LwSS
GTpzJpITCeQESEJ06wenlxk3nQ56FGoBKy9PlDUZMwT5cWfIGccqGJXiHf+ZwEzCZNm4jTQPtAt1
T+Aj69PXp0xFclIhoG1yTYFkzqT0htoJb1MXyUTihweZdLuXTyvj4UCwIZDdqOjjWtPmTM4KJ1Gx
wyQK2RdK8LVa45UkqKXLxwhEIeGubeIKrWsQY9HYwGNCbS5ifDPHXiM2NweH8krdfVOGkplezT3h
d8htP4ojpHznRMmGEQQaa+1S2I1x79bAlH4hi9qKQx46Ac8t9RMdK6gRdyb9I1wLzE708F1j3shJ
2xP0G/gdARSJlooQBpRjORbBtk7xzKHkRdIQ7UKDUntTBBlq0/wUTxV8g+2EjjeWsmIX1xF6Kr+W
h6P9Eq5A2cD0Suz5NwG/LWxvpnr1cZoW0l5xzPL1PE1D8KT5RE8hcBKFJGfXbapwqWAT4veBQYIR
/QBEZRvaM0qzhtP795F/eD//q6/k/gK+7/bhGjGuTDeLfnX+zX0nyguAqgBK1tQMD29qOozlXUuD
HPCdjbH7WEawIhdt5Rdi5dkzRRnnkj/eQTu7wJH1QoEnjMLYGZeFGAVvH76+8Ram7a4OekMYXTx9
qtonXTyiKfwqZBeMy1BYaRSYN1ArNNPi2LgHx6gcvUIgE0LZVabn4o/bGbPCTompHMeohZ7ECumL
h0lZUthDBgi8x9ZGX332npu2ziZZgv2xw4GOmLsCo4bNLGsoQSlMEi8CXS6PryWs5+mjLOoqimUB
2+fyjQKAQ1H9VJ+4+okWuAhRcjIXoKFdFd365ImAwjIEb1zMPyS4goiXpQUYeN1e6OhLEY1lLVQP
EyzilXwJPsKO+HkME4OXx2DGwfBccdnUW/RHUmVrSd1afVXEdJhB9cOrZ2yPZCPr7h9z5dqGYxeb
SbGMEJBvvw/qHWESqV1Ff4ocJ3J00yuAs17OqzKFlYkjNtkNgpWD5vk8faIjjyeOEb3nW6jkf/t8
A6w504wNMXgx4+YQ9Pxj97w8PEsI5EYkAX1QTYXG9jIs7CLvkvRJ8yooVH0i8ILaMu/azYYBoN5X
jmGskeuyVeC9WgCeBj7T3BgPcti19BtKbc5oJ4kKudn/tIeUSi20fgW8H37tJgOMS5bDsExaLpad
zwEHQxTfcm/1W5nLDw5bvIFoDzUew/2uk5cgRWNP6BAtuMruXBy48XuWHXjMmiPkYBjhKCg3M1E+
h1GPigg/KgpH/MqWogG2hR2utazj78Rirs4vSOmkhpf3LSoU7zFEklwWPFVQeWBq9m7cuLmcUuZF
20DkKN2wch1cYHsNVfnyPEEJ9J3EUaP2mC3iztsrtjCCpA6JbF+Ljcomr38TTkBa+FmLAvAfJP1p
IBQwGPmj/TOfQNxNmgQV/C8N4scIyes9iE7OZLWst3yuugPYIhEdT6BdAgaZSqP8CB5hHGH87Wxj
6Nh3gvN5zDnFbAWEoqV8CuwDpOPCQjNShbMI2KNTuJux6uDs8WADrrVVQ7gO+MtyyFO3xED80cLT
iX0aIDrFVDBXxyeCmyvUuxAEWsfkDSq5ki1loMBoGGHev1HWdK1V/SqYA9rlstqEN+MUpfnbs3y1
+mcfXMUaoa4hozxga4nup65o6kNyk+YCCuNsx2ShulUpp8koYgqwHvJjrENwZsv0rZNbGwcX9D9A
DsgwKLkhBdi/7HUJx1GMze4hkQ6U1W4QG3g8oY4NJc/Z8j/qeawAQdVyBszDvvhOyRotb55ZPXyp
IlqifweU47wc41WK7q9QG9MxM6BBr9PyDf4h1ot0/4lbfskH8XAFlnrFxc+UCs6rvamWzlBMrC5G
17cUWjQyPgkfuYABaDFLo2Elz4xirzMZOoTgT7zR82BAj53hUOdd7xeEbTngrn4ImyZF4TkRM88K
iNhqjhhRko8yl2JiDmHQc9SSUlhdbHDA4tuFwxXkHra0L+LEQSLnURpBNpIsS9eTJKBS8OaWzuPG
IZsQmrAzQblcFH2hdryXFUNkOvV7DxHaoaAYIyHdhGOE7jpGjRMjbAIDoXnJUKPps5BU7rcuT+MJ
IgrZWmu6g5taRcS0/O7/YbD9WIYlv/wjG137ql6pLqPyoMYmp27X0SFeVH4EYrcoUuAoFjEDLRFj
3aSKtSLhn1s95m5vyGwvmt5EJY7F0z93K1ZqKuFmZuLYrFPnvWOuNw3eA4yjtiA+RwMWvrGJjyFx
T5xg8MV321qsLyxiLA9RRbk3/hM3fpB0MgVcmwmF4yNTUS1T7ENLMdpQFKyPzojnHs85+Ccq0GBw
Iowl4ttoWD/fClkehg8K2OGx64Hh8dJ2CCvNfWrqSaW0xdj6I5qx92xZW4qXez6uqjcvHawVOmF0
oeR3W6d2rA/zhnxNm16NivOcCrV+x1iORwlPKX5lkCu+2tsgyZgqRUJRxEfbVRym96y7wNHyKFxY
NO4SX60GJbYHq6lB4Ypta6Fa2NUNbV4IYOiut14xEjzaE9m1Sl5tHeEn82XAgbAr/l4JNCtxCWQN
oyJhOtV8UXlYZr5tQEWn2UW83Jm5ko60AYV6Xkzq0566lhSy6Hs2UntA0ct8sBDwBagw0lfjXAHq
k3Ytfa/ooEpjy4PJ1Wb1QgHSeh7+xiLxVFGRbEUbyfdjN7mg4EDZmvlrTZzkeBV7WDx65N4sgFBj
VY8rrOKWSeBaEiyWFY8ytSVdhKv7ZskAzaOeUFh8ehNBOv4vSLwdippegVawa5QITnvnSIsxMwG/
U4mbg0O1sB1le6L+tHw4HlYDs2ia6fhKvJENiopvUKjXCfkCfj0chWIkspKMke7TmSykqLNduXzs
TbmUvx31b5vhIInDPylMr9fgxBsVLIQO8lMl1xEIesGtKOVnQZ6BXorqUdFaSciLoDrJbkShFFvb
5euebJqVSh9avXLUzKeUbpD6wkZf1XyihD++2SnXLSX6pq9EBCBXxqLQNF1kp5vwDrs/hCywk94c
r8+GW0iZJY8bJO2dRYxqTWTTOz5y6e7i0u2/IG9oyUQ4L/w88v/Gj8YojX7cgv7pQFKxzihxT9FZ
08nptfzCM/GaviQLAj1HSLzyfhHWqEm8Tj0wZTJ+uXb9fxRL8nhAcALumrviLYPZB/Qn2T4T67VG
Hc3MhdmrNrCcr+erZ9gJzde9l7N9DpNSF1NQ8niun2xtybXmzTCktZaNBCpXP+S61oKbdA3buhkQ
dVczJXcZsKKYZWCOesYeUK18yx2oM2RJVMyDq38WspmqnJhwh5OR7jsTyTYoqypaEHCWBAyczJGz
shQoD0fUCYVjZIO12BiyZrDgi+YcWwiSXyDe4oyrhFR3Rfiwyl3aWLjDVXbwZrcvbH8a5Eq30FFU
9cJ3vOth1TXsnus0AOBMU3l6bXB5ff1r1Bczb1Af9nKNfDQj27viY/0lra4HTo8bCv6kNGkZ3aMT
LZLvqY1jMbBpZQyr1mPKqnmO9DLond6I4+ftezl8ABzaOL3C8IrzUwkv4HtnCrFNxfjJvL2W4GBg
/ah0dqshYmLiSv5n2WkywdGl6DBg+pwn28h88bDDnLxJLsV5/Crtfw3CqrIQDzbdCw+YTv6M0H1f
V49f8qWeepFkKzur2pZMyWF56UO795TM9zKQMpXmBgDDAtGHTKycDA2fr+j6lcJ2IlFH2IBg4VUg
NmOumHDPY7ReLyMwXn/ex+h7CFjOBuOTkTeUAiBsgoRRmKoJfMdom8rLcOsv+lPaMf2dBpNRAhPd
fLtUfJBkurePT4LHxTic+bYdZYmPbHlY9Qa/of+Bg3SJfLafdns7XSdr+dc//rr2FD0e3j2P19js
1prHR2+fp3EEwzTI4LN2XJU0EgY4pBD93Tj6E/1rWxEOQg65hjUaBDgmMN8cNgo1OX8C4IGEHXwN
Cs/myuByZOkzYb0I53KNSWt+9OtXHgjxplHgX3zGh1cldQB1a2/XhneSoJeQ+ejEj0pSHSvU/pdO
oNWKDUAdaXX7Ox62tsahC64nY/1jDERY/YxwkD4KjLe0vt2BEM4hEg3ibsHJfS5iwQI8dIvXtr9w
i5pNCk8A9uttpvPjA1IXVGxDqZJgiDjMndp4E75ybrt2ayg/Yfc0M3MVV+KRDISkuJV77Bcvyusc
IK2J/sl/QRZKKmCVlkcKvrGNLxCIwV3AacPBhqv/N0UeXg/+lDqb8W5DAuJfTMbmHfIuMks+BPrh
XzUr6jpj39q8koY2Jue8pZZKXQfc1bWvz3lBn70hYpkpLOlnMPpaKoLZ2HFOF6W+WgEfvna/ASVb
Q+2zlkLJnhskFefO6Ohk5ePiLw97OYqzO+Crodo+7RCMNeKHyk7lEcgPnr7eJGPNe2XSSUFOsUT/
v+unieqjXqNh1DCuHbICOa3gZ9wGTAP+h/gjkJF7w+d/ChyMozsCYhYp3FrOXc6QJC3aKp08li66
UxzF8FrJ6YVfg4xLklG1nWpZvHh9khJbSp+cJ2dph6nxOP7/NZguWF+GqHOHzfHAGj+3eljJX4ab
AxGnlzEPQ0lBeZPM7UI1gmYqj3kRvUgs7tJDoiQh6bdw3YMhX6LEHMicq9Z4LEdYIgtlDjiJdpaL
kHH/lncwuPAASt+Ebg7+sP1et3AmQcHo9LlRjcAscR/q3FmeawzW3S24lSQt6v+40MWiOYoRp+lC
DUTw+K4TKgSEctQxrRF1z2Q6O0W+VUCKciDTRQmgcFXE0bSbyxc9ckWedqweL6WgjdMtqX7/jeFG
md8tji6RdlSuS2D2LZveVd1RIZQUMpeSWsH8NCaS3i32nKdHRhyTaKoduWerifCj7MEM2FzQNCSy
mmaLVkMxRs8Qt+ZB3W9Ta46fP7ZlqkHVw4cmI/b+IKue4H3r9ZBXYd8U5vMZDQRjM57zpyraiJ7a
G3HGKc1Qqw+PmKOKjrMSW5FfiDrOdQmjJNxI8dmqpJyqPdBgp18aU6eMInryDo6GVuENfeLGJvsw
iz577rbN0t6r7N8m2rmnae9gqCDYhPYSCBHr8r/HntK2WDEv8gHWkpHYlhGhBIS/7/EKTqvrJLCO
PqVvR/NHGgQC6OO7kItu7aN2CFxT2uAJ0revitYVy3h3AQV9jmkFZ+ZY/cV2dPdoukZTxlT9B5+L
/5GO6Cm+Zk1G2yn5sPZ2xbB0ZBGl4TbkZ6pzbbAbieKNr0HfxHelBieI6eqQvlWfL0DB3lBFl+il
fDsdKTkfZF1kxXz9rBA5qToVPvUQCy7MeQJCGyJZuQ5bhPrB0pegFP84Gt+YIy4yWdAYuqS5+B4K
aQABC03V9MuTMXafpdpG0B2TZVLJ0B7wSkA2G7Q2hGKtxf9t4+uYgXZgKYUO4R26LV7KoTYh9OUo
RNHsJkXIcZE911iTri8csgkSwLuV3FrybKS0t56GRdjUERCx+m9m3zn64+mSYzCLP62B8ciVIBmQ
1NWwk3Vce0Rrt4ziwYKzG2U5RpuxixAg2/fQspUKmBu6DswjtGNg/ythpUlXX11tMk+aBlkS6+Vs
UV98xM1WWkLjnhSAp+MEw7FsR5NwMzp7L1/upBFC0O9ti/eCfI+I/k/SkCf9CZ5GG3eydLj7EBal
2ogboW0Vt6xO/hkt0ovnAy5JmZw7KDmkL0BSpZOQmZghnZIG9ERayxb/1H92AL9i1qQpZSi7fovI
JWoJhQdyWC4hJZPt38IhVlGneJJGK1oiP7Io6z69oFLkq/i3uD8uY5cW+Di1iwM3so50zphHjY1d
fFl1da9SuzQSlJEdDAIofy2xI4UBciZN8jxVqAJGDsT0/rg3yeGsUIxcsc/B/15WwzqQxk+9dLAI
7obf0dnVWJi8cZ79NH0WOPYsPhHQ/7HixmaNJ1oQIN4lPgsQSaDexYmclnLHl/9Tq9suYLYtdi9c
5SZIXvK5UpxR0IN8cpEQcYowWb9ICCFatcwUI06Ua5KVG5we4sEricsFjPuGpdPRRA9INVMYzlRd
mjNlrhRgoYU4RVFaYF5Bf0Z4qQtbjIemTbwWe9bN9NG4uLqnPOB2bwrwmcxsMGcZwsqLkHB+G/8P
SECyVHVhVVoSRR2swfhPgKpuNRN1d2Wp9CHSUhrv/fL4PBrpZ70GjHbIWsb8yD5eWHvzZScWAyeY
98q8szEKp8rYVlZLXENUxL8x2+FT+daS3w+yQkcgzqaUmoOlTcqTIrlGghQebcHb1H653wRhTm6m
88+TqOwJgZZu3wphzNgKyzPB/zuVrS1ZLG7lGORMXvx3Xkv8WjSv7F9T472cIKAFMRwytlLf3WYc
+cxdqoDdDfwevL0vuKXTFxaLkUdLLbvW4RSAs45hy6ORFhXuVWPMJe2RV9Nu299tapMZfBZvU0JV
Q3/3J9qbOOA3zPDuRHWgppW1CoJWE/wJYx/ojNg5agnPoIQZeZGG8STTY8QWIARgoXE8PyL4BJJH
VpmSFTNaILE8ohOQLGw5cxPkvyVGy64m6YpJt9kUyXeV7urUvx8LiLKhukEzbYhicdnIpbbZKmRD
Jyf5fcWRj0GWnnhtsQF4mp6AfC1XxeTL7XfSnKXmswfi4ZZsm3V8W3EmkUhazWWRypSpql0HK0GQ
xg9LMiH53GhaJVmSVVpVTigyE6eOQ9YumSFp6vpUjAmaGi4ClQSg2YijlTnpo76341RszuL1uUv4
yuzESaADoA5XAzIgUY85nqkXA1OW2dw4Un8fZJsLWd8WzkBZSzudr8ITGgMdagYEC9Qvjp0eXzOy
6wHtJMXETOdZfBhxQllMkrP/HkV3oFW/qd/Ll3XOTcFjjAKYRwZ8dsTtdwi2MrH36MHCGziO06oK
MCjZvre2x32gw8ZCgrBPnh3M+AOMv0CZMr9jHD2hlBh6x9hQ9H28DBK5GxGfMvP82qvkp7DqpUNC
cpK/0S4J+aca2KkC1astm8Jx3geLB+dEiilEr4iuydUDU1eRUYp1M/zRBbQGsil1ba6cdePn3V3F
dCr2vBjOCTFtWtHBpLjr7eJfke9DxuKOosrd7Rh2yEnmme7Hs2PTONzdmaRwI1PmSp15YYyoQ0PJ
CmUujJ+Qrs5xSKi26S6D7JDGD/cWeNssNj3N/0YLys2ndCAT7tHPWAH7taML7Rfcgc0+/s0FL1y2
JHcetP1ygXGXRl7wtJ9bc0nUag6hqgeWXzx+4fLC4930TTRyNc9QYUi07vUvsz4yCMLyDf1+gtQM
WZNnqakaoPfEuZPDVqZWIh8EjoQt99n+kKMKEpjIpal7EYFfFK7zR5kq4+Xvt4AoretrlG/qobep
ycWjWf2rb8ivfwWjNtTMpRkjkT3183A2Vn4yb67l+AWGE9Ddnt+Kmh/Zcjqfw9RqfI5ghnl+RXzZ
hCsZ1dMb7DAWkydihCodPyVq8tAYsMORcTfBapLdoeQZGTpEf4PrQ3FWXdries+vkUyLGUjof+14
Wj6ZRE+e1y5OFEGF1bpwKoKt0duS1aOWsComA7pyagBZZBqXWfzkl6lV8trnfrUBIrTQctDaH6v0
lkQfjAgJUuXZyHUauGJL7g0ZOQ31JhFM4j+n3b0kMaygvxDTKFjUf+qoWgyIYU+BMy9V/8e+KFBN
RFIsuMm06oqpszamB1LIjjKXtTW0qFcEIZEd41DevtUO2Sjib8rGUihuztaika6EZxr8hAQ+P2Sb
+/Fv8VdFm/0oT7QkZubItumxQqXD8Gc8wIM86nUvqdGXUzH6+CPuKjlXdIT4VMviFVLh+EJWhHN4
/4GecwzhXhsa+kqvOuMh9h+WswfRBhS7zOm38KEkM2P/N3ZScJC35rXxJCrWCG9AOq4WmoUKWmMv
sGpj/0qqKSmjbZDrCrdX6QspJOMW+4prZvkMwq/3ofV6hmbUlDyDuY+bqHI0F3vBr9CKRp+23Ltj
3lCijZf4F8QiJ5wnaL8vLgQF2cuDjsJ66B2ska7j5BcgIVuHhJ6Bl0P9nFdcKYLScylCC3cNsRjz
hbyEd55fff7twCSCvxU3sCAGIKjiGkgU4LR6Q1Ne4alpRO2wz8U6eSdS4nOByA4Tkw0x3WnLm2uE
MCta5fd6+FK6tWNXEduGzVmCsK0wH+BTUOV0pAB4/qG+W2pUINyg5XRU3qYCI3IJusoOPMe6AIzq
WvHdWKtVS6+OFYQbhPkKXsm426rYmN8JiNbZpkzanZEIhS9SSvuHqMxoN4/+TwpWtY2VZ6owM2d7
0ufx7rMsipHp2mDc4kydyNqQZEQjuOq9fv4+RAF2Q1JDV80LSGo2zlq3iAUS0Ua0biuM4QP4mj+e
GQN6U2VzohS1ARLErzpjDncfPpDjoNvV1UAdy5z/IBEoXrVu/x1jTqXFwKInCmvcaWOlqKkv2X+N
d2jntxfVL04agTBx/h3bGR+v18GoKkN5PRSh2WCTSx5fLc6aqDit9TMIydVB6sdyLdQ3femwemca
eGXuRJPctNGqAQFerbY96piOVMSrOFpREKXVgxGc+oPu/4XikF3EqqGrSUKpR6oW+ez4u3LVYIZN
P3sRf7P7/r/wDqOoL+74GeTZt8UL42H1tI6voVYQMix8YzY6sJFSpEOHxhubFUw4SZod7NVdGQ36
kD4qKQDgJ9xXIMj5Sh3ydwUDFVLQ7EdPYFTXl1iZDjQ2Pk/3zjt0gN36SvLXT7qAwxifuQziEAla
LrR4ojk8cZcH4CoBlpIFd15QTctRofF3DKFbHLPPJE7PYxYhXJuLFnw0i0kxB+elPrJ0y9tV3lSJ
qK4E+YTK4sE2OMiJ4TVCd9AdM4Md6z5MzkT4VzBIbSEZqypqUVv+CxepDwShXevQA4KB2T7cRiw3
4bsagWzmMTBUJpyNbqeuUYLXX2w/Sj7ZVt9byUjGBpG5EvaxLTzR9ueNxwP7hby0hvB6xCr13dhP
8uot1aq0ciW/rvUh1URJngLs8GB4WbtXndiI899F1YKzm06mLXn5JBkaDAgch8KepkEGpP62y9wm
ND7D4PqKSdDsLOyHbc6cu7NFz4NGBatOmBC+WM0MCTTsJ7kD3mi36WyyYiaIe9Pox5LBGYKW2SZr
iivCQtvuclkN37DtHlQ2cG1gBzZPl8IqvhVMeWeYgiUjdQ2hzVTV9ZJ5KZ1bKVbxUoY6sgiaByS6
brR5fxRYN26qIMSENKaYrYHjSDjxRNi9R9AciA85L2MFrzhxkItRhG8O7D3WzW055omy5MWW0g7S
HgocgtXNc4wQf7R3bU815W0RzpfA1g+9fjoBrz77Q2eULZY2aBpS5F/ZRgQp1cFPv9cTKLQ+15Vy
Bd6X0SMe0IvwkKMLCM6dnsQWVGQJXE1FiQqcA61xSsUPQ40qLljnqzTJd7mg9iVfOOVDgFvAddwY
AqkP5++7ZlXcIwkk0e9IDbVY60ETfwSD0wYxXhY8fUXmBdVj+/mLdWDzDElkyjQYmWDx9eiBu7dx
VwD2lsGSl1YXv7zbLL4+iTte2NRy54IaBl+vcHOx5JWmLBmaNuKma4i3uGcDxojVe18mcjBJ7arG
ZbpbBvyCfc/roZ6AE/ZmJ5Adnb5aEMycihdFNYcrGPJrLnpNAla9efnuYRGsI4vyM9wl5v3nBPok
OOEDLuFPULW9XhEuDI5vUm0TDeWXYDldsM3E5Oo6QJvt7L7YzN+JTQk8fAu/Bqr3LbA5DBZj0xJZ
A3/zJP/JijQSZTgCWU7hdIuM19pgdlMEVY7O4oO6agwE4khCx4YMKeFHBC4GrPVIVEGrLpeJwOkl
8Ybo37HxaJtqBIIsBg1XanPxztsMZc++s0SA1pB48jlu4bH9RbVffaARhVIGWkLuHnoe+bXQJVB4
HQyexkjCRuHYiiJp9NH18yPi/0GaZDRPTLMDcK8clY9bBvyUXKOBrA8/E94FJzwTfJLVRchoJU0s
KLpkydjrlpMQf/KUM/vTySymUH8YnXOoXBfhMgHDZDdqq1iB9qTQmdXH3JzrAe4hbB8II2XkjE6M
mX62Vn2cEV+lu9NmOeRWf2ZNIoHarJQwYE8plawhpasfIk2SkMWMuEhZU5HvuHI6C/Ok9bxosGar
KKSmI2otrWrVwldtMF33BLnj6d7YMHb9lV+56JxxAd40daGtvOe753n5PAhgTwbfpCK75/ZigJ+0
KWBjOfF0i5SN9jmKeGImrrrVWBsmeUFVCFtQ2u69i5j9HJ9QClXAQ6Phj0omc0eZf8gDaZTyKLNn
QeDFCyMCXBkEC6c9MQxnD+DB/+X/eXb7guwY/8Sm32JukZMojjqiiAdKSs/yYB4Ssu8b9JK+qrr/
bFLJRK9bSiTs4QSiaPukqmig2UmueKKPff0BwqC2v1GYzZPC3xU6Qymbhy9f3KMN24D/hZ0zymQv
5wG8OuSxdFso/gxyeeULF62z3MTuBPREk3SwfibzDPtlRjAGb80XDQLi5iojkOEpfNus8HWixyRz
FlQt/EDmNb/P0l4O7paTHuLh1TH9ph8uCgMT48r+wN31YnTZsa9DUDkxyoBkI59Cyg5MdAmHSsl3
b0Xa7kJ7vJHi0C1qp4lBhUF4b+AOoKxM2Ob2/jOLQs8NqCeYAOGMUB358RUleXVtdykrADf59ywu
iQdyymWlMJYv8mR/yk/ib6Jf65M0aD9T3W7fhAvYuvTRl8pA9/fT2qEz+T0iHcM8qrx1MMU+bY5V
Z5IODkqXUhb+dITkxbuPDVMJCS0bW9UgjlnMQ700SYvfmmXKnc/IUqsqk9JCFBV97oSkenAbsyzE
8ZuWynvVSajWEFYhaL3XfXftsIsVxrJ/qVHBrZ3VQ3figKTP6CsgAurUiiHa5EBvLKwyXFvdHiYs
FR7CYrW3g3W656JH/5/vqE53ZTofhDc8KdZ/WpYQMkaxni/duB3927iVJYS7RjH99Ex9T6sJhUq0
DrB34lCDMtK/m5cyJNPN7+tZrl/1GBpvNINqcMiEdx4zjqlTjYzO/6zrYdYhkBm05RuiQjkppDeE
BrUclqjP7CA8NqvKuA2sCT/VQ6YVkvP+qL7IFCPdB4CRioFKYYtmrpocbx1R/pZD/dqHKcGEElZ9
6voWPGu+pZhpEq+/9cOmnvg0KvCdf0P5qgej1T4lrbkBymxWd/KJ5Ywe2Bm1P3EkNah+P59TA904
7kdNzgQEr+SOfnb3IRL+DZ56za7FIS9o4ih+V4CnRmzOPzK9Pe7BTeI3gXuJ6RLRZNqpVvDs170N
uMFC7z2vYfvMk/JehxIRovgBmevEDxfvAB9dfk5uZcyWfAlW8e0aV1FKcPFOR2Qfbn59BxyvGTqh
dFyRnbk33R1qer2Zhq3hVeswO++2Gacc6dXTsb7oPGQ9SnWyGIIiUkFvkvSx+nPIizt8M4uMS4Kz
wAfECQRT1IqqtsrciEetNM+HIap6+44A44bFzeIxzDAU0NHWECOJFJC9KOdw+XjHH+cIZEeiVsFh
kYEU2RRTKnCH9VFlXOwN6m5z6AAZG7kJgJV7gyTTTzxhE5raz62MvOuu398/utQ/oMVZTzKzl8TS
mGpcqg6nfKMAq9IY8X7E9iKK2mAhzCNwjziZ6BzRkvaFXc1RbpHv5Gq/LJ4kyr5NK30pvrD6cBPu
ASbgT9iHw4RPljOXjtEZwmK/c29dbnnVugibJ1iZ0mVY8BDSnaFbM3i+NTWvvOiPXKpVTMBFZs0y
soCfREwKHntnVVuFCAp2jpRIFDjO4am8FPCm3gOJFqGUouTjfmhNXIDnuXlj6eBU8tlGkuu+BJ6S
AZnzctMgT2R8xnNp0mQTjl+KaYhBI96Xtwj8dXBSQoHNGvFV1W+h9tcRR6hGXON9e/GcZBRYStGh
AXxTwrKOyJU4bFOJcCHxtoooAsWRFNgWNsuycjkNAA+R5mLv8Ke3rU6kQr4BYl8Gd1qiDHYZHVS8
fJBdBmcmj16Gdivn1ImnO4lPTUNSBpB/NW5iwLM5UddC5uyBB97B0TxvioX4wb2okyDLrG1Ft6zK
SMuLWqirJCaq09h8mCDI4R1U/CWqxUZ2DMgZ8D1IaIKSTORSfCJChj5M+jWsyVQCsz1+uK+oovqT
ZSK0lIX26hMPvshOLEyu4VCocWQp/+MsdUHK+PLY8fi/dlI/k3/4mEOULG778rpwj8sERiMr8vTe
T7QEKa5095VaoG+WzRNaQGzZLp6yyGJZk6xrDHfjejAgEDnnqIPYD7z8CAA0jg5fE0QRVCSrVojD
APlH4K1Yk/japm2wUTf0W/Bf4yKpYhs2upMW7KaUuS7fuhPDQxVMZNfypZL09p5es33t/heBA4+O
FtgWuq9LP6N8HYLBd1yPYVnrlhEFe1XM9qFk5DKoN8j/E1I/tou2sxlRXJaWYllIg7pV51zU+dk4
gRnFafUymKQYpOjGiqjbEDhNxkpv2WJpzItnRn1ELvEkOAkHJgV+BQpVykjROhwcU1NyuFh3VCzf
D2eQ4r5BMlWoVtFGVDoiWcKMnmy4TyzUE58fKEPVESwJD4fJ/nmiYaBWz+PCWTNYtoSCSUa4myNw
ov/X/XDKGmkdFkBJ9y+n/57YA/N9eyqbYWBoH7gd2F5p1UpnNXg8sL2BPtDO0VkZiXKZ+HhmRA29
rTb1zLFZO3HQ7qlxbnxc225MPWb/reDd7LOCs7IKoceCgUgc+aj0I5SY5N7OTF4ME+46fss2vqcH
itYyCBCmZnrfxybNJaLjdDIcW4mOm4c8vYMWHWbb6WWajLzYOsTPMfahQmV4GLLhuRlxXo0x4d34
N/gf3xBSS5y4OeBBZuDzeBHY/LXufxD0r8vZrnKJR0nctIBGG14sSeYd8ryGWHOaAXXagKxt+um2
JGWlV3YAjHoeVWrDvKFm60XUeNeFqaTcF6s9jakQ29729UXKOh19B061Ne3Slt8DzNP2/urxilCJ
hIgPMmmNMnEfyPCaaCzyu/eTxTuXIA+LlxJhcbkT8mEHatQ/a9ieKXZ1rI1ynqh78QJTZS+outL9
OlaX0JKU+X4OdzOeEMa9YqLOhvgCc/2kBNpb2kkiRN4MUxSzf/G3NKaCtHtRzCY4o+fyAOCWTjzs
I/q2A6OoKzl0y+6pT3nKT0JucK/29FvHMn7gQHS3nGAc+f/rQk+qQL28nHYYPN+7004WzV5rNjS9
douTUsN/MOKQoen356QSpOiRvcCIIU1EMn9xOlqT4ohtM+o5V05oQ9q6fqWao7npEIEY2mviVuRN
Sj8wdetjesbgJlKNlg4KvnHpkSTCh9gPmv/FJVrcYeL3+PPyFEU9Yy/3u54NTdAjhOho8YZ+RiuB
MKesB4O2b2bQ0hk4BjQ6n8fOqiGhkv3P6O8j9a5QhGy3PO9Rv8SN3Vepey+tvgge0aJCkDDXwaVT
2jd5Uasd0MoSiJHuiJIsfaz2uxqVG3uLZXK/XG/991sDmdyS0SWa1/0ilwPLuRoa9DBAH3H4w/qx
xLj8swzufUyhSmchnN4JHWPE5n+G16pIwnfjbLhqGeik3JBvkyqtFbI/VtGsIrpMGBYE52WOmfCU
RHvHeR4nzm/qSPHL+Zy8RffEK0o9rdyziU20dS9smezBC9BXwDe0c48Xd/rHV7cDI6mgj5Oh+gaU
CMfJEM/HElv1rkoE64zDLABcx8yvvp0fbiCWVtQ3QkNJ5zMtRVuaWUSezUSt1KU9vLBqhzGfRHu8
d8puY32WX2GjsbBw2VLQETKVVfZI6dc3VnGSQ5yBkh6S7NsGE+o+GaFGPa9yl+pD4suBEBRAkEp8
UCLR+HvHxvM/JpdNjGDdec7J2OSUjAN6YV98xFTkwUe3PTZzOVaHix1nFV0Sdlaph5OmBrIhtCHl
/QJCNiua8wOK50nsubvPE2AY939NmibxVqef7JjcUC4C151LzS+X0pH/JzNoNkJZ7onFtSSVR6gm
i/vooxUSIIjXJ0rGEKiKZmczgC2cdrUnV4Xj+UInd0LiJNxnFzIkG6f2C8Ob/mM+pyEwSu692SIo
A1wmUadltWwOfam2Pud097c2H/YY5n8izsw9z8gsTu6RiWPS6Mz0q4hRD2Pdb12cANsP9pakwXQa
MCGqAw38L4MGNdgKTawUX+X+jaSuItmmP3yMIcx3jQr8vIAdBdTiMA71b3yqYk7kzoTTFr2zjR3l
yj4P74jSB4Te+07xIiM+BlXR6ujcqhVnlsCSXzWdmBo9YkVwvbIuxTGvad39D+FAcYGLXnAJFdg5
Bio/FeTbvlpTZzC7YGnhqMoY9lcKNFcNyE7GK0rWiBjepNvPZyCJHGxwN+11P4dXFuH07BJo57ba
5gZ3L03WTU7R6hejubeI+e/A3G/RDd2A/uww6meQGjl6TEeoqpnFzCvc6HZGBAEbkjdmUAuyFrmt
YObvMxc2xdvYlQuFyxvS+bU/kx/ug9eZVgYU1lUoNjnPl1A8iEZ8ZtWP4oqWoyKPyOCDKB8N57rf
GAQRFuUNM11gbSqALW5WnmcTNj8QX/nJsMPGJYrhrLVfJM/UeieIuYFuQMujfstVOzDxD7nn1RPd
BfSDdio2vJa4jse5ByC8S3Ob7n/Joui7LUCZEGkbM3DMTzQL5hQIWP/zhtC5Wcdw45Fg8M/SgK86
SDHl7R0Ni2FtShF4Yib1LfuF+sFkPdn9/aUlZc0dPFb548beVoGoHpFIQYk2PDwoIR+5UyGC4STs
QB1ec38EKgUjeZEbKNs8+OR6vR2rF36bk4vHzHJJLYjl/ug+5F9A1LChY9Fh1R6fA1CVtzpZtwAR
WP6o87CEqBvQzYmlcC8S9KZBGB2oFavqa+HpLZrn9gHsEoClH/0jSoL9bX4I6/6L2JOD0hom+KNt
T/hfpOg/3MsOJmlQLkOo3YNLRFz7dAfNcC68D10deQvzYeXS/xMs2eGXkScZG4d7cDu8iHN/EVJd
ht92YSe7jdDPKMueRV+0YT2LV97vmnT6wbvPTNy+pjA8BbcwpeUtdviPSzZ1+dZFjHzxZYpJwiPk
G1klIBp4GB6Jj5URdOqZ8oQY0Bmn4Z2PdMQPxwDAyxiy0dW0REmWbEht4HRFyecxwFOeqs2SqIii
DcCb/Iy8xD/M5eBcsy+aaCPL8SJfsLFal2hBAvSMHd7ZmJO66T+MdXElBnvRARlq1DOxWK0Z+/p/
J9GOUU1KaZbc4BUM17jg94uNM/urRCiIJ1KAAk9LALlYMUMroRr/rNBfEgpAM2Fg64IAtExED0lp
bHcK1M+xXw7vuCAslfymHOKZ1TvJ/ysCiEoXUSJN5vZJtJ7/Pyc06aZ5Amn9RktpoMI34R22cyJD
XG9inHhHPwzqwx+JFhH8nsulLg6/4IiRQlmd2fQhP6QAkpJdd6vGv4Hx3O3IGyeJ7GI6XMRqKO/S
crp2Yw59lP9DhDsG9LETfxKQuLGzzU13bGqOThfjd9uxdw/SPShFqMMhg2C3um6RrB+I8jQfnESx
7SAbBnnNb2VGfr3H3V0ZTIOPFQjJ3wHoWkrLbwqBZPSkrZdks1+0lIui7C9FmJXRgQ70mskfjvPY
xjHXwWAA1JuYucWquTTqfgE04dr63j95p58Y3b+KgmYt3zDgsReatnxTF6iQqSGdjZ2cTQN5AmsI
mwzsRbmcqE3yvpNhLBwuT/nNMMvZuzdxOXmDz2vJbBEng1lIrqrRwi5NsiplhCBvktkaRX2hQpuj
VA56SzwwBC9k1as3zdLKEzdRhAtc08tb2idxr2yjijJ88zwL546zEglvhZMhZZEHjpx6js0zeDUY
SimfAWctmFxDYa62sPadV6yYwybdaLLDv1V4b0EQ4amAIR8byLOtzsq8fB01ushzL3LcDfW8VX9a
yEt4S1MCnyS+qGRusRrQ8WVnX5aIDkLsjEZ42BjmHiEgWTiBVnX8h3D/MXomeV8dS0BOPLNwg0np
YGYMLdCCXLBhiGf0VEHW326LNHf0KihTFL64KDIBktH7d+1BrbXyS2vR34je3YWVDcjKO0z8eZVm
WoCp3XbJMlsDW1GK51SxqrakgUU6l6SsPJA2gEUfMXN4XHqyU3rFP2K2fN4FK/onult6cUeM5zbU
RGJFmBTENkbL1w4Ir7LM3mjsylgGcdbxn46XJnGn1tmb/+nPQGQsnBWGkzd4yy6ECeu/KYP0WGcr
qgWuznEyypuMn4GjSHTuhUjSBn/DW6hNnlk8UyM8R8k7unJs2MfqTuUib6avDh867LjUnHoxL/wL
EA3hAz+QHY5OmP8NASh3+IS50r1vzw2GJAhr1CnksH16zIXgCm6+lQjbliE+KscLrpt1+o9sj0pw
yWgctsU0Vil3FXg4cwRVYOfrLbJ5bhHVwIqa51CNm2b4vFqKD9DVvt7X+G5pjYwhCgk5vP/+017Q
YOxAl3cDqo3+W6RgGTfPn/ZR0nd8QokYUeXEcCUc47RyFHFQOmHH0YS9QRRJQmgx9PpTRil+FCZX
I21Apw1hGi6GtK9V3mg+b23/0/x7YuBwyivGIXlsJZHyG7u0VE+eBsUUfkIQoh5LO0Bz3Wxx2rDg
u6FaTifv6kS1kg2OlivNww4uhWpkfhxgh7ZiM/pa4XGwXtDR/do5ec59YA0D0ofejHZYAeqHKIAS
sqSFXCCIHHHoTy99MPQg9YhTASn6P3ape60vRj1ZK1AX9kLPdv2vXd60b6WnUhHT6Pfhhh1Zb8Cf
YwsS0uMbb5KBGutUrIWaiVamW4Ej8vuAWaP5reFIFW9kRZLggKCDS2vkW4UlPvyQaDNhfii+dWxX
2Y5MDyjspHM+g2LQHYjdj7KMNxQ908vEtkAzQjj2iGY33+lcgBXaDtpptSzqWfH1YFZ1UETrkSpE
BXEO2vVa7QRiXT+EObYS+/5nXT8QjGDmOo6PmGw3RSUx3rKISbPG0MKZGO7VaVxtP0BWbKChlIZh
76nZZo0knzxHG/RYjBhQrOfLfZ6HtQ+uY003fIcqgwfeNjIOYOBF2EQ6AOjknQQAG/YXd6V6L0fl
IN4QHXzQ1xl29j3OSQ1esKBOe5j7ZxC0ogAnu2C8pnJmJvG8PoaURaKdx32nldbTlzQPiVcghUfo
Ki4Gd1fBI7as5hXYco2NB4+G6qdSaI3byIOQCbY7ZDbc+2vxz/0XYZYjntxNsPO3icE3PB1WbsSF
vMTuUUOkljcj5ZnnXEKKLrVr8UpE6yVCwXGieG8Qz9IY5R2OA9pav4JAHz9nLo81vBLUVqVln5tm
4FwpWmYylbs86Eadivgevs2NkzXV5wyJ6c9eUEhnsS5mCeKa/J71S7G1x/qky1CnYqMDaP5XvZJR
7Jhdm6SLw1QNjVS8m5SRtx5lyTuvTwROZgkeGRUlikRx5sX3z+kfZ+6VBoGlQtdw5Xkn8gB/SNS4
/c5oRSdb5cWiZp9uzsix9zA3bUenfu+earOn06vzUuiFgvaEpNzyoF9NJsAn9jwr+55MV5in7cIr
P4Tev+sIycAvafPxF1eysNSXZfy/uH9g/DtQwFOQUdMF6sNPiToNT5KhJPfmvQRkH30eNfsOCOud
fFHvqU+dCLIekdIpMYqmu5Gp9swm/drdlsYrON+mznd21QQ8Aqz63lWc9KTuUFBbazM1njruS0Vw
9G6hH0Sa0AaUgLq4NEjDUHS2Rn/K6k9cHLtoyuLFIrHBU4fh6BpHp8UmklJQKr+qS9J8I+/JXKIf
La7q+xQsuCHorHD+f2uCJPg7ts8MFgdApSR+7zSckfW62JEeq6LQwK1lmfKLS3W8D06bi9plQCBj
ZZswz12KwecsbhExQY+Cawy5vJT2fAHSqykDE1X7kHYwIpb6tM+SJNLiPQpTsrwSFXhB0uv5Oly1
F93AITm7hEaZdKRk6+ornB8VAaBxnHYV0pTKLlFwNZO3MUB3JxKYreWPfj6dpKK8kZzfrlxSY67v
TDsSXQS4YJqhlYNRuHuugU8w2TkNGbkz7+0BWiKRDjbZG+pCPlUhcRK2wUTNbzSUGif+HErLrO0O
swVSLdlCNd8iNVdrLPfPcOmdX9xzdDvKHm7KT4wkfhY1X75egCs8HJaW8qydJ6LXJhKkrkk5Rv2Q
++Nt+YpD3R5KWwLTEWgVk24/kOZpqscReXsopEYBok18OVC8uEPaM8bmXd/CevcJkJLD0Rx3HSyJ
aiY81sm98Li9cdJejD5F0lcP+DRhdyV3WLANA8ZEV9OmfcIHFOv1ntuXo7KL6AXVgoABKw6O6ifG
v9bFNfljK4iGOduz86CSwvt9meog3txKDjbzv637LCIgmoA7s/WX6fkyd/ce8ScFZnIkC2/MchB+
xH1t7rp/ushVRfieyVTOuKfpZJBDgxll8y5wsmW8ZoAopQS5tbW8wgin2/PPrUtCGi5AGD7aUY7t
hVBrqQ2LThPzPCVg/ap+o6ci5lF7s406/PtCQMOva6SRmRNVUHywd8EHDnvArWN1hXZAZ8asnbLO
IPXGLUbcS8NWuSovXh3zHEPRCUQl3PwJ5HDAWlnbozOeiHviV0BR50EXdWysHdTbfJ3p3+v1uR+n
ILG2NLCJZEXBnpzgHzCimn/UcrdlaWvDEaHqS40ocHvlUkVXDewLVr2+aaC6jLVvE1nUbGHqHa31
+lDUJxd2QcJQO38GTdqTtDvFXlpdHUgKMPIBQwiPE9PdgLqNwqKrtpJusjAO/57waIo9HfAR6xdo
irswEvq62F+reRPcxk9sNDDOm4CLZvDT8AFp+jq2sttQ6kM2tdPrLJ22x2lXNjvyCkVKiOzBsrzZ
e4Rbu4RGlIp0HhBT3X+yNGDR+NiLRNWuMKz0RqsixZ4sdw3Fy/UiIy/ppcj0rOzg+7XAyQVVH1zI
XqMhBj+eTCiA6OICsoTQvg3iK1UiPjklZrNsysu5e6IM8srzzZvANNhOTjVCT5ectX5DbbQ8tYVd
wGH0nV6UkNrPM3Rv+6xg/2pofiEfMd5WokDDe8EIN0L6ym80NuQxHR32hZpQJDT3OACHQVG6B99u
XPRNyz4bnYewYhwl+xgdLPkbcU6F1YcJhswpzHXDgfjqIQLy0SBF4mgfajO5Q7a6T4Zq0QD0JSio
B92gl2AVXES7y4KrtFyyvYZPlNT7TmRzHz/Vkqc5YDRGHJwkI8MFFiyGrKvB67ksPoLpyyeXyI9Z
RjGQxmUfqJwa88igLKlDTSkxXIk5xyEoqkw+K169xiiXRHfcIJnhP2XlsEI9+gT1ADouh5G1lsct
PJgxPqQ/8KxHrlCN2b74Z8nnAF8pBZEZ6FhtlJ5BEz4GwP4Fug8Nky64t+HW3uv5bgdeaLQn5vwu
YD0rA3fJO6izwjSinYGWCXO6PGvpE6V4mzt3l8VQqrK4TuaOcR4lOzwzAN2s5qsyX91Vhw8xt8+D
MsD0ro2AT4nxyqK1NxogXF/gAB7d/8m9iYsBg8zWSMsSYfj4x5GidAVutcjZ0qKYiSzxxCVQS7/v
R3gmRNWS5FSv9dkTW8WN/syPLxwOq5DgZwBQlXXwzCqFjkNJvGNvNm47uzE20gViFM8X4fUqpG6F
Muj1V3lsWOZ3LPlvl94y3ARZ7cIYhD942wq8+LtMib50lu/foDrLYdf2ZsGEaakyQMYSdYZjQX1I
qQzpJ1CXWEl+r3JR+fPC6hWEyHkhC5nlnzLdwicVJXa4mUzs7Lw2BNRmWQSuV3qhhBGuJEv03+W5
DjHRkWSxukoUfWwxVOcxXRm1NJqJ6KVjmN1CGXuLsPHrADDe1rRwyXQ2gBx455YXk6CLO3FAaspN
jmHDJVFL0N3F2wZBqkEO2muLdc4Y58CCxK/EC1Vj5KVbwkCVs5R3RG0Aa069qphEtAdjH4vgbuh9
vTW2U1MnfzdALvukZEHDpjWSQ2outgcFyWih4YMOHyp+QQIbg5V96mpmd+Njx5rLpsZYOA4b9l8X
R6n9g8eYBuRmNeREd5NWU4s0s/jg/lsFslhaaGz441N079orY0qkT8jJ0AYK36niBL+1L0UJWzS8
RTWW96gRo8z2bhTSHFXppofOwgSoUouKauzHjC2wkJxpRrm3eyll4RLwA1KXElBHDtona9NHK1aZ
34wNpEDxO7js8lmu6JaJ2uiSGZHAQXuK39Qzoct0FQcoAeW7h2ntx2viJ0N88uAjv4VQP683/A+V
vfRy2g3TBWpowJrotmB8laXfWSzz+UEgsk3A3IN3Aw/zjkjK0gi9yxrdNMqhVMCMMulxhBCtrJP9
ckrnrCadOpZQCM+NDOXJBz+S12J/NrOSa4kYdRdSFtWVhaK1zZGfzkRMPNB4jjTM1Bkrw1CXGOqN
bXatS6kiVjIeeGY2Z3/OdbZb1kDU0JlPm3OWJ2Wesl8tyPnVMeFtCbBR49GxO10jpA9NHsBP+HsZ
cFG6yIvhU1eD0u5i1+b31L3MxX13E1kYuhTPCbcy6xffMaFw/GINWOEw1opdIOkpeOF+2hsWtJfn
Exv9xeSVcF0nBo6MCozzb5pIGF9o0DtpTf/2gcQFqFDNeYvmhwMTs+X/AkqogoNm591+c/1pv3LP
0YvV6f8PyvF6N7scUqf4HiiYDo8mQkqHjhr+7bgcGq1tiQktIShb+AfsbWMaoJ1vBYKguZBQeYFm
ydBaQ2wV9v0LVssTd6yvwVTqohXRw4+cNpJ5sLitjQ9PJn/YE/x3djaWVAbOs7Uk1W5We/YjwUuC
ZK12TYBSbTJJlOJZaAwdvLKghXN+odwOnzciLAR3j8L8NQ0CTgTTCP3qRUm0s0gDcDbbuB1d6Ph1
6VPnVDL+Momfix5F8y3JvByeJ+jgaIv7k0pM7scDjfQDYjNJTJQdHx4N0Qh9btb0q18pDUMZPnGi
8zIhqUf8DW8nF/cYyueRv01YixdxKXHwu+OzPWy4dc0sQQUn4Q5TMAUPLwutB98Nqt8JvESxgJZP
R+ctXRfQSJwg7zTc/5S7Gq3hb2NZ7cAxSjGc1+F7FjmTdm299fc0V5nlbOPg9t8ellRvGmSmouyM
PV5yHpOqj1Kd41QRgXTbjYDqM0HpS5wr8q5KcIDghkeygLeQcf2n5fyLnhoRrp4z5C0ThY1IGMos
+a3o0/Dgj2XkLVee9KrNWNSzg5jJJTfDNAJoDITQ5lnubynlc3Aw97O30vY65Z2PH/ay7ANRcclK
1c2NV89Kn/naQz05usL8AL5YcwWh4RqGvkO5iqlQBNxAxsslcGTaarU9SBVU/OdERc3z+6CxnUXq
sVdH9OAjuf/cXZ2H3PQyrAgBL62403LNDGag4hNrSXrgow0JuBVlOquCrsgMo8himMHBfGfDehY3
f6YTVQaSFMTbtlSmnPkTn6ArW08SsE/K9EEgQaH3DmszI86KL9RY6BvDfNTAXrMrKhcT3w52A0TD
fmuTvjO01ZndllrpN6sA8Cy9qQR82B4MXRYlGvLx3Y/A3cIOLptFBS94UCz1VzY9u1wZEPN/FtYi
2IG46j3sH+VcF1WD5Cy1j3NNsRO98XRat/PiQNGZJDmnxrFi2z0Ly8cBjMVdiYUowbMoSaPzLHK+
vUb/OJzmJvfritsMIn8eUTtKflo6pcqa2qA3yiR5zUZFu5TiiJSUVMeOKoPdvDrrz9uvdU3KTL29
4D+h1nA6i0fkSHTV5NnppStAXL7nV26pjaBqCXKaX/VXoYmpGPu8i0o2lsh/Y4KaTFcu232Xn7kS
YKDyXHeJkoU9Dc7O5nLuH9q4deeS/rKFtXeiIlLa16yPrz06U27YVQv6koiT6TjsapVi6XAPkcMl
LsaDWKwN6m/wsqBcXBrL2EYh2Kmp0OjR2kzVnakVu3B0a1w8OdZR9ZaEcHoaEVXDsYq0dzoLrXHJ
bkmaWsQsgwut7bCyqDQWgRwH8UMWca2gxK4xT99h1damtAqC0XfLtyBIuqnLV14tTKDW1jtZHCkR
jt5Xo8Wi9JWheCOoNe5DCBwqbnn/T1E3+gNxQ++p7jVaZvm2CmYJ3iaqkWomu7MfxteGCB7ndXV5
mHCl8EC/vvhfqqJ0eyIAkIDT4Qp+ujIvBuuylUUl5u5rS5+oX89elTglYNQy8HAZWN+mlpKN9siJ
Gb6gnSNtJqlMiwgaiIcwHsLtwplz8gM/kUw2ALBR+X2M9CIsDhYfYHDsRkiYz5g6tlBcn6tTvy/O
csvK46DvmcOhiAq1iT3caeXFmPV3Vj4a3tOtTgkJ9uHnC4XINxOawC7iFMU2XgTfIBm0DI7KY08t
/JN9g7hpH3fF1E0qA9DaFm0hMourEx81Sh9AWtV8e+UryisWgtPbyxKrCo09EJ0KouaxjoqIZWV6
EwnHFQa7qHraMxKwzzdcOCIXfxgd/FgIGV7KtQRIJfo5pGeOaNPpo5IyNXBLVHqG3DNlVyjoSYKw
VTn7yizuTnhqfo6HuCyc/YLRc8ZF15mhS3gxqIMhdYLCxG48jT8T28lcQYXFx57olFVdf0nuiTTB
eZqS9fG/BFkXzMn1WglS+9BD2/WNsfOkSEHJ6X2A23cL3HjA4B2pB9lHXZ8Gveoixc+3Ri99ftej
7+D6tSEKG1pwFyJ/gOx5PZ7FZJa1psKB5sNPrfeQFx+h9h8L9xltVxGf4iodcaAJGca8IruWuSww
bBAkn0EeHzOMR/enkFO86CdRWuo30CaCCDnxUQ6yAhNAXw5uiDNFgsd6Qnbi0KcQeDifdclqH8dP
Qr12ABVgyxAHYRanzZ2FrUzAbqReJohc1R4jNFQ0l09B+CWptvvm8yolYLUmRBnyHzj9YAfdANJC
I7wCJF7ZuULF7DGxiM8Eb2OrS2v2P1t93jcwYT9cZRyBktmv8zZcFlXm6DGfeqJgIaS7NCZ4zX2n
sUFCptuxyURlNBprfBnoCilJ8TNP1Vd+2wuw2MaNhGGjLUs2UMfMFKEoYcaxMONir2fb4WrC5yxn
DWXWCOOmm3RrtjdpVlVztdS5niumgJcMyZIXNF9LMuew0Qu0rIgge6wx+RFR0y43tsLWLVb+osIQ
ChDQDzkXbVSeHo2nGqOexfAPM8aCXoRFh5XZIBAVMyHEIEG8h6K06Gkm8rb3GKl+Pu8T6jzsf0IG
9igdIhuT6k24KEPC3wQn62GKm8yUOniNWyo0KW3CVufotyiYP52QmSWqi8snutnCY/eHJ4IFEACX
kU8S8KA12tu6foaqVb8raUzaRYTceB+Q5ujJO7PkxxNKnsY6UT/xIyEif2ZJH0CRXd37DlZx4k0c
z6oRWMo2WpLJ+ybabaFLV7twhHDO18hWy27YKH72L6VRasMDZyBMzyD7LdXvKEcnkY6kLXTz3GZi
44LapEqpY3y10Wnu7N/0tFA3Aim41d8oqsnX6r1+V4lxOcQ//9xw77vQwkSPmUL8Rb0Fo8JnQAS+
I01+j41LSXHZxjenFfJIKUjxcaDhwqom98+pHZXmck2NawFnVKiTWhQeCKelpX6HxGtf1ZwDaZn5
T4rVM2QGaEMD7KFzehQwm65zfGZqNUFC4m9p4ZZ7S09jYaQgVXmdCgly9AmkVYfSG5Nx52Y4wIoR
NOebBepUaRiD1oyFf4zgk/gzRVdgB089ufeK83k6KVRahD7Asb6wv1UQYGSNd3liOjeGaYZPUdui
JfMOeHidBVnpvZ3PzMSVWiZLMyIgKzOaEbcrEo9CW7DCAVTzjE4oXcWYx3GBJTqKx5sQJ67hRnq+
o0gw0CT5Qz2bgo2QwBxXV5tEaCr2frhQn0yixqg+EBFa06IkOyQahc1YnNwMgxffnWuY4+8e3Fih
2ABOFit081bY+OD+pVKyEjNFEFyzPEhDE1ekPc6GeYFDQwNzEOjVdQhn199n3VPpjw4oLvT/J4dg
Ad9rmHnK0zYp01QXEOY5KRItAiaDvZ0AIPBt3CkWJ36kSkONe2+Yoe5EM9qDh8ho7YKY36P1eOWM
1F31wV21pEArQ4Q2QbTqp2/O7SuZ8dM3IvG/+n/0i22j6xIg9/TF7xd6uWRia2SAqV/n6eoftrc9
n46oCGCVIEN+HHXHBQcSox634vb2gSJK6elnxoxGu0dHnt1NGlFNowA64Dwts0JIcFh0nfdE/vAZ
/FTtsviqdjPtaxczljgFo9PwrRX9/B2jcVFqLAabwy+wsS3ls4NS7xJaW7VK7tKNtJyekcfoHroC
y6EvjcN4xhULL9sZ11rRIVtRY3wnMhpfgNayhdxCXg+uTheAznKge/xeYoEuMdKbpc/nwXf5cRwD
y6KBSPhy88KOiQwENnGL22uT3XXiycF7rOwdejiUSAFCPfry3gd1N4tV2xYhpSF3aiAYNui5fQWp
TEgxH+LIGKB9CC79f6AKKZe6CJRdoiu32xtNDAJkEpD/avO+sgq4xW7r5ys/ZYE+7+kPQsXn5Vn+
OG7nwCoErR4yTCEAqTizEctu3dvSQBc/A4FVbHKC4AvCpbHDWNHy/fcqL4Hk6+l3Ah4cbMNvK8+d
4Lpeg7DyX6ozI9SPs+fSr5yJgE6ysgLX/EVncDoHGQeATNG7goo/YEa96c1k+6wrmICYK54EXJIB
46QoMpbsglnw8tay/i7IuqPwc3foynHGKoM+EP+BaxjM8183QWMBSMjg7nerW4VS0p8iy4mdPS3j
MmHcSljabRgeRYZ/fBbb5LSf0x/gMo4DfLYIR6F/oe8tMOyH728UaPGEjjCdazfPmVqktMAUx5kQ
XsMtUYVk8BKJVE77xHc6PkPbtwmlsRyAaXsa5s++IWNbpYDme/dMSL7WYyOEJKmXOFZi/s0qpfhP
zSaZxlZicc5mGzIl02uYSH9V7RHOwXUuS3CX7569aEHdpBFHF6ERqCawHRCK+n03SDiSj9whV8hD
8lIAo/tsv1IuMPARFoGi5Lsn4kGoTClu3pD7BmlgiIE8ujw9/NgCl6/OeeZgI61vgKj2xE2C5NyS
eRJpCsjnHGpVl8E+Gkda6n8jL8+2a6HA8gAyqRbUYe/oupatGgplhMBn5xBTXqLSyveU60SdAO+Z
s6HO2SyY7RjB3XR0HGJNnCRZoXrio67eUbfKdMAz75RqjApvVOxK7W0RXNIPoZROHcMwleusWJdW
SMdWlrS2T3qtr2nvZFd4St3qN7ypizIJrWwFZL+AxUxt3gVDEMFWX0tHtm9+YyIe6Q+3D5jslrsP
csc7z3L8K1h+W5Ypc1jZSwFExVbxIxUXC0eKrNbiXS3eu1JzaPfRsNAVjg523BiN7QnJ2H51eVXO
QnLR6pqcVRMtEyc4EfAvipvbFxUCElOns8iLC9DIxfUFPUA867YoFOHgjr5UFYBzNiWhRrDjSqu5
QRs0nJna3kBI5+aixA19DCoqZoKjpnlxFkeUPMd392dEoI7NUurzevS9V7tENDOYBZAaSZGdis0W
b9qW90qgF41MmEs4yXgLrjz1kEhMnQBN7kLfo1MMhcZZBJckrTgODBawiwIAgo/gNN4AWe4U/+ne
qn5BvImv310AeRuTuHcQ+4N7FXPTmLIR6x6U+Qw7b9c8cDNoy83KD5tljFmfSIalwgSTpmoSTUmf
7ilTGPchyPatIztdt0PeCMbcvgta8JFeLpZjC8fmd2vAlgwqjqARJ+TSqLB1kLaaQe77oMo7KNwJ
cK/gvdteXvNiOYYWEMAZ/MUOXWkZfKnIf1VVgRQJuS9Wnn+hjFuTiNCxD2c0abS3W40WahME3YvY
72cw3P2hFzL+RCz9lcBw7l8dKY4ZIfQjxNM3gEPncaaVl1qQuX5k9n2Q/ST9RzRUcI2J5XAe6VYP
IijR5TnNFrhqbZrVaNfuG7a5EMyyDKBY1K2ew60Lo27QbPVWMFpmSIQ0wSzlszUsAiW3RasOX31O
rCJBderblpyONcB6XyPfk3YKPLlzq4EPcQQzGTnrPFTcsc96RXaOcsxf1l6Bt7wqti2/PR5gjuz/
1tLHxlo6tzSHonwVY/Jdj2S/4Sxyyeaj09lPKkRhzpuLpDhK3So/IuxUS154A2sm8Oin5WYY/WoN
h45hJ4pyUYxrDiSU7qF28GH4t5uNOFtuNotb4x3y0ILvV49GrdZW5tDdTLj5zu997DF6kYWHuhwu
hgh7/IgzbulL4W1MVG1Q1vzlu80CMjW56C9swBslpctAIOzS+aEx6BzTENhpASYX8Vnml0g4ZsV+
a/vO3Uk8KVb/Ub215ZyltTnsNA7p2p+sJi8GDs4kFDwK+/qeZtu3Q4bKpDPGhWAWz98n342sUgBC
FFl+xqkav3Ai7qIj1OX+xHLP/r2IjupEsFmn2NPHtgSBRE9VWWTdYxK+ZIBG6ialWtIN5QfNpZdH
d1CRu8PPBHpXevGQ8sf7Tk0EWK/ODr0tLckGki7bmcgOYW6MMkKHlZm78FbIXBVQekUIbdh5JeSd
KRKC64V88aDqKar/RYbFIrq1uKAJdS1mWJSkzjNBA5SyUtmJUwbS3ErONhG6ku4652rAPZD2AWrS
SIeqIj4RX7OsRTeeOoGq/LPo/McRd7NWEOb3SqBifAaLJeZcvR5NrL82Ircz93B8Bo4OktUhS+2q
ErJb+gWg/nQYydewcg63A9wdktezhynL/6irAnRBRq3AHvHdr51080dKHlbeFmno6HUpfCtR3L3h
MYLBn10xK5xFWIM+NvIbV5ruc15HAR0r9OdPzL3CiEvI89XQkfL7hOEZBmhdqA6MHl1AIggHdPsd
S9KhMadnXDf79j9/Yet5u+gzvM7NVSaUMLlY00Xa13pzO1A7k4TMZoZM3DpUWz3z3NmAEBPw518I
7DOU9I2ZrLOpFJ+b4gBfrltDWsPKQMZ7yCj8OTwKHSW3SehvwKvr1q0zdalx67HATVngk7rcVmB1
VOYh7y3w92jNjwOwYRBGJBxr33GLXz8oo46Ad0l1uRAyz8cPJSkYX5z2F7lDlStP3EQG5XDS7smS
VgpYxcm9zD5C/pBMWbIUjx9dXLmvc5B1BhOU3h6gGuX2ne03Qldd2vviOD/8LYEODAaIP++vtQhr
wKnPXHzJOR6pSbfPpxrd/0hz8gaNwx1Bq2U2VCJwnf5+rKenHxsWTppBqBTB1ItfGTqAmS6prIts
+brLzzzlYBLexyhiEz/KBczNW/7dp4qtxwyuT1C00hP+Q6L/HRxNxrNqjPyTKjP0U368sD/0Seag
O1bwOUsm5eKZ2f5qAojWh1xxFXTo1MMaqsWhOoYUJq5nV0ZetR895zuRaMpakbKgW6P/d8llb5g9
0oFoZ/mQkliQR2uvBhtD898HzCIywOj/YNECVnx23MpnX1jlAFQDzW7QofmoM7ZtDset56/JLADP
xJ2ds94hr71ngpKM9iCxuCzy/I++ToOHe25Vn4+tSqOnXcrRZhgbB1Q7Vi0/4b5p6L6WuD0ngpj1
XmaNlRb85HDCgxw+6NXCY55jtkUktw4dDvNYjffSaKmP6yXxRDZOAMEbvR7imvbu/m7tCIBQWGT/
b4rT8guVPrpG27Stnlx1uoUzHC/GWu2crePEDn+vvd96LB64MvxatpHvgPmkCSxh3Lx9NoVMK7OE
WeAVI6LNaWwwndRvT+Bsv9D7o8og00uSUFygN816Z3G5Ti0UMBSqvKLl+8Mj0KMpgQ3f0w5gccaq
rX5TuUR4nJU+KM8IzWZqqY3s8wRj0eyU47pq+4j5zUU5xhMSZvohNrKOxhfOdSMVXLrp7829rcVs
uZ1qtuqrjIjav8zKciUTKWhR+WYCE3bqcpHFPUd9wh8KBG5WW3iZqIOhD7ZprGmxdDvMfgSOs5h/
3KgT4MpVFOP3S8z8iOZJpKOnsQAQuZipLamd1eGAdc1//e7n26i93GW4ztQW6f+GrU5nnG9qvfBd
1mMTpcMbySCoNGLZKcpRmWEVphcWeizE0x1wVktj4LQuuAZdBE1rPa/j/ngXUvBRqyj02jdzo0M8
2wIBa0OUozjY4B7oYFtf7dPkv9N9wWZoOcgQ7FRtpQK+I/v77L+ba0YOi6hCyvmrbP7YTSuwJhQx
+8yO2Yv7TB2zUVrR16cEP4+zJ+f3TU1N/SCVG0Wg+SfWNNlFqItUqSY/ey5NUTmwiIL4umGVR4y8
dzCFn7ZmZ9ysoYMoqzfNMzX+FGH2GAovs5rQm1oYZH3RY+9pcPWdCPs1EHUZPRTtt2m2HcoXTBOt
y+26JOn48FUp/+3IjFiFfFlgWwjyrXZfXD5z74ymSU+ccoMvLmZpTGk+KifDcP6SSDrqwsjMo1DK
sU/CSWgbEpmjqL4OY1dyPPlWfRSN1/6tJIzMLe497dzxgR1lg9GJ7P9cxLknI6R1QNc1rWedxNZH
KInIiJQlySa83mm6ajymluo2J9IaWWEKS0drrqHWdeSjQriwYGaMrI7MaPMerqnVzb26eFssaZx5
PlMgjbr+s1N9JfFeK5shK6qi1Liy3JagDozcpS0hBOnpzhBpzFXPjUzBhFik9V0T1Ac9j6nA//xO
hRx5xi8zwtdAdISKla7E1Elg7R0ZRkE3GNgxksUVXtqfEjC/5e+T+gmXAW5PlIn//rBLNdSFSEEg
vr4+HplHhIKlNbRRDCeeUFegjiaHrZ3oIZk0r9MSqR9dZpf1nLg/Uh0YVNsCN/lfPCmVU0+6fqZE
VQ1aZNoynqE7wNqS1d+UKrPwpQx3yHrnRd5IvzvW/+MZxQLM8UWmQ1jbj/rVe6A5MAoFN8cHu5ZS
03TAx2zALGlmhkGkGadxwRJnc3zaAjV8NnYRoa1PyNiIbrs+pmb5ePKbF21gQAfCWW8tHLKfCWSY
CBVTC4Hl2jLdyHPgIb0znan2Rr+E1O8dFD6XsGs585LGcA2acp5aSxYs0Li2riW5k8eWGZ4jOd/G
ytTPnZ+m7tY8zdaZ/IbWUDtrpWDRuyVRUgidNYQZpxyKsQkC+5HBqw3nTCz7AyYJpMGt2jIsqHhH
3tzn7/mued0vFvOymRVXnd/t4p+HHGm5UAD31Q4KLzd7lAHyxtpQO73aPRIXkYndsBMZ7MUAEAjR
sUnD4krrtVgCgE8v1Q5YthTH2iXdbW3Cd6bOi30ZlLWFrg9nWhki2lw0OJj76i+Y8gqY+wgUCTON
yloea00cxjzkvXtOKNd7bXn2+iPM0zbsJUvt4ikQMXNfHnkBO9xhr3GDkolbUDmMwwEuV4STHLGp
fPzvZeO2AlnfWjqaUXlepjkFLdf6YsJNw7CsvHsOTkBA5HNRo8Yu5YpxRBNfjlfcfn1sYmH4mYnN
NpTrlakgEvHQRGpW1RfUv+LLzfQ3Tze0lanhxyQFqU3P7sR5HRAdMnGd/DUETMwOKyf7Ctj8HVrj
B45F+WTmbK0flcCZ8Bvym7Mj8wHfdAc7rwbPruZeRUZa6n2qmC7PKli/FmQbY4SlRirKOh+Iw2R+
5rt4/Tt4VaqwL23F7xBwUriIJsS8OuVnwb//ZSPwCAJN80DPQBya5Hn9IsHL+Ew36AJAljqiCupJ
Gcmh+mowBxS2o2wqygBDz338IJ1IoIN5y5tTfq55mNXBPHI1izBMJU4SkmPekZalKh9wcYBjROwj
f5W1MXRyP+IuH44vdvT6LeZDumN5lL8TqYIS8AjSkWKDlc6WbFe0pHzEdzxkTlPmGWeW+AqApEDM
xVeWpIcfHyA40eV/HQf1zbttHHE/zdtL20mqFsByjbV2V4adL23X0yrQaK4PfsE4KyWNBmZ9vYiA
iE8WceDXe2TxEQekx5Xf+my3u+povOv44MD07YpOd5ntxeaeTY4AjLxSX0dXIgmzWv+0uNPcqum9
bADBm3rvjp8+dbNCZdHHjN+UALkcEEnrn0/oOmYDOkG0dWUIBN4s3YOBDP1NeDCm51qhbrzvX8Wv
JBT+QgEFbSoUFww05WCyoYeo5wx4Jv/HOciYn1N9eh2B3VjJLfpDIU1KU5sKFQsvYZG18+eZYfEZ
OnEMufw/eZ8CADDawpd34//l4p+JHo6haVGODiS3nqcikDfsv/aez0rt1VIMwAVv1lQMBrdOTFoH
Ck9IFqkcy1vVz2yRulwD4ziQyiLu3p5lxN0oABponUeJ5k+xTxgBM3VDLKNaTGL79djXvHFn7oLu
rUcZENp6n1wBoBuKNAVXm4bE5mk51R7uXJFqdt0VCcYEirzCXddShW/0XLZUqTmW8JletCQxDpgw
zpjNnjdwSLzT0wvrNwHkeTXOtThTgXU3YEB6BPschpNv0pAN93CeAGzK2WymjXhfkiPn1fHkm7Ng
QnchStgCYs+rCGwjRx5HyQmEX1XIFA1P1/ujODCnVKYIi51pi36lvSsAw5I7DrPtVMmd5fzoKH4h
XPKmSw3ikYIlSTB6pfMlyHNGRWo8DALeulMhbBwy4dy01rPY3HX+cVh2XeCjV2aa2B0U24Q7FUmY
6iucA3QG17QszpzKJbDHcbOjGPtcvhDVJhVrZtSuuY3wPf/AEQBgCIC3Q6Zt+/ea61EkE/TIsmb2
N4ZtZhMcqiiWUb06n+UojeX3Rt6eM8D6p3gRfWEShwMdUEQ0cq41pgCc4TzP50KAm5XhlYX+NaOh
cQhhzXPHR1k4dNkLrd3trmYRJfDX0+iyElW5KWv696ocftIMkmZoA8ZHNELLDb/Ne81/Jr0Jp02x
dAErcCDDxWDfklR4TfghS1METWVWDKAWXiJsNTV2CnJm66ImULeeeVRMHvgplBTW/nFAekVgS6yj
DmRNs7JM8t8Otw7wJ/ji69Zdp/iBs9xpSykM5faJgNLJEWoaYpWbHHUJSMiTND3DisWpzXKKUe4n
ATlbWUC89GZzGK7Ctt240DYxZGESmimQ0rFjviabMK7qWf2NQO1hVQ79DQfNxgicLXyT+YayRmQh
1JMiFwJSFGyz4sZZItUuS+Qc72t5jJE9fJzYv+fg38OxzA42MsvAkd61kox+BTRJbegLi/80pNbJ
nf3bqzAVsyTyGOKNv2QKB1jOrzS/SKUtgq+7ByFGdAt7i0AE4D2TP/EaRR/nJ3LfqALRQsRSh8XC
2/ygDLdyTtS7H+r7V3pal1F3NRQ0D0y+pjyL2pVCc1gbSEZBgwhmhFHLU8PrXae8Du/96vvsvGO9
AfDh5FNesyZP+BUpsUzXGL8mco43zCyWpzhv+zytq8Wgh6QYuilmcjQ39jsCZRnjJCHEGVYCoN4V
sY65bXCfZaP+9xAKuNadwBy8IqS0hmJbJfSzwbCBPO0F0KTbnKznnHo6h5Xy3ZyqTnEoainHs0Tr
DdOmUIAW8ojnNB8tQzHonlTfNHn+5tBGoGKaHp2762ymrIOuE1YjaYz7DvqN7TIVk52uXOAebPKY
ZobNBOhqtlqO9fqFvv6b0/tQjrhPSUrfuzIfpBwQbaoFdz9AC6+S8Zm6dOkb5QQNG8KBjKTmb401
mX1gZ5inIX2+qGHSDzHxL0Hpve7mCSuyyyz+uB2z6F9Y/bPhnpvMINgxnEgz0sYZMZDhKNHUPo1e
avtJO/NpBfT6m1zO/ZM4RGW7yYKafcSQuySm/eU27CTz9SAnMXj25LXFy9DKVDlsTayx1Zq+KZK7
kUP8AJW0CQBmMfaURM1rYjllWclEgSKYry1S/yxi0Bu4dtJpQVzSlI1VqH4dpPALOUvVvNwgIIVY
6vAsYUzWHfFQ1HmuGd79mAxoWc8EMiTN/3wy2ykK1uwbsRPcqSUnLIID07N3NKcastAUIxko1pg0
u1FRSUjdetX7FMgi5Vgr6gBP6t/gKQ58EwbQxMwHU4QkNpe0V4t1b3Ie8d3GgDrir+t/w8HMvu8v
L7jwY3XLNXwMvkkh9dRsf9dA/kmPxSFQ5Os0iqaG116vmnhH8WLlNkJhSbWFR8Ij0QKj9Fc7Ruoc
6oBGo8MokC9tCuGxcy5WnMXxDhwyRmLaeIoAD75+fHpA2QIaa9sr+nYLm5qSN71TRQ5Lf51G/ugG
9qp4cM3Z6c1xssEFhCvlGYNEEJcRU6jj9E6q5+5Qfuq3JSY8jqyrRlZtegcjn0C29Zckui9UX43Z
hNRvM2dB54Lx8uSLKzKi1X8yu8XSPSlCEFCT3lOPNhTzqqt2+bMKf5vW4MlBD6sTDzzeCj2gMb1t
PzEtF8SEYMYwbG+ReL0tSHCj0Ezia/VcmlESDLl/C0QDMuC6Uj3nHySS71Btkcyu5yyKk55yrbBe
fJm8WLh5uMnHDoTQWyuFxdkWf9hG9PmGtr0SYtaxmR6PhLENo1Hj7FnJYWE7xplueNF1QuvQyhCP
qI8tZ3mkJzfoITbw1w5gYUiXkDyodogEx4HinlWhY8HSUZ6W21ya4DtjggOA5gd0JXC4saD8Hquz
DP7P15sjObzA05S4ISmAC/+orvgupLz5wkI3g9c/e/WHBvl2157Okhm99G54Lq7Kz5/sLhhDnfsw
NYmPKhLEthxDnhMiMpnkk0oTqsF+8TFJaogdVbddLTfTHLEGGzAw64+wLst3xBY5vp0q/JF3lJWB
kR981MMT9aaWjyTWgIklM1/gWLl82dwlb36CHrfWlTOqrCjNPYKEnpeDr3zAcX65wrgQGZrUekwZ
QqBiEPWIVukKtT60Ju1rWBE2tRSumyIDSU5hGpe95C8sA82G1wEN3/8noSzoNRxDBhRFMu0PMpuT
2ht8NM0Wx7HxcSr1CKr5hrl1lvFjC4bw1kN+6+8nttd0KbgMKyF1Xs8RtqJLuRm37xdXjBXvUm6Z
G4JB2LwGpuXaayLa2bun/loGxBs9ZzhWRF6T8V3K8S6NfJK+r/qFVRq+PpIEGfFSwQX2bVIbdpeI
N90XlmX5zhMf721yQPSzWpcDFgrXa4mo03U59+/RZiVLTlg921wP4zD+iahe9OxN0JSpN8JWenvz
yOZgNNZlhn1esSC/F3z+GMbMbUH3NeEfND3wLrjxd4MU+mjCdugIs+zdBzHHdchHl/zZTfX3+C+U
k+J7ayifO8FeWXbMK9vwyacbp4aL+vjZTgK/pAvFchJg/EpLe9+BQVMaJTiy5g4zgL415ONjlArs
Beu2ybpJtClihFtXim9kM4pj62nEwLXhbTqMPUcLmx7DuTheSLBQw3/tMh5y1tPHtUCmibNN2KTy
77a4e2wbNJAiUfLLu0NbxY2AigrX0RIGMnTPhwMIQt/+ul3PN6cnrfP72fCanO1ZVlKA0KIOs80a
43pl+2NtEpGGj8W4zswNiAWz4l73n/Of16ljh4fQSecW/bCUeX7Xvg74zcXP6hu6Bm879qiDHVe5
hykUjh+7fwLNnMmU5sDttMaT8BLbsgy2a+/k6ew1H104tC1+bGGdPTPgVZi7bTaS+m0HTrw007qn
jSCKfIu6smfEugNo5h2ATTyq4hqzNAtec72Q0vD3eFXG/wAmiOnFlcW73kAvcj0nXAa9zHTPHdbY
21oXcNlGY+l+qATgm7oMMN6EvvavMRq5rAjcWTXYUIPti5WSz/ZbfVFrx+tMjcuwH9Tj/onzifQM
nOevDTfk+NULfBv0es9j+hBYUP9x71GbwYHVVDCHP7HAKJztb2JrRlMknJEUdbVnZUuhXDiLWagZ
i10Q5IIBFhWh3yoYdtSEIgMzs0w/2T/Jir5gv65sBSf3taEEV4AwgZNy8/jRZJ5RDGIN48E4AVOp
UP3Or0F/2KDqVc6THj6OBHI4kEmvqK2cUBXXwrj4LDShF+unu/hTCgZR/LP0T6B+q9DDohcEVhTs
OvexdG51qstB+UN/q4V6Q8uwvZnrQbK3m2nAjF/+3bnvWfX8uS2vIqxJIFT83iCRx474QzAOm8l5
wESvLOaBL004IqMxFn+G8Xe7murYmVxFivN42BhjQoTLZ4Z96TjZHDwV5yYK+a1NU6uRKIWgo6P0
awacgF9/hqcKdpzl3WN0sQsvp+Vat5iZgVtoA8xFnojMwiERKAO8RU/XWMY7eA3rvKmKsOAqANUQ
uvJ0PUd1FwmRi3oK5OXBzpBcLmwi+AUv/XBE6es0/alnVPUK776W8ER4dU0G6S9AqpbtawbpqdXj
fuVoJ/pxy/AblmcCRJb+i0ccZaaSDV2kIgexbbxtdjK5r9Ok1IHygxJtWnu+q6NjoCkDqZ57MEEH
+Zj6VOMX6rE0WqBrxvSMls16u4hDWfDUA4zvCKp5tFO1iRSIE/hkfu4rQJ8bMT3sJl7WURh1tA1n
H8xo/PdW0z5uYzZ8Pq3Pr6jRfEH1k/zI8ZJTNpt3uomu/WZmDf7BhTVqfsA8BNBjg5y3R3iEDssb
PUpCxMYePUW3eFfwGAHQ3d09gFN9e0QlTcazgAu3IFei5CasJlLo7CqCRmiSbTeQwL01J4+U+JVg
CfA9DPABGae40zVN5GUCK+p+XUbSYme6KrNn4GmHf5toG45lZoDnAhUUuoh1oQPLlA0+VJfASFk7
hnpz4QbShvAOr1wBaNvbl3YzbL+S/zXdP+p5nbvfI8hoo8N8FKB5d84TxXAnzlk2bazqp42rvwqe
foXBAsZ35MGP1r4fjDF+WcHw9Gx1DmwDMnevn8FNkwv/uWtcivXa1B08rIkns67u55iB0cvrXjRu
TmK5huUVhwLLS77UjEOTjJo2zN+0jPcIJX5e8ziHTYlljmw3ByFdUW6SOyH60YpJvRrI8s5fPzvq
c+98ZYD+RmK7JrdpQ/MngzQZ7KqmC05exN7SCEdObtaufBmhTUNR96wFpvVXdi0Z8U6evQGvOYCt
uzxsk6aCprZx4HenJE2BZxQvNqtUTXIQODy/tO3B9+Fmfni1s4WkZc9voEkHjAFKDO6yAmr/UwL3
XOYF8ubMjjWkNuYkOyx8UMRaE1sAakvUgQ1kaTSkw8xSPsQjkIsKzVzXv6dy4NF6trPYgZQs7K13
oKM1oGtZECZu0osRcVcMaINhkbBhuYXGfRoJEMNxxKVlKg3JkULdn14M7y+7GrbgHTpj4t+FZqsJ
T36DHtkxDSwZN4m1I/+1zCa40+zuncacxOKkpW/7SqtM9iSFuchG6fODqyvonq4/OveSMA5OdVb1
IpJOd3ACHbBxQ/8kLz4YQdfsDdBUgBNqPff8ffPorFtH/F8GUs8h+ME/RrQ9kWuKqVytgNRBmFoo
JOzWJrmd9TEbpSlGtCmsC6f9aNcBmIp7TqJaz2SI+dniHHJZqzulItMTf2pQyM25wE9PLtT/ZT8u
KHMUdb0ZkQ0WF38JZKRQegawH/xuBIYa7OieY0XFNy6XJp5AdagHfSEclodlNd5lNibjzjpFgfFP
efL+U6Tb+JJMSqQhxpIBiuOpeTCOWHSzq660cuDfpGUxb7IT1JvCriYmmBCEA2ooVDqzoOAqlceb
+7cSmdYJQVyEZCDJb/DqFaFsngSiv6sL4HAEEi/VehW0t3Cyyhh7ShyXqo7rrs8BLfNG1iRnT+IV
rjnaUzqTYutvhmWnUiT4J7xEo6qsXzh7E+yr/lwpqOjheNYxy7X6zgtcZw7O1KCgNFxGGT5v/j9G
U7K9f/DKdJL1SHt699Kr3R4YujHsjhc9IsNRr3b3hpYjVyDviE5v1JiAKnJWsrMLAVHDa8MHkFIV
v044EiTG6KrLLml+8coPsImfh5BW680YMOuqLsB2T05sa8KPzlMOd1HTPQEah1M/XZvybeBw2vBC
M2JKEJb5C4I14XDc+uGhacBjTl29dIzZyFCA/o/oa6xqxnmaFoHTcnBCws+9oUwUqZq8/VawqW8+
VE4Z/pO6QqMxSEt8HQwZRxd4pPDgHTSvLYvI12R3RzobnK6THWc6OfHeKJ+U0xt2l9L+70PGMcRd
LiQvEPYgsonR8imk4LWNKdw0d4MdFMIbynsAwh8eQyrjI7fVJUEQcZvTjkIKJ49LgqAKBIUrSYVP
1ZpiBzbEv8tvTZFb3qSzYwPYg7BGrQa4DTx5u5e1KSKNT5jzhr3FP92ef7XpnC2GomXjpT25Acld
xWZduSZbWGai/VjR9y8s0d+aWm59gtlCVV8yviOkrc1I1UqqRYENwLSkBSJw2Jl5w62MHKHZ84Xa
KSBZDJLXqw5Gw0fuXs/BOc/bFK7c46VvnHmGxKmZjY8symUf1QLbqV73rWYja+nCfQabSHdbC31J
S6BUt4sRM21LLEgl7050vHOTSPK69dQbJGneok2S+VaI5abbCj6FQCy9wzK0XhY5HF1wRszIqId5
2EhBhYdMzfKRzySUUk5OoGCyCS7Q7p1/BjSQZzk4liRJ/unki3kLQ/leC32oqCTtjwMJZhuLdWHs
/U+PpOdVo0M/WSTn82gDfEmntMZR/u/h5UqQpo4eB/RbKrYlhRX4LhJYqQgI5Md73adPSXM7y7O8
gf5GdSxo1WCO9OHBEL+iDMkjCKIRmXoyYZQkZs2nccmIv6rd/nYmddv2CNI4Zdnz2JoyoQOuebQH
6UGu2sKPfh7bL2CSVFSTBgNMeLmpTdfohrd1SohJjlSxdLKrowtwGq++VFYoTR0WE5UVEkQzL5LT
OWSw93dAOQTqb+RnD35xQqMgQWYl1u0PVQZH67MS9WkOQ1k5TcXMGntUGohvIfkshRY63S34ajBG
+eBH+mV3+nPn8b5IzLmeWyRmtrRAwI22vDN6H7CfFHnonWF4IuDRCir2eGCDCdRjKEsKuqBIh8fL
InjZDNRN1Qag3RM91NmI16hqfyjlmyx/oVbYYAaToSfAfxWFQ3/EXXmCqsHeoP3bO86H6l5Gtl43
cztj5zn4yMYs4z0rRM7zxzSTEtOi1wjEFYzehaT5E4G4v9xbFd7sKpFLBzxa4OzFgnH4s7pXLaX0
xN/IgodForwofu+Ys7V5PdeFcQ8Kf3BzTCGdIRkGN7bFnrGN2pdGQy3lpBJoRRaPKgcp1/Dlbe9V
hWvq0WgO4zzIGLQwdNvlaY0iuqddUgQo0QgAsYDbCL40PvNZVo/bvsXmNCut+XwYgbs0BsgY3wkz
BhxrYLeLwWCE9SrWKjSvdaqZGdy9ytVCY4qvGM/wEKrzPB9pZ7MOr39xJ9rVWSvka4bT3Xqtw5JF
JxF0ZzULEMrW0Yk5UlOuiZceaxl8MxygqGPX8osmTGM/fiRxRa7VzT8BLGygV3WxF2/wnNS0c10w
X66Lm0em459uwuIOdcRiqE1XROzsil3lvNdB/GKTe6D9vcUpEcehyUp4RgF0UloQ/p/SsXbzymIq
dQrr3seBIIW+6sOYJB/+fpy01j2gtvXQTKy/gFGhzEAbv+nPxzZKp4qWU537gIeQ8UfK61qeKreJ
1tNgE8yC+c/ghnUKh4wxlJCcfZsLjSAkeAJD4IY916xgWIf0D1Dmv6v+arRTZkp5KF72XWi+/7vw
mrrJFLiXx4/aXfOHsoa6aP1rOtIMV8sbq5LcsSsi4eNhwWz5fZ1ftcNAhyeNSIV/Uk9kZSmyfPWV
4DCSyc1jyBssExypYQspBTsaduGOv7sabAolPH3pDI94tg95eDWYFZUyIALL9tDprExHrcZ+dokY
ZO2Yg9oHmMUf6UPh5cV828wnyHWhpKjnv8SzNEzhyiccsFdnQs8IK/4glYOwxc+HkqY7Hn4YTR6u
+zsgPUsoL3DXpr3vt6AO4cgRvn9AbAZERNH1QBxMrqTeiXZCgDfqAwdn3CiLcRIsJn1UH6SWtHy0
tv4TLvyT8FckKq0P4RhuNBCYow7p9ELvvsoc2ofNYceaWXqfTqcwtlh8RiKDgbxtp5CRZTnyRN3X
/oJJFtAEpblGEX+VT2+xAcDnHtnWlDQ80NbsWF/bfY/8X4Ap/aLOvW7Yj/I285E/h5iaXXGJJtLT
vRjiltGJZ4YetuzNpLlok5f4ir4YeQM9SvuiTNq2+eWavo7MIkQz9B3XEM7wBY/9edaVAQi5Qo53
XmeGxfO2ZdFazrB+TGzozmRz24qbs2UwY1xnSGo/UwSq9ENZ3kDLDgH5cBSXc9vGc4HAiLH9nFoh
xxbSJaMaYW9DaqsUAmGDGKiiMdJ63QWQNScizkdKUuvc+MvxzXMbZeefAUJ29CFz5xLA7dc33f5f
ojJXkZqAZKT5MQm8TeoGwnKXOoj/aI1EK2i8WP6zSz6EHxWT571xMxd91tvAn9ItzvJ4L/i1SLnz
lxIQt4OQSFksiKwsbV8gI+YRTFXO2BY7YSrj3ne76zL/4Txa4DSOH4QhOGNOOujN5RBNvB7KqJqz
WnU4r2Rs0RHNwDvfqhqU4GAywMn83tAb4w2QJqbkyBLDkX8oQ4D7QuCoxaE8NZ9xJz6Ht9ye37Uo
kI0O9EH9S53sSY2LqXgsoiDBy/cIulpKVoaAIbz/AIBsaXY1vj8lsOoLy6n8lLEev/9RQfPOJdC5
PMufLhB8iJ4+06Px1UNr3UpvpkBiMHmjMOPGebMihCwsWQH+ljsTqvgIDLTHxyHIwfoseJgkM5sB
Dvnj11s9DxW+Y6QZVWGbEA1S5yObCozY46VUBqYi7ae+tWL6ERy1bVZ4iR2HOQFS4AUzTYMi1l35
QLUqR6Yt51uPo7TovUxNWGQhj4x44WkuG2ti1eWtz2tnllpvfzgdLMfy5Ukq7Lmt5kBDen7A2xsA
QrtEaxhLiZOXr/nnyxRF5Hjfp0hQkzj7o+Y+6YfVcmVNWOeOCZmS3k5xjqMY8vigXDUJlwUvI5UX
xxZeim9IVFddbuPMC/zXoM1u3PQ9a/uX6LitQsWd/Ak9Hddia0gSLvEj2hAGpi28/fwMAvTEY+0N
Pr/r8/bsQ8/pr8d+2zsJmn2+Gson2hwvYKz407X1GCMUL/e+99C453CgASY/kKqrffmmMuA0pel7
9w/nTGAseEhF58N6F6gEVAvww8NJuUGQjfzFW/hNf0pch16JRfHc8o5hxcE6PUtmiYqLdqI58aV8
oKLXbegzol5b1Fnsn9F6lPhfo2u9rcySlWX/BfdaFWUb36EU0kWXIDE5pY+h+zcJ3sIjjT24rVA8
beVas3NtiVmZGMyqkcYmIMojOHdJOSoMkJZ4d28xk3dh3h4wU0FRM0dQUs5AS1PooaWxGT5rjXiR
iEwDKg6uuKqiuLOrLudgKVJaB9Af6an/SJaEtNQZVtuyUml15N2zbCmxTQ+Loq1RzAtfZXXkZEGf
slxprsQ8S7XfT8/qkSuWBSYN0Nu6f3CNYCyZB14V2Nu6FFHijk4FHiKGsAK6WtyGCtcQW2fOgovk
l4vkznSTZEV01ZbHzqMc4XehcJvTk7bOwid+0DYuEozlDsWrFOwwRCDyujXPRaNlGPyvffOWGlFX
URT05n0IaAyY4oHKc5F5t/JwPH+Y8Y4XtJK/Age1hvZltxEPoCCd7f1Huu26mtL5Cs25/lteU2F+
SxldFXKj944Va5lpgJocZbc/vVfo5jdH4mvcqXa0XSvIOkQOsjltg43r5oeuVEdE/w9qTNzueJbX
+D8aLyR4laNkZKsTmBuUC9n3njI4Nf3yhe8TrPCK59UJWonty4eR1oIDXvVYE2HRlEWLammtgVch
VcCuSCOnaNSf8etJ5oKyK+H+biklL4jeOHuIrTCmlVDy54ZWAWITEbWnfFaUENwxjzKkzaELRqHC
beeXUPFgbh7fBXDm7C/eKn/jMkHJ5HSoocKZCD82fsu5IqB05noUN/ZAfRE78y+JfXmkReeKhrlK
TCsorzvoggkunlffFPIc99bxLCIKMSm6k6Nxvf0BiZVky/4liRWYS9vTcnVwjvHxqBWlkhu+piRs
t1+0uCOJn5kHHyloM45GMk7tp5T6R8Q7O8hDfaKCr0IFgnt3wBXqTaYsSBBS9d4oaHyvpDCa5adS
LjcaHr5epsH3aH7oNxfJARNTEg2n7GeJOtBbZ5NQRGvls+qFz6+GInhjgL72d9OsE7xwpq7n+hDs
Bk8Zyc3/KoUTGYoK9mcxYe9CFTp56j+rs+k1urQ9YbEW0m54B3J/zLNzobGUWRSQRNdmZhV6+4Ho
ncGPJxOM5kX9RdTFOJ15kefo7bZsVjqQEoGu9U6f5ZHCkj5vBKIhnG7BTFg7rsZblFLplqsNEQ4H
Q527vY9jlcjBipvcopmry4A1/bkkPFpX1jQAaX0ZOzGh6MB9rebQTI07TCBPwt1TnKzvwF1xEV5o
WG8M+/zv+gTTOJSksu0eER18DRO8tO9ugH7yIlQb3A7whpMrOCm3CDpexv4X7528YlrpCMxNmrcI
kdRthbm+KyQeQzmsY8+BGWAadSa8KfoDjlMpVZnfH5eJrLID7lYRmpwwmb+eBh3aJ7Lgyt4kXAl2
b+7bxQ76t/JGrrvaTY+N/s8njK7Nxkq46BYa7Mk/EZCEXnADZKmkr9iIPwBYw33s5sgjE4gYvrdR
4g/CLmGcNDrKkoXYQ6/0gYAtBbH7bOdVWqBhHJkm+KmfzwkzW2crGTtrCOtxd82JjiQ1yItaqW2q
uGOMUDsbau0aih7ve/YfP6h4Y6XwRyOpReIbzi4fuoLL8FspJyWAwiUBpe1LpJKnDIpCorSdnH4L
Jizgo8uq8nya46/EqYP04A5EthU2SbxiBBsTUlKQk3dFhl33m61lC4dEhXmB8zJ5WkekffFfwuMi
NfflNpiVyvxJ9oP2ghoaQiKY8RNNwCWhM3LZ0fkdQfqDN+Y9nmdALIRCNafKSuBMqDCa9AUb3tsQ
YpTWxrrcFBAkLyA2MVZjOcEYOeuCG0JD/R8aEBSqdt3bZlAlT4qkVvuQf3/3EV1It3lh53+If9wN
dDnaHLwSAYXFsA+2OCo6bLA4x8hxAi6nTlF0A3DDIrjbqr28ZmpZNfoGFsr9mSf8dxfUACYDfoi9
pELxjUDbr0YlS1rBQGNV8kTjS++Wn2N+9O9y1CEKLNLkUHL4X6aWZilEdhukRN8J6OScf+agsQYB
S9ggzsxkTXeRG6gIWWjyvH5n82v7u25LrNK2qncb9jxi+DmADum8yLr8/OnJNGmvUzxPrDhMikva
pHTn5E1ZNck1Hy+EGhvY0eCIuI0iazPJJvviQFm8yG3cTjNOZ45IG28DMJk4oWonAzBTYcNf+Msj
IIPYh7O7mdMb0au8cCb4YQZbrz9Lv6wup/CnOqL0R4V9VFRDCyA521N17dyeCbiaU8rOsS4nbzLT
YVrHudhnbhnYTkGi55vUK8xwddL9uVB/fH88/DadDYAaFU8rpZvLiAEo7yejzL2/lD87670qvFgI
K6bLzK2M6XjxGW9g6QXDTPZMEjWtfGnXKxR/iMepJxpOcsbBLeqUeyxc1sJ5nY2vdpjD7fLJkro3
ZukRev8zHux3trGNw53lv8ER0YDWMIdZduEC5/vlV/QPKt1jY3d+251epSm7vzzKUdx6rNk/5f0t
SSn4kCtKS+s36uZiUFi2ZuTK0WqQLaBYg3Cve5J0NfuhSOdLx6g3eZ13d5tqNkF+6pABhKNFVWuJ
uyA9+nZ4BMHJlCgnhHUGQZhegpopUhPencMn5PncJiUixnwfAB80FOjFxyC41dnNHeIwAo+Rg2Wy
J22CsexOOaxEH9leDJzp7emkVWa3ixV7vHOY/g/c5TIBdQNd0h+ibgDEfbLvWJxWUIkbmJkA2Xwu
UBch943Ao27lpJKHpz2fUm/omfnq11qO156DVu+JtVMfQwC3wRbbPzyKslG84gjz0rI0GXDGWka9
QZpvKSHRrNbD6tjdWL49GhimBe/20JxEoPOaXTXhbnY9JAdYMA1BVhPWFkd2P/L8lW7pAg4UE3ID
yvrQkYGkF/4/0dSt2ut4ML+pk6JV6SFceWp78a8LHZkN8Bce0xD//vvUQGWaZpq9lyqkgZAL8xw+
pwvmIxpv55rgQeWjJvMh97XKz3MeCS7Ta4hN0rkeuryn3j4VkVOsbBG7ZlH3lPijbMhqfs0A57Ko
d8ggQJXvv3xiV8sgroeU0JJg/mb8tS+11fvSEaQC1/jpVFOzV7fYM30BTnnJ3quz9SoElMvB6An2
ZXyJhG6TxxpL2e2PDC9qyAcSsfTZGqWyDkOHsafbFlgwsXpT4fBIbptvhvnJd/2JZkFBtIU7hQ2F
G2tUTCsS2sXjcihZ/9yXge1JoFcA5rUtjVE38gKitSF3ME+d/if4BFauGWR/ltlPnQWlhVRKR2+j
7SfGl4svFyjvvmRzvn6wHYj9lmSCFI3ToqZX5IJ4GRYOxB3mZdoF7Cdg13gksmpBUDN+nwZn+k+R
ubs8p5xeriquVUa2/t05fdALQiF/YJLqxErAJd5w1zl7mqu6UUzYP17faIKw6PLC61rAza/fXQeS
3Gl9W+yhF9eTjtXjeAZLYYTV8xkNOZnk4q6NZzpLCPDpdvZ2dO82k2gyo7KZ/1dFYvzplwaZAwNT
KRcmLjgvw8F2ORSZsQFyxaba3n7Df/3UcDVzaBvLH47zzUEvEoFZ4RcSmERx1luS6Ojoc5/5Pb/T
dhc5MwBj2CNhZCdOKna3oJXyHqPqhaSgXdkLMN2sM5CQeCPvWYjaUSqHMdqIj8bdky3CyeRvmT2e
DPBRudeC1/h7n9b+uYbRXXNaEE5DPN9r8YAyUrUn7+wFzmKA+w5dZpGJ4yxgPXnprzIIIZrAnSyX
td0b1VHzCAkygwWT5B96AJdtlJ7Trrlr8TBzwdZm8mvCJedEygOIwk6RqSN/9yYBUGM63H30AQ6w
Wcd/pOyogZKQVj7wr9M5HrImUtIWh97/VdEvrjjdPbOOlem4KqbU0JcO1Qde2cq2e65qLOXFgqix
cv/MKWl6riODyGSR1gjSup0pA5xbUK+heqgC3l+oOhgOI1599ErQEGSWgWmeYY5bhhiZr1bKK/fi
l+OiZ2xLFnawiJ98dLNVLCT8qr+nvJjpTgG9e5XCYT9q53P+6w1D1IlCQ8jItqNvyG/QjfxxXf6P
ZLfcIeyS/dGuqtep6YdDsqDVgHNVkhUtNz3fAVrrNy2wji8pwuZrHDhQQg10zSi4FKgLbzAWBspl
nCQ2qG8RlbkOxts5/WklSzW1oNPk87wcAVXdSjMH2R/J3us+dp5zQRbOrhYQ0cPHCQw27Go6+769
oyeL4CDHAnkPaDJ0A3QSJN4U9LRsCZKfeJrSk+0L0TabLE7cDYozqVH8XoHFNAO4rMaSdRUDNo5D
nApzpSmakZr1v2I5+h8ENTt7aA5KNohMOtvrGRF2q6yfBsTtBzL91mDB+mM86r84kT0KxJo5YnYR
OkQGZHmn8iKCnltAk9eL3NOIrctI+ZJMaRllsTNpx9JKYdsR1xYDE7dyDerrdmzymPP7oPpdWpZw
gUus63WA7GjyLu90h8/HbY2Zq+iMRwjI9SFMfuH99P43V2oucJmkpngmE960ZfDi2kAYTLPafAhU
gAu/1Ho06nt0gpd65GpTuhNrQghuQjCQojmX+bS85s1TmyUJslEK5gjBGPywMWCqg3jxKLEr5Jzs
2C3l1CHsFyvtZ4O8xdyodPpGZK4PY7294tlZQy/RcG0KLptckf2/5HoU8VnTrUvdL6U4wtBHhlkx
l++o2AmoK9hDKv0DJtfnNgOcRanxPhOE4IUJDKtns3mvuN13dXPC97kd3Cd/qUJHIBgsjdT0yp4O
dE1dXXZaYSHoHb83pqT3LktFsEF4nI6Jaz7Zh+2rEcStpmEg7o7WCUV4ffguDlFo2nJblHGqIiTX
Lnv3eTUF+Yr+MJFytsBMZmNqR8GZF+TY8jquuWixQPhue3+34Tttiq+ZdqWBJ1cqwlETpaxElUys
Jmx9UqUmLy7kmw9s8bVfdKtZ3oX7pGvPVWAj2D9NS4B5UKfc2KJ9fmTDrd0vKRspJWIfp25VOTg1
5gJ4vHp0Nb30pdKD4D5vOx9/S48Mm+8nMM+guZiBW/PnV0lcStCUaxbz39QOV4lXyQuhAUBkvkfY
Qcs/K045iXFzffe5uyfaZMbSBuUIpE18tf7N7tMovy0isNyTWNhawt/GKX0aG//44K0ePIPIc8uY
2PibZAPv4IIThsaoiVKzWCcHjhlbDXuc76zQ/EUG3KcnXCCSXQoJ4cc/92bYQ57XYrm5Kb63cIm3
Q/tN2fr4zQMUBPSr9nrUbuXBBShLZ3b+HC2UxfP/kuUq1ntybYD5CGe6hbegofYdAvJgh2qkzOga
BZjD5u8BW/YsZlOHSmIzvQONsab/bWdpmI51aDACiyN5RfHwfCJeKxtNE2t8Vjrst0iTnnuu+zqT
9ZAgUCrMSWYpd92Y3u8xH/UIa5hu/FvvcHAWGizcAoWwdt5mvhTEvkfaaE7gn0rs8PzonmQn6VO0
m/zX0VKqEWog3CgQrzmBBrCCDqOtXJYVjmXtd0i2PH3Lwtcx3+jPNDHRJj7XZTb1vhtEC2k8WDqp
kUWVhYh4O2OI2Mz9ZmkKnRp65lQ2C8Yb/wR0upY5M/yqpB4xr5V2LSnEU/2WKHkle8CJy4QOVaPx
SBV5uX8rV+6m6NS2ib/i5DbVVyETgZwlTZP2wNXqwDvyfVi+vPAmn/n1WlJZ3ozJHZ0HUrLt5xAN
GQbNsbpLn4elBgQDthkW0o3q3d58nc6ixg38vB2DMmL13Q+tds53CUW5gPz30atFahXvSfCVuP+e
8uqjpL8QIxvl7wKbiIWvr11MPqxtaiuG9uU3ItAh77QmFelMgoDm7JotG0vDkxlzbPnWS/nUbpSy
A42vx/+eqjjUReMTRV5JZIzf5MUKhQfiYbjIw7dCgaaKLJC5ut5rhP6tO3fenWGbc0w4VoTjZtgY
o48kY4sPpUaSbizyAOE5lc9JSBw96vizKfkruPCfKNgFJuK3Md237TYh5y98NLB9n4RMhfBNznWt
QfbVkEccA2FrcyXRcVbKXdCWesWG6u+G3CNGteAX7mfaIwaK6loBl8SaYi7YsCQ5aDaKleMn/OEr
1k4C+YurgioiFPsXRLp4zOxAzA/DqFNAWVRSWYerG9lVkQtjunAQPNzCS9NeOJ+GSogrd5zNQtMF
AOdgEz3BEn3vxuArBviPYVax2TOQAWSLjhr0k8i6LFmzkk8RZ9sGd8z6U8IHAM5PWHaA9+KtMeI2
ZOgcROqNzkttZVrRrPIyLOfaunhk57NIqVbX99NLvzShQt7pmg1J/SGSzWMsCM4rktd+341QnqnS
zUNzYlB6cEydYWCtHKHf8LIsuki63/SRYQC3cVKflWBpZ24dK78E4OCsY9tLQscm5Jk1mow0myCf
0BgGX5fhWfo84VpT9Ya9FGUBdQOq02L0wCU6MN3d6tOnpTdIIXhc0cOv3gbiolhu7AGvY7nm4Lo+
d7Zb210+Y4668qxNOXuuvnSGCvt3F2yPFkRefz7U9h78WP+DkavM/UuGCjUNBhXKFgAsa+PTgqN4
OvnDs+sCDDufKamfLweYaWFH46Cek+fWywp+2naW8Ofhe2lgto3729jg0GHupB6q/JSJROagvwLn
IjDIozCuhW8ngW2lcY41l8QvrKtWm9OX24kDXZDKC+1UgUvyhndmBwj1vbtcSgprwnyrM5/Ku6Ze
WM2wje5hX4AWXHD4S7ALRH4JpT0VsBHIeONf3VkTdCRrOLyReUZKsxcc/A3M01mnoI+5aGYdbDSo
+97l218GX0fOxIEKslJZjuKBUsmXZ1NlQQtUCMbXecvgu3812Hq9jtF1qd+0K+EVyb1AMpWgYU6a
/ZUq3WwQU29D5aWa2d2YiMUO5bovGjguq3P0T0ZAX79dUUqccI0ZqQqDUFdlYdaCLpZLw9in5OPm
3w3+40pn4ghZL/GT1sqSdCjs7AaeP7KjbxFIusvJrOenOcFxUQl1p5HJ0dkACPzHcTjLa275Tgsv
g2iryWnt5j3WWYTmpfOnMzH82vxwH5GhdZkLgwZh3yBYS362Jbisf5FQyjKAIbp9/yBSA+VIrY+X
fPp3IqCq0/0JtTp7xZapdzpmWFCjyeO4QrRHWioTxdNorrFbqRsyeyGog1VqyYtmPm2M5KYdN4MT
N3UsSn7Y0/6hUaF+6LrYJFz8WyiN3y7oEH1wuani1JzJoCWJHeYO+NHzjkYikLYAYexrWlx2MFIk
1D+hAI0Mc8+6eoXavD6XHFXcKJXY580Y/GxTyYnZdNTuJi/F6Lis39xQJzLowjhdC6mZNU+Z1cLj
7V4xfbakA0Su/nsGEpYbiPrCjIXGqyFV8gCrW1Fo8hRiAAiTR7KI5nAix+sh2hPwkoqxIK5PJ9+T
VfPuAfv7/dZRFi6zdPPoDCcUKhBl02L1pjov00e3Rs6zWtwu6sl+LsIxx8zgIrA/gyl5lV6ZrlOv
0SxTYjKrTJVZbYP3NWExO8CwlFFxW91MY5s6FK9R8VMlSejLg15hW5hEpM4LXL0N8PA9BvkWC1y/
xQVxEet5STkOfnMFzd2NYLAaxKXrH4k7wWLVMniLgckWQz/uk6jYIJRc7xAaLAYrhDk9bR+L2hdk
N3WIbEVMfYuvWZxCZAMa/mvF8S6UT2J7PhHlPjgrNHfLC9FvRlU1yILIe6TIOS1g10pvoEOkoCRr
lVmGbv0WXLPLfTdiSs+nU8tbgxN6wRNdIMBN/jm+TUWQhM1ia9s02Q+ln//s0D4DkGfKwgDaMPqs
QOiuaa+E4rtuojyrtSfieNmomA6u9Ej9eABQb8i1Zt5+lmQB4t63bcL7lZfVA9eKP2gbpzWU1FOs
XmZCTJIG3+zGRk8TE6wwRKDgHkGclEeF9JZ3i4T4AJwJ4DG0mXI80gBQORPw+vbNnt76L0n+wnAg
dNDjh/MFpzuv1QjX/DytoLcA1U28Iy8+bF6BDcd5YrjwWhB1QDm79hRd2lr0No5P2TdiLIUT9tU/
jwvg2nVr2Garp7W8jsAvqugZsodxAZgqb/fjHZCtAdIt9bA2vJIsE+UNJErd5AZOsI4o47AjOQqd
1hB5twIFWuPy3qF5pORYI8fDczwJbYOMWS2y4hr98bvvEgPnSmmtg5vFvyVY/yFdoIVSl+r1OFsh
5Bb1dFONSmxL81QP0N1MOIQb4u5SpZghBavQXBsJx2A5+3QJFXzpyQlhr0qXK1U4ZMuDqFZl2GEr
Jm4iRTCQqhm2d4SxOoOVfOz3PVBazoFnFGSR49Wy/FWSqCzelW+ug65kn+F3beqqXCkjq4Gs3Cbv
EFjNT+dy71r5SET9XBkzNS09DatxRXmWmvEbF8KUkw7xBjjd2ScMew1Vc7FUDFx7wuDR/8zMFR8X
MLO9mebPQjnrcOqUIebm6Xzc9V+nWJELVhtR3pfCP1V7/3VnlMtAcf6ncFx5TIYE8ouxwQkybztp
lSUR7ldp6P6J6GSWRKF6MwziUUpOP71ry7l2oMmvp6o6ypiT7darLJQfwQn5XrWN17Gbe0F8QfH9
KXbI9c0ZD4QQtC1uZpOHvMCsL7ISd0uz0+x+1p4fHOKYE6OcUl9AMtQGOAYnmXJISRebg0w67hHr
bVQd+TAHX4PBvLFl2ZfDOjU9JMwuJGWH82cFo9uuKTalxD2qewthWRXZyjNeqdbNtum4Y2+DnNdD
OIZZczcfgHCTcKrYdKYfOMnPT1/+m7QCDjhmClvsFVHzCl/46VVEd1pdzwgJG9RxMxaDMYSZQzEk
8k4LqJvcTY8Nz9tKRWg4d+kq9Jxz6aK8Rc3/7/5jr+66gOUO0NExeYSdWm+AxOkXJDlL0T92kYhd
gee+6ji0VA+ixAGknhCknZDrA/fbcTvDPWpJv3lAhyUc15/hxT4kDZ1OQ0PB5lwtYPZLUiPyZ29H
A2XMxYk34OCRvJn/im/do5sGwc9pPlQvHt/4IdeQTvK7nHdETBfA5c3KnbzJ+yaTNYwAojFNLGWE
LxE8EHB59OhQ/+dVFIWE/Xog7xmnFu2PcKybx2JBU2KIYrUfB5K/z8PfCYZkd3VDZY6ZBvXO4VNS
j2hl6sbm9JVP1NsJrLf7Fk6A/IPOksl/Vz4+o3vOi9g+a3vLRVUJ5iV5M9qJBPriJmvuIpCAmm4A
jiJtMxooq/Zuo2yAZnQedva6jyth1sq//cMKLkuIV6JPhe7LwO6RAwVMFazl7kEmyKER5WAYFwZ/
+fGiV3fmCN7rBmrMqFoc4IdOVRRJplHGJBT6nGuGt7wMjy/E2ikQV9evQYb54P7AXccYgo4svNuX
NWCGi1CYayU5duZ6OlCll2+/96PPG8edwxaq3YxQ5pIjs0NUK8XdF17mMQg5kp51FY8OSix/JnrR
o3J1ZSaDUqvpUCDq6w0PDE6aP4TCRTr9v1Xoa+Um6BIZnt1v0ZlhnZSs4I6ZUkzHjqrtCXolrf/l
vD0llcxunkInjv765Vq/8jsllVbYD/wyNuerXHadCfYq4XDDESFGdrSCcAXKomGCvbmALIntoUMF
DLL6f2nUQao8kiv26FBMfm1dMDhZxmrZGY6ztkh173yBz0iJnwxGMz94yYdbwBr41U4n6HECoNgV
vNXCUtAofvCJ2f8oU+5Z3NK1JAOMHT1pVdNxodiJuKqM+X+jr+2wzWtq9q8h4RDf1yZ9sPhvdH4y
Jiyb0QP6qKdXc/0zeLS7y9i1qomwSf/3msQtQOtz5KedS2pDb9e3pT0HRRS5reluE+w1atu1HBoL
3CbYI1PV53KP2KCTt8bjUwkLnV1UCIeQ8vuYynQZoJJGjq8BUaWIEYbeDw+OcNzxqGdm/cAvSnE2
dKiUgFlyt4GVqdRibEX6A9OOFTsESazsIEB+IzQtXPtjC0KSo/TRQ+A/5rHNr9hRHUYXZGTG9w80
kFu0I7en3Rhl/OFlXKUoxfUKqzS83FEd5c68S4b0xxLMDpVn3gZ94xG1vF5Yes+9XoTHExYdPkxO
Iwg5z1+DPMoKtHzR5wuMSK38gpxZPisVjFcGhnVZsK/XFFM32PU47OlOtun6mpX4BDp9oV6y0Yrn
i+dJ1FxkuNfa7ovkzo3EvtiiQtXUpxc4V/k+GCpmPPKnlFI317KGo3afFJ2G82osI2VHM5SbzVlF
sCAseYjAEAw0cxjAuIVOD4guMltnK0LqFtoZ5rpyX/ZE+CjenCuaI4W5W3GmUaV4nVyAsbqwgYGb
XnKUORGiOOMQc0T7PSHoHNDMG15aiwvlbGqRBbY4QOJ30B4vKfSv5jnj/HmEkoHn8yfxhJpcBao3
Xxevm/NeemBCnXn4n/DREu3aPM3lks6ZlxcSr2RZOZ9bTqFZ86k78fGf8m4H+pdFCDdtZTpsxGhD
KchHpClKLVPBVGLfUPgdsRA8HYHV9HZQw6YgLGbp57do49iW1zHE/Rx7IPFCSL4qcPwq9pG0nzye
bpKBcGloTrelJsQM0SQGCJpGBVLOXHUz2i2QMslr9SwrIp0/doXWTTO2y+UO8qN6LJ1hUG1Ec9hv
xSoToCDucBVEWvv+9sp68iRsCFJ3ve+0EmEa6AbvDjW0u5tIEhGISphnvI87FToNdaMAWrk8zi/6
w3oH7vYJArHes6Hzp17sJ/S9rt1FdZbHLOp8MS1PK8sTV0MXz3bf+q7wRX1gB/Q1RwBw5XBPCDyR
RYAGccbCt+c91ALhJIvf6QMztnrBP0kerbdEjiAYM0L8GdD3I3PPnrrzqI6c3QgoaqSTWVTmUtXJ
l1xBSd2QXVJIR3VGNDEXB9Mgf7/VMBqHUKJ2/D3KU0g9K9ywbXl2QKHelvf5bDYSE/7rgeKqMGkM
k4PqgInwiHutN+iltj2JaUipGTa3T+RL3p7Ik3A0mWSIS0iPIosuOxbAe1+pFo5PTQfpK9NRiiG5
EmIuCrxZzDvkiaLaDWegutddLtcIC8ZVBt/2/eOcuvrxljTEpg6jg9LrWknTgKnbXGwhHfb1UI6W
Vvc0H/AatXNJSVvXLwX/5LyPNvnTi5l7QpX/uBq+5UNye5aqN3DAHc3aadae9m2hBQ2cbC2r57U7
MrKSfK7gdOgYtPfDZy+esTEJAwGNXuhUXklM1idNYEn7unx/WrRPISKwSzm58DEcglus0dqwr4TJ
T9laieF3rrNtyRoCcV9cXd/wqhs8R8TFIgsGGZiybyzuNk/vMd6Rgr0DwoKqNVGHBQmRnr88B3mG
6S1t4DaN0TaW6qwH3xDyt94s4Q2v0uLaAS3zTZCskX2zGj/hONnYtEDH4raLhU2gRAfYmowkoRGH
W6/mcPM4hMoxsQJUsiS+SGshiNSxyBPahL9VoCXPeElOTWfyUTKghXEFrJNFwyM//+BzEDWYLBA3
Sw2z8xBJ8IRtr75rOopksJmvZpe52d3DxKOg1UwtBKSY+rUPfUGuwF4W3S7QoKEVXEZVTEFLdQ1n
SuSczfBGEpVUotOjYxLs6vzJCrA6o2/6XHIKvSgyDVk716nLC/JLj5c3q7XHZH6P8LLU3Th1cZrQ
mGmmSnIVUnlzOdTBR8897GWf26nMTF18PoW/VTRgGfyy6NM165RXrZ9DlTOSjplPahbNeqUlUoDW
4O7wqTj7/lctzXidTczCx6Q3GkaidJf4nXJkgnPHpC9OFsYva+GNcFz+w3NI5VtQS9lG81LhNdad
/tK0etzCiwGZS/2V3UAbpY+uFRR5weaXQku/zPVm/81SgJovYE6+5Oo0EoCHgBybJ5EKNd9tKmb0
T+3pA5gqQ7Dg8TyAbWHW04vVAI3IzH/JWyaC0OcuQjBQwcdPY8jHkchcycyGDqQUtKw47bmRGmTG
vTd+haSf9CmQv4217jgupqB99NyzPrVUDUs5ZgXtq+awAL9fQx6OR96mqhc7uadkdIKKgAc1THBo
34mya9kZwJh9y+emBa8mb3e6idHuyCHTZ5HNCnhPGpLROCyWNWMO6L0eYPRWbi+M6s+i3YPrnSRu
DQbtkr4kBkl79LD7JhqD5tgfVNQcHfowhgif0FZcm4ap/A5C/v3MtQ9dmMWdb8wTDFcV8V2RtiDM
8C2B+BbVqkOomXfxYWDK6Q7BoKvrwhM2/bQvao8FqjG0+kIVQvQGWjCyFLwfaWtYQW4XbppZ1R8s
3HjihOpJbzU5UAJEnUryfLeTsSygFNB0xouDrgky9r2R4uYi3v1mS8sSuyk09f72iDbIcMlM84Iy
j9Z8y8vC4p+Hkchv9i5RIkyr6+xEB1C+UWjNWwRgJi95L94QFPiUenwgkMJCDBPwvGx+NuXLW8xV
eQqvY9YbJ8Yaa9Xo8jRDhGw3CP14PnL6qkoIxA/Ak9KZfDSaiBW8XkWewArZG19QREUhhVAOLATo
kS35vwM8pF9nvN2G6N+I9xoDvxY7SKOy9ZcGrk4myM82m2+cvcadaEioQ4/ImJ1diRvotQRMkc0e
talKtzjJApT7mbsgLbUZQtxpNOXPxFB5G3u3PzLuz92a8NMa0iMRTZaeUhnblwTjNEp6FSNv6lDv
ZN0mdxD84I1txfWkb9jS5ipibnQMktxFj5VJKxlVrNimQvfoSu8ahQUx+ZR6cZSifoZmADsNfHeM
FqSa02Q92aS1YyvLhR90SRo0FclrANtgmq9V/aKbA34SKIdOlq1jdq9CZMAPs4fJCRT6x9zoeMu8
lWgTVqyaumjIUWAsJGKA00XGB8nUfFhWxWK8zwYywS6rq+RbF/8lzPdBesSq0tKkyAl1GrVxWhk1
6Yel6dXooZQjH6IVL+VH0p2H14WgeCgBz1qZTNTidQv9rTg/mHjh8xXxXHzI+47z4VxI+9ag3i8J
wYs89KYTcrqY4XqRi20/ERqlo5+Ka5X++crx9JPlF/6N2HIVtjQ/Id5+zx61bWR6kOk40MK4zXE/
eRwBYU5xcPNwaJpj4X7NYXnxTRamzpAa++zJEaym1F9ACi3n1yFnVBxxe4ZW05T8sJOQonRVvQ78
BIER95NUpSFaMArF45DC2iapnhmxsdyMEdWGugwF6h6kqpQW28+x223pY5KjL6daydsot/nnE2zz
5wWInxNFQlt1uVJ4/pfp6Dnfs8Eeh0WA8BgNM029HK5CM+NIj7CSnhuh4K0RY0RRdmlzTw2wiBsv
VWHTZ9hTCj4qVT/tfN8SsFsjqGDXODC1OoAfI0Fp6xBnH6/KXXS7k+V2/gJKPDkWV/49clKOuDeI
PM/B75eX7lRFVA31rcgZXcYCw/l7j3kUhOysExvAvtf1vM4yRYrARkuYws4Kt428oZfnuP547hVB
pkXlrfytauIncEG62EUpgnEFg68bqlzE3hbDOuW7PsItY5MQJI9yAiQL2S9KJva5DdepEeVd0SRA
wxCPd4eWKQh5nGrJrjjWt9z10lWoqPymgHE+2AIKldHKbuNyX6LXUXcIbjVC9k/fj9wCUI2/Ge+C
WDhcFC7727T5CSmPrKuKMBGDOhiL9ym0chYEUNxSsM1+VQOMXzyt5PZVOT30DIaUYQE+kT4dr4PD
f6emPJTfvcZLqCiaBb6IXDZwZWjc/bvvcuR56uDukLpkRSlBtle9b4KII9KpZwooFvrW1Rr4Ut1D
Jz6Y0C9pe2f9YXgF55QqE6+4t77EuTN/rIhuUHWC8mRlSY+MnKzvJFlfoVTG6FT3KsoPdnIw9ahc
/PoL1/3z8yAR/0HGaQG2NrbLTYLsDZyZWSb/QFtoAk6ywYUJN7eBohZOnxcBMj7VWlaLlWjTEwzo
6AelNBuA+rxMEEGW9y2TckdIvKSMiJ1/8/ptoPrH0vYkro8c/iyAaHfgqzzonha1XwnIUp2QLwsv
DKNn40uUtJKHMmVPmhGVKatrRixBDbjscLV7q5yhd6Qll3T3FiZcCnfv5O1oUppMR6DoNZpTa2xp
PNZj3DHhDtkMCwM0YjHqfQEHhnR7+PhLVkotcHWedVe8tIm17Qb6snNVBXWzGjrZ+QTfbDddbfTN
mH7ly28YWaPoY2zhVEzlBchdX7gIu2mhec0XQ3hfzK7Qpc3wyLIW1IN0N+5avPEEvIMAljILuZT3
X1rkIYEo6DHCitMedSvyaVnRgXhiNPxIgKoqhsXWFdFcdTNwQZhpNh1MDwsBLOp/II68NP8IxAoY
ajKpXTXlM4dRhq27L+zBHooy7Geg5pDWb27mcnnk7Z8l6yfAtasAG2Gf8yrMJ4Txhjd4anO0NH0c
7LpbuxYatrlDH4F+YjWlv5sdK4CUcfZMjOs1xFlauMo26K8n0ufvJKY7vkSIza1HV7kzIMY9d6Uz
rXRPeejavxyE0LXStzh7YROSijl7mgXeziOvqAlTwaZ+FKktiHaXCnXAyodwm7hAvBP5CeM3fwTl
Q52H0cSfVEUqR63t7l1eJcXNhTm7TnAF2lAdXxCdA39XppCXpyfZ+ewAy8UoykSgR4pGAxkUSL+q
NWIR4w9It4Xj2v3pzA4Uw0UBvzi0Y17QC+9K1QVOHvsq5aXI6rmQ7g3wDDfBoI7umTWciIBM5mSM
C2B36Of8uePqnGynaSvW18rJFotOBa1vK7WNsItuzXWy+KxAWqJ14CESSBQnzKlaCwF5cfIxlvBs
S5d+yKFt3zTXfoD8Txridx8r/QFEMNPQGFgNLSEjF4jQxk/gHbeyUbjy9wZRSU9QYyk7KMVefTfn
nu4TcWgfGhKL3YbMDluodX7WdkObc2+tSYI4+nLUcqfm7glYz6CDddaMtvhz33pfL8JkAjPVEnya
2k/DH3bLw2qIoq7baw2N1p+EttHSmSx6uJunT47z86kEl44KldQc9EOSSqsfns5o9Sr65IGJJEFS
3MHRMbope6u2qpOnyc0b7+vB1Bzr+rBeHOjKZaQ1WABsLfzKlE7YwdBh0jqp+hq1O0IYvAheNGLQ
9V8Z4F31X8RDa8Q/1yecFpzOxgvVUj/+4IbvHQNylMQJXoWiO1voH/Ae3ss6qNah0jNHQgGKE+CO
qVD/hcH6aQOxS7HuRXRL/g3sl/ft+vmYdsq6+HFe5WzfcP1RBemqE+MLzU3QhLj9+py49tkpAyad
MW21GEMYFok5RW0DCAxz12WAzVNsffJJP0I/4yyHcziaFoYoyVJv6BiAnfrO/5uwrHSF+3H0pqj1
DDszLxKEH/oPHP89Xq1L9rZwiksQdg+XzShmMd/Ba6T1+h8pBwAxUKLxuZdRCFXoW7oXyBLM68Mh
cWYyueF9H1KzeXGKByeEjLX0y6gjzbavjevm9sw5zTt3oTrsSw/KWiSBAL0CDUNAArDkXJo7VaIs
wSQCXIFJY0vdT5WQcek3tVgir8MKMq43ucCPNd1x4DRSANiljT1BsVVbleCu9yQtEaR3Gios3Ioi
gAfn7A9fyJyZ+SZtq6rhA66/JogAQ80053mlFtMrDn5wrnaYdQEndFOOKPhAO6llWgGDY9kZ2XXx
eyBWcTTWcdEB5cUj05P5GmkcMw/rdTfLVk9uDFC67I4l2zvoaTrv/nQeWec9oB+r36EekDZOWH9K
RwUBe58LMXK73zutYpS4SASt3U7VOoee8RrIncnk6MdDU4HbIufukG4K5QSZT2eJDo8qDwMJTtMX
LNk3WbEAy50QyGbkOmkx3QdCKpJQDzQZhp3/m+Alh8bGvCXmKeDpk693yYhtKHEHe+7CzGoCQa94
WtQJP9oSeNCONwIL/Uitqo17Ohs8en+w4DWzOXPQaXLgKUB6K2MFHqxbIB8JZo6p2FHnh39X95qR
hJzZmwrv55AtS8BRIBg7FKZQtsr7ugyHPVkzz1HJNgRY4Zgv1rcJwWHRiI2xBJ80v+g4r2n//OvH
aLVS1B0WhrRAclcMYKGEXHLG3waEmtUD08CpdRyoqtdZ6Mbws0nCqihRMyd3kJbAot5DMV7vM2ic
dl88Qj4o+wIBfxkges/goS4MnuuX2wyJSABkji6ad6QRdk4/rLQj7s4HtPXOCMbZdhN6sz4GGbR/
Mf+0KcyZoUOAAYt3EMcCX7H178HgSxNAwVSFqgpsSd43GiHmbwpLY0aXhvJHp3JNLncht9Ocoelg
lQoqR6XhlZbggg2NFq1eIuxwhePbZTMhsIa+p1b5mbLkCSr0krySAbdLgoHxifUFAL0TBem461Yz
sCtLYFkJ2O9NSzl5RedoCal+RF0A0cIL55krQuixNiq2tebqfOLwu7y+GXEr57VzS/4jlLcRIRNP
gN9nvtWpbbjkSNj7d3ILnSdwomeFR4kpxmjATydPvzmVjUFINlB8EAnnt7kICB7tlUd1K3p4HqHU
qQSA1zrbKYyTxJ3w5LdgrOdggJxQpi9ksyLMnW+QN3XJ9fVGAHSnMaFexX61Ph+PHygY/0p8OH2u
OjVO4+pwEy3jiYHF1flp2AXA1xvfGHxQHgBqnU9mIoHzhFFJNdgpLWuxl1UlAk0uLZvrNorxOWAO
0mUEnqff8SFWNCPA72XIzzYlm08FAoAWTapbbSeneSKIfQvM15Y2fYU7ow/o5FVA+WvN74SduWA9
zhKqCuacFRFEIK9p2rcITCrUy0aB1dPXI0A39QzTrnBoejDC3bZwpL8iohmGgnfkzasxbrXjFwN0
f8t8UnCUepP+9EVpzudf3gwiLkkzEyfp3m1wKV5VYK3G9cJcNFEnCOsG/6LAa3uULzwr9PK9N5IE
ojjR3vSF/DljivmGwLYeYOy2ji+JSEGtfXKYwiX2ZKQxHaBl+9uXLO2UCSyAwMGAfaldUcNs7o46
fYx4+xNtzRoCY/4nyWMr1mEb82LykXW/W/GemDxubPXsg81DHJFbFSWddojh+73+QL0VZxqVZsrM
hvk+3VTOytKD0m2GW+utPrnjJpuyzPTUZIrKPsi8zVHvnU8D5qG82N3jrxMaiKaPSmbfPIBR3g9Z
DHl/mwS4F2qWhTq1ocFz3FavTKcJOVIKKtxIZBa3KuskWHLREIkZqoBUEGDkBQ8GmJ6DJ8l3ErS7
bGM0sMTKOjZyVW6hPOk7bOjSipcFKakPmFZjXa/shQb3dliYsgHUa6MDfbxrEnoGBTAAtBO0jZPC
/v1/uJ9V03n4JjH3/gy/s+/gRLRmtQuxlns3H4mQiUSlVnwwVYCExjxTrD8hR2/heYR5ePig6Cne
d8Sj8gZUIfxSZ1Cjzq3i3XDoYfym+pbwgcGaM3nSPiCZ8yUcaeovurtNWCCIB4++x8CojwhmQfv+
jZspGdrd7ziAFzkLFtFPYA6j0VtLjNLyLnPnMH8JZwcOw0qyDUfJRGS4/Aa2FfRKgPXJvH3LyJy4
rfBiKqbEHHv+G0eCWbt+lFj6GcdZKpe4v5mdvh//XjHMR+0cKAW0zoIo3GKGMJBx2xaPh0TkF1Cp
H3MOb/SF9XsTpZ5ljGzhA3PWo00HqY7Q/TST2FnITZDbhaIWCHR3UEj6/jg3bMzn30TkSlF8SWcI
x6Kx89lZTCVAuE/+35r7/dq0hCT6fi4QTM/3hXs7cn6dUI85DJb9gvRV/MSLJnOOtGDKWZLq6Oa8
X8zNDATOEJxDu4BFIc78BC0+e81kZOmDPLSytjm1OusoO3Ub39to1JG0bubKUnPxfumzwEnu01n4
hNZTq4t23O7plKqeTcMGNezDdiTqaY6zmRwujtCwJBi4Q9J/kZH+3FSxpwqsJqpFf2RQBWTm0LQO
ToCTI3e3H+YZCnPna6ORotX8OKI3hFHUM/LO6e/mwlXoSCvQ05ACurGX3yYO9AYmPGpOaQAsiN68
UI7aTsrONxRC8TvBCV7POaz4sVg+zN9Nso0oMY34dY2SUIC0zNq6Rd0wL8MQ7JoKMeJa9190yznV
U4e049Vwp6izvS1Fyb2yejDW9FNg9rfJswRMA9/OeAw1KD2kdjDzjG8gFY5pAcDCwSSfxBg54Z+/
PK+fGPIN9Uos3UZ6//EARm//paE8XT16vzKNX+st6rV6/c16tDxkWk4J/3hU61FhpOL7PIOlAvIJ
G/IltblNp8fEAuDxuKqewtwp1jKmkn6F7w7ExvT4PVYi9x8c8McSd6jgEYx6JWIRO5cC8X4d9Bk7
90IfOJK7bXtZI9jtn2GPn1QlxfpjYNGmk/IcimuOGoKnsU9WbrTjslB69bRxufktOxBmV7O5vimM
zj3307N8LTHtylB0YleaZWNQ6U6YEwau/2drDBz5v6mehzJU6c4s7ASdPXiYofD/ZMzFmfAdxy4o
3eju1zbzhHfnzlyijxQQUprM8XB/NBx0xSXKkoN5qYRDqpaEsIf2JC60jCRumjvWA2waWSk/PKTG
6hlha1jNdV15IBrIByojMSWaxt8zo2Tj5nuKN52F5KuVOEi//7fNQUp2t4GMlBmRirnBT69pl8X2
gL9fa9CoV1cm921RwSyAbfbmTq5vuAR96/K88NA4RAbfUKwbnNQesKoO+qYpS/YHSpK5cWjwOIl7
Ban+Pe2VhkEafhYnU/6YRQUS1YzGtBdFEqPxERCmEBXA3GWj0V1xTtMgSO9G5NCBPRCGSux1L32N
CcpcmS5L9ke4+NZ0P7z0UFBFECn/ra0+JI/zrcwfd8xmGbmDVcfiR+b5/aF4n0gr0/Hfkkv1+sXo
Bs9Hmyg+WkyVQ/54SFQbZjhXE2dzDkpGB44pwoVJZDDc7naXjZQi9U9qwe3lR/CvEY1Y6GE+iX8J
syTXXSabALIqBClu5a4jrfGVesTHgdZkMYg76ulj9kACUnEm/F1aZ5ogDNpVf17CmSGxuSiCNPsO
gd07TcLBnKRQO/CCfeg+gQGnst4uvyq9GEN5vhGzWCM+/O7hPcKxJCPfQ6Ed5fV7KipM73gL2qpa
msJIFfhEBEUFdlkiVKYY+2rZUCyWznavbmrFijZE8+FJkEQghFjZvCQGVoEFSF5GUJRdnJGdC638
aKRtnaaYO80+GcTAhpJxlQfJb5CE4+ivF0s3GpH0DNRdzGlF8EgYDJtru1x2v7gT6XHka9ajzLpO
/cfMdp7lAlbbot746VkALBOnTy2oH4K4qoGtiMCHafUbnNswCGppUP70lzeqA7JaHP0ZS7nPUXSE
cuFS8CzowJ2FY7l1jt+rdqFRPQvEmKJqc40+OvBHmsQUqyTkvuNzWQ6/mJFV/i0uuodTah0t1z6G
dtofIkai5QCCttxPJQKQ1k3xi+N2gH4Ky4J2GtLEX6cleceVMMXrCJIVa8h+2jG9wxt+TGJlUUNH
8081CwM+7o110FsUtwkjhNyH+jMc3Ig9J7Uwim11dRGGXm8zlpaqR9eD0WIjVa+u2Bt0HeRBAc21
SpejQIyLF5HzWAwvP9vas4l27xruVuahw+lYi7BLtDBqrYuMxCMCHJJTWmkMOOpTHU3CEHwTbDmD
XiXKN/XwAXCT7zX5mgAOXKblVP/XijvaDvRscT/ieouG+zwODMQhUfnHWZTbbrpcrFDHfJjSaAoo
S+GxYRbJKPVv9pKMDF3p1oIeArJRZ38OLdogSJPY9nLQUNGJmVNuCEALDre1JYbVdD+cmvRVkR3e
22b2q+s4KdhcrteudvcEX9FJBMoSezGxi86TZuNA4aeJWb+8X6mr5MqqindB4Xeqb5tO8pDiCyPp
j3K1BHWPC9X8DFwqqQS31NliUUQ852foZM1H792BcYEPgZA+58tNJ1gSGaqzgadcMNVxmWBB7dpy
Ek0zn5b8EGx02VVf3G9i0O8NGnf7ixAa7nJnH2VPwoZU8JIVYzfGAqHxxxacjTzWxVle2aYGplAE
p+pVqvDcgkpj3btZkSV6QHs4/ByMmsjOd+kus1CFo1p8Bxd43ibLdodUBHnAKYNbieQfSaaxXBlu
cP5ks/ZQCmsh2CSXVIn4srQbAopRJTCISn9pPdT9BoHbWED7xNG6AD83aWUESY0rqaXJxQNKLgiU
KoICKTEKHBPmfGvhPpBeiCg4x+PzmQYpmWWweHxfo9c/8g+9qMCLlHkKhld55Ax1sP1oN8f857dS
cbKBVyFbf27L0WJsgR1zi4/EE59/EWzomQ9YBt2/bPpW2RNjylmjZilXBJtvG1xNIOa43DiCVQjT
67GBzduaJzw5v7kQuLX1kmdlRvtozEEqfVAaphEN3G2U052FoYsNLxUxcvn/3arOWDnuC07pxWsN
kC5JtsSch1PB6Y6AshhADZWBOcriwLqMpydzaN//HVkkN3QLhBQVJ+fiamH4gzwTW1uUGaScPdKY
V1QvaElTOMkqkdKl+YnvEE53SyLLH5yi23P0UiXFbtwtd7E2gfMHk0+KMX02+dFzYAVl7FBH+li7
7yu4AOgzxxLCiNq1pUqZR9GFI5bQz/BT/rhyZjlBK8sDJeVwXL8htiHPI0IdTSBWLefhfdhj+HuX
VrYnkRbhIgI6lWxOmWf/IS5N/TKWjAoF0phNdC5O/VmFP3SGw0cLvPYhCHWegoy97IrRB5fzLCEx
aHhDTS5DHLwzJo3ATagfTtNiUFZ7vnmr3KwbKFQ0c+1jEHeVJkOOwQkMvHfH1NTPjOmJYws8WKmU
PAZDbXI9lksHY68pD4LS6FdKwFkJSLN6+NMWKpcNjYlh+ZLxDERXXnRfpBycRkUPHRi8EQsKKZpV
IjkoE30meC+1g8BgZgI2qLmlgEKIbEJwux0FHddDamYGxBctEPwGKuZjPP3140Kn3iXpTYSNZKRk
l2+03YEqR56rCYeIUATxrkcKF4JIPZ2/2Gt6EMfAdSPAnyczALzRKhTBMDJEQba3W2cDqS2QeSVm
Q831qg7ANHmWEO8AdujGipJsKWm3wy9F1Dm2UUzKXOqhV0ytiRU7I31M8hgSPUASom+qIYJGMeiL
1gtuNGmlBVj4RhpwPmzVmd2Pv7zp0QcbU3PWzns8DY2CIdAU5WH1J+LcGzI/7xYQc8Cpp8bNl9pV
xSjaJhWis8+5bVbyjfdm5fAe5O/KE61gIrBJ5abda7mFYJoI3Y3puz4NtcIs0T+gaeZh3nSJf4UB
Wnhw5R6E9TRYHr49oJ7JD24DGYCrN7pcpkvhUj99R3+iJSy2pOd1zUaSHTrZkm7Y3ONWebX+N2r4
DVkooIeQhlioyz/yNpgj+C3fbT1awQfrPvWSqNqnISQeUKlSQrCHtB/aw9DMNUcgN7Yn3lUlL0gO
TISKQelL/c3moe48USNq9IsBPyXs9eV+ZyTIt4lTpQmm7gUcWGNQCu6BhnxdjWol6VSZFhzSRD0W
eooTyFxXZF85fVrMDF84yjZ+DBUWAWX1EkCEyGk/0nT6OCmYF/a23ascl20d7lLUtwFvHVrxYjuL
y1+O5MdeK6/KmEAs4lXncBHTtTchcnnLDsqVJi6foKvkkZaiiKZr9foG3oTJn0SffBfHQ9ckFRLl
t4ct6Vf7/GamCEH0JWNPZS2nG4d1dQMy015rRJ9gNDe5HQbVhhdO7IuFbyJQDDf1lZ2q8wMs/Bdy
z6K7IrZfweBQhPVL3jD58KGVt3IRZ0rQ3lx718tvXr7WcSJ8W6AHAJOuW0gF4rJa+4uZxa+y4DBO
JeHn56CM3w5nz2VKKRhA4xOlDLet1TdccVFTFsGuTLUOybGhJSBto6KvgTAW9/8niEJCMtxBZQml
ZQN/rXJpzCcw6WFfawVc5eVXXYPTGSkVpmNTbslgNMgxnmCb+qFv5n8baT7MB3M3wBB7PQ3/fIEp
OB6Laz7LgwUsDqApsbxaaXDZvxKigH7YybOynVeIR8GyhvjDeaif2pfIEvFVFT0LMqoxpEJMXwpu
7wRbwGUm4BkxEg9D967a699p3lbBXvjnvJLXL30/PjUCZ6k3ZbHUdvZo8/WT1wzzNesb0lBGVZFi
nVDbMTMbVh4z+BOzp49iHBr9i9ank87rfqgtUqx0s0YVOsGKCky8nqQCyk1SymViohVLOX6C3KH6
jAG5hwr7QBdy3c37ios8rc4apukmNiEVIHPpRj9IvqrG2AcaO6ZFdg4fsAlufuMrdjeUbY/wA1wZ
TlLBPHiOC3hNbUc4ZGr6GYo6s/Y9l6tL91Rw0xhdkv7GGorXy018OTg/bGsszHyLBZrRt8DUtbZK
ky7ZvmKRAf4Hgdf+kfgWZbFyw/edL9D0vk9dgb4B/5zNRK7wi2rxCJMSSYpVdqByH0SFB0TCuZ32
C0ojKZvrrKWkOvnnsRIiDgDUhayAUYxzXc54zKhtV+FG45X7M+2L//RhciH8DcZAxj6VkEC9JgF3
1SQaU7BqTiNsk8BTeFIU15P+QSm7wgFnySANIzvhm8+NJX668h9YXWS/FRPBc2VlyfK9qi4ZB6LA
I45tfNM+/lmZ9cN1NDV8/Q9NWu/iKPLTaJAWg8UCVR0iGiJZ5HKpwQ0BkcK8Mr35aaOgAZ9bJhtw
27UCIn74a7YXtpbOerh3/X3Sjb4bWqVYTNwpa/q2hc++ofxHiI/ZnXJVbUJPMJGU12tYDlIaA092
O+H32pnjw8Py+La3SmEPKAx9x4vyKPVK5BkezEtmK1hZ9kJMe4VGwmpW0LqYVDjt5UYGmaRxDi9R
SWxrdRH+Ne8vItNy/B44fb99U+Sh1wPKUV8RxTbTpBGW8xvBgOLOtm7Iv+/poEDXMACnPAMhscaH
io65cxRPVYKPwODW+E70K6Jkwu3Gim+tpN8I8h2wKzXB1hOheuIH+n4QBOVKP/zcAbkq/A8WcVKL
6IBDw8FJVD+0QGaRvJj+GtSCOiNzv/xuQWzwpDVkh1ZocKDql1VLRF2o3uTJj4FTNc6gLNQfJsn1
iqmp2Kg9qZKrEBXjvQ0t190mfMmMKOG2Omes0bB98fR2V7hwpwn9zL5ln7N7eYTWRR9ZHMcsxToa
Uhor+EQ4DgMmS6RCPr2fhTLrP4w7OOT/l+wLPCwtacmh++7R+UsF6tNLLY+rgt+eB+QznZKUZ/pl
EfM8W/FLpc+IkeIEqHcERCkxk0yntGWpOCFOYcs/LfB5SqlQg+aea/c3+1KX2y37gH6cTnV6trIk
64htj4mcszQMlGMCO52xbFQyTaGaW+Ggq2ajBEHxJZjLieO+3mZ4VjAH9bgPejAisjDXh74UhRlj
vIVcP4hCjPp/jEjMSysFxzUCk56QgcoPLAVAjCCGrr8nKbeQ+UtCxVxb+UTOS8ifKn6Re3p1ZnrZ
WWECtosLJOAu/4k6dgjL43D6zEh043/BO+7/Y+dGdyOdJ0riijEgYZ4BMsA3Ha29B3ArNb5IyVPy
lPAqZ4ccgaOETgCvx0sEL63g+eUB9ISTVuS4KVaV0UAOGf4vlTfr/UQyxejxPShFUPkdV4F+gCw7
YeWlJskzvoPAqITD46o1WpSWv+AEa+LmWRr7Ce5iptqwX81eXLa+ZQYIox/tkcLt2kmu/2rg/MnK
W2Hb2z7y6LgyKFckv+E/1rDlCHfxO7OF7GqXsSTU97JCL4Wo8lFBrskhn403ZPoCo3DuONV+Hr3o
KeOpeeKUC2mYq6Uo79NYfRMB9Re4jzjDVUgMrM7wa/SEC2ToAIsULAFRa9l0uON5ghDGjI/A4YmO
AzwtP2mvRDi8wiejYUvHNdi7aGrbc2+U7mLQTvRuy3GhOXo3ATEc04kDOZAzQMSRS7G8aNu3QCc5
wZZBE9W9qySNVN/t5B+xlFIS/lbf/u/by1K7PR3GbaCVtShRTlUl51SZfRuwGYMxxQyOTUY41mrI
2JDVxLYtI2u7LuvR3nH5CwyIC+wcql6bnLfa2YIwKLl+RGebQ8iCzCKcwyMsx0otGfiCRyCmI8Yx
tpxJjXz9sgq3aigVGyqSdxCRA22ytB1GeZ6moiT4ddk7Xx8TP26JLh+ANkWPq2c+JbQdPNpaVGQ2
Ec39hP4Ls+Dwt1Lqg2TYCBmq5+buvpAvHrx6H9gGyxfqPyt69cPo1CSt919KZG5SopQKVnMcxiWL
85X0P++86QRq9oh7hYNyaKRGc4Cn21iH5/B3twxAKE+sm2m/rAqqnDmGdwpaejQxfifbxYxBdNOb
RW4o0Acw3IdzgJTXKC2v3z+UVvijVxPcTIbHdnPe2sXfnVy8kN1AFw9cLUu3ai8qkxLv+gRZqdt4
KJSr0UC4Pyh5P6DNgh1+OabyC3wRCOgDXhPIyK2M6R/HESu3Lw/ay3UZBr4SZx90h9EnzsqYgXwq
5JDh/73knoaZHcqzIGVAa81TnynCqBLoFwMr9D8yWDlFVi1JgehhuzFdyK5vPj1rkGzszpWnNBhv
qJokDA8jgbZO2tlo0629dMkjL4LCEUaDsUiAQ+Gxh9qNzaFli/L3ERTKPUt/WLOrijTga+b4yHcJ
K+Y/M7Yiz+tRpB68lRnIp4TpvszcsbSvFwIZ6CKwDzR0Xt89kFfXt+wzHLzDOIAOwpB8L6RA5gFX
djUKUc9iQHxwGFeaUhBfVgOg5QIGU0LUmbZWJWkZqPCofMn4O9uejm2kL5xA1eSD+Je/I3vVwHaO
G9FG8QMwfbll2MWHy9T0xaiGpXCYRlPmNtoRQkhL+/tj5NfjwKjDnxQIeueCRL/u0aSHDk+WLuus
N4PazI571GZ7oIms24Hml177dN0Wvq7E6bG79h4Un9Zy3wGLP6jfFbmzEnPIJNwUFGzMq1iyCGrS
r/FRaWUufhWXiuTROINuAJmZev27mVYpMzNmhaNZrjFyKwSeftcgxq1RCPQ4VIJpW2GkIdfgmURZ
ewOk86h1VTaZSKtAq6Y3biAjZiwbPv6LaDnl8ayzHRiiI8aZpYz6q1s8dZ4G2m8ugOO84jQOENUa
Pfl5wkTwo+4BS56gZUCy5+kUyZu1LHrIvQPkgyFw0VJmU7JqTR16Z6NpIXME94QJxlX+VJVX4iWw
8U3FrpH0OO9q8K+OXfrHbfAhwhOkpzb3eP6IiPxMi9gTog3nMLtW3Jx34uGyfTmkhz8kroK5/lI2
Nj07eX6C2rugHKbTpJ5/RYo/0j5kN6NYa8vLeDrUgX0O0H0vI9aGffnjszOgWXWMSzaRLmdhTtQA
x3AWS+HA2Fj4jBkpJ6tlsj18ptyz79wLh6excKRppzQr4ar3V0XXaDxBGatA7HxE/s2mLferFiKp
JLfrbHdwrlxR83gKACBiKheErY6yCrNAb/YtBZG9pDxPDyFUuWryfxME/lXkpSzAUgLibh0PGTbg
XvURKX51muVBXp+7jjZGdoqD0qKIxcrDbJLTZNehB9AFQ+y79LOjyufWgTKwjPH3tLRDLDrYAist
+vapY+nR+JWOt4pUOGYKz2JXiLn6wSV/D+1I4Hgtmi51yYmU2uisQoZeY6i5rpCE/CpNl5AlHnAj
3cwZBpKsz1xB5qMqpYnV6tPNjDRVYmafYWXpgMM4wZFRZlmaWHUufe39yPoyOqog4ORYJkNpC0Ax
kNIV9S+cds2Lu0WPqnnFlWc2iiCQrBtLF8eJDTuCqbyw1F2m6fYJPmLorgFzVT95v4EHpQZghyCW
pIIqyPypdev3EQKSKi9+lNDH5CGBGaaq/mnmpXkM86mr2uvoxgMqO4hPLuMhLss1GwMbVnipuhbd
zoYKNtoovDuDjQI1m7YhY/ZdzXjbke7A3PSOH3ONIV1baGIzvFhKGQpkzCt2MkvRsjx9w7HWj/cZ
Mrb+J4InzqCdrZGjOHWZJOStQe2nfXfgyV1q1WCoS1kU+H3C9t/K1PIt0kgCQIzPEQ8JgPnpjtBs
+dMsPd9UoYTDnnVadVzBxl2rAVsSOUscZ1f7333O46OkQHbommyDaRFHysGRuiytG6C5piXrP7Qg
w2MpF4JGSb4ig/qnXRjgBVmQCEw5OgIVG+jPqtQm3JX/peqVNaLxsyvpscECEDjNI/S6V00nyrqP
9y1TYimA0aUqZotVqlCwgeXmFzMcpfNvL5MabVIzwdeuaQrix+iGPJLI/cir2Hw7atyi3rbieQ4S
f8v6mF1py/KknKHVWBOU3Rv5JZBppuANtCVXvRwbzjDgY8ljb6ERPyH8ZY8Ew9SkdDCsO8v0gD33
vM7mgXrYj11PXliV4Czp9WjfKebBJ1YedACuV/1KByBJAElR8096gkSJyRB1mBKovYO05b7joHFm
1uzx6NWpSLBaIXA06cPmbnGrIEQAd/q10lVNV79mv3l8st7LaCp2z7cFGo7gKLl4Cm28DH4SA2rI
Sc+bSkGuUIYmocjCmO8MGSjEKghN9TOeE6YbUuQAlRpRhNjd67ecR30PHUo4wZ1uFpeUdviLiwNV
q8W/5vGpZ7rk532w+ODxKvqQNXwMcR2UX97rbZ9CBqCGO3VLV92yZGdtrXRQEAu7OOhAf238+86E
5cbFfkRvQto9MaSsBxY633N/5V7gcK15ZPsiFGuIJUQSDkgCv8TYSSrof4eUxxO7wmM2xH1fYg/h
ksmf1LbjnBohP0QYGKJRbS1ladSatPP/o31/JW8tTut7FcKgTH7y3YuLuwvn85jX67zm3ipxyc4e
U8A1ec8utPUoy3PV6LecbwTH8qGmhDzBADE6tkrl9kL49EePPb+JXzAoWTm26m0TuIZfDqYsb7Rv
VoiKLFInuKPV6s1IvqWi79iyciDICLV5MoKiviERpVVO3HS3L4P3YC5uN9REIqZp7ncLfBcikONy
2cuxB2jeSpEHa5LsxN9ww48qDJXq0I8xdE9PEZPhC4Kh9EhpGAtgRto9gPHnjvIN5qaz4z6VcREp
KPAqbya2BRqSz9yszjD18A3aom176qg7dXUDZoKoUNbY3pkyNWoxjrI8jcavRGdO6KMhSPyqA0Ts
+RgjdLyoMUQ6HLyPLm8q7VeqA3cgps1z1wQlJ9CbvLfBZdIKR4jejkhZiO1PAkG9K9qU21td9K0u
dMtcWYzLV8vSFaqeR6Jq/YKx1EIxIzU1GUXurzjJoy71O3SJ70UCQoOPkWU0IVMkHrzJ3WVSXl5p
g4t5nXtbpKfK7OeTjKl/yBgU5F6K5a6S9uWquuyrHq0XxFGyQyA9xnIcAuaLGgFrh22fdhEBMvap
zCaE7ZxQnNR9TTGEeL7hMaEOVUvGv3NYB1Bl/a4Qp2/6oM95DGGQmwtVsCZRmNemNexN94VP0hvB
GPqQm+SD2fKUXv+kTFr3QHhke63Rb7KKtzcsLoFFIo3NCm5NF1DSrcbP4Dpi3TRlEgTcqWtd2jb9
7lJ0jJqZOcKEVoQGI1VbHIxrsAo6FtGaVtJ3Jun/Ucq9aCLSFC/nUl8GpkVjAgISuEY6KYuhUBc0
t+ac3NUuN2dkAx+z/P0P/D/bY3PJOygFsk2RlTMmTW3KWg6jVB04Lr7YvYlo5zaGjdFjGWxefazZ
Vb8hjs31lu913NmJXoh848ZimU0ybAdWgdineiUqs8sdWwo8feyN2ZBdZczakGDYqdhhnigwFRiu
fHcoGDsBCZnqpfWojJMZWPVTbUUXbvehcuQfWjGX7DTcgtYraFSa9NFxgLQkfGAV+XYnw+Oezp7R
id+yduby5gKw8EzC30+OOz96Gap95faguMeciIAifvnjnMTjmjY6kjJ+XMFcs8IByE1TewHan2Zi
ViN2IEk6RRLhn1DwkkHsTak/Y1tp1Im8ewKdvXQVG4HD+aCM9hV8k388hzZtWp+lFyJPEv4PPhsU
vRVGCMkkg1SgANt468aqtOd5UyUCGiaNb6JH/ie3uLvRb2a7Mv8oAZhK52ud4+R8CO8I0FMPhwPB
7D5D3gcrllfxJ1GCJ/qGeJc8cfndgqzNhh+abyuLvyeUstSxDpsT90hWSucgIS0/6HQi9/ZqsUi0
wo5xUrnWNxQmgoH71RRz3uS1MjZlBQFFvXwUzRMDaVpSfF5jPMiwp0Q7JY0INrBRSai349hiGXAs
cIn/5Xkz0TI2qKI4nvAsH7pGetdXkmhBzWPV0QlRZvrcFmeQqVFn/S043IiY9fTdPaDBqXFmHyY9
d7a4Ypt4z1Liv3pG8hpubRXe1zSw27MrD+MC4bUxcb7ogYen84KPOXA6788qeW9+28kYHV26qxrQ
/K7+qZlN/Vi69sLTaIfQjw6SWg188cPyfQdA2GbbdN9p4Vden+NoyaSXU8JiZdINqLeTQSaDfg5D
VN5aYoCELxjKTkb+Hfj/pFXLSvo3pEmLNYVrm4Jsb6i2OJARuydjh+jUFV6Y4QtuCVAgYhOuIGbD
or0F+P7Q4APLIKDPGkPCweiYW71LvRnAVV+X1UXRqimm+pi1/Vbg3ROOaPQHKkhkhk+Lh0LjrD9x
9C/mMCsl5YLaxR87OeYlSR6Coed5J/q1gb506Gz40NCXN7nlUHlgpBu3G4hGSvuFYapqUxrCoH5f
fcsE1CqiabzdVw4e+2J9Csy+8crCdr9vnShB/M1mp2ZovyS0H7Ka1DFAqZ9e0Jf2+F2NsHJ0CSVO
H4M48PN34rYnU5OO61b1dRHY+hOU6QrzHTcajmm3Exkvf8RmknxM8zQO6I/XdUnrpWvZc9AJnYG2
TrfSWyyvIxLhbaa3b3Wb/wTushlq9RD/yAv9P8Y6t9nlQzzJaY1i+S1z4kMlDRHY2QdV+u1/zA6Z
R/6o8T9IiyhaUXUoIfRy5OcXYrhy9pffWRl4HNQYEdagvThO1O9wiF0zEd7eECZdXPMPuaFqSjXK
WjPy6VzspVb4/V/U7P5bsfL3W9rRlbFX6iDlLOka5gH8iTmI7WtL46xPA/D6udlZWiPDnPWuTk80
o/3p3BWiAN+l8Tj2gPyaZ3Ifm1yCSzFWzRcCbTzH2+FbfqQoGdTArbHnDE1XNV/DN9Dww0UVDxDX
mmHHpNvkxmNdMU1gfVKSF63VMVAECTI81hwFC0Qe2TD7KuKiJoZb5NbDsngFJwN3AXo1VV1kxXyG
3nE/PnOjSDrwQ4bWJ+8jK2P31WzQZMfdxsALqQQhIJ/XjoSFJ1CYJ4Yne0c4Lsej/qUhGH+rlbzA
gGkfx2c/89lWTBbr95mpxcmFxEfqZ1yKz+Xc9PWgcziLDqNx8ep0T9JynU8mScZWyRE2YeHkorQk
k4uC3uIoIDGAr1CiSsuBYq1D1bRBYo7bqbyLD3bH80LdcmlEekvqejEPoMQKKoRFJU5yNxmGbLUY
IyMRtE4R6gYYRRVixG0Dz1SIwJ7BXKqOegSMeD4XNqj/pyhL8QnlQ/JAP1dJKCozVOGJUXxuR+E8
Xx/EFlDMY/o2+V+UelpwcSH7Wkvaa7wWnog7Bt8H/s2dbd3vKiXJ/hVGnuoziesFIlnsTZmfLdzu
mlQoI4Su7yuP2wKo5bgg4BPMy8XBa+ArqA9JaD10YHPO2iPYwxBbhr+3iXxg3nzvUWJBdpI0ZWMN
SndajT5t2geNskFPOPJgCmSn1YSdSx/ccy2jP2tL1Q1s34pYiONEQ2GBCYlfVwen5nLvokAAqvp0
BGDI0KpRD7jDBpFGsnSfShzd3hht0n9D0RJrAZ+H/TPxMz/liORnVVhHSF3RnfrD5frj96ZnaOtE
VdBonjnx7Fju4IVTAHftcKN+mBeVpeF/l3/Gwf4+ILum6wzxi6PRh5QiYyajhaF68KY9bUr6xgMc
tk4whO1+c+xRLSJtiihFhss/CEkSZpIIi6/K8e/vQ0ly7FT6gU/njTRQOxfEu+c/iW0n9HoLVgos
yusH+4P0c+4zLL7XeST+RctO6VyH9O/S05d6XY/sqsjGKyOqXOoBpMVrhpQGJPRuoyYRvjAubYVS
6yt97KrjNnI1TrJ/pCmQQrv/KOyvADvTrA8dFJ9tLeblzo0ikijFZJzzNyxHVpTBzZ66td96k/TP
hdJxGEbx9UXaULDV3JJCqwdfvGSEXIjWwdWOBy3MhwFtQQBt7QxfuQXMTNFpiqWoXcX7tHBqCKol
HL6h0lwztS3ZDLoeHHXIwxFQiZRioQVpmaT3cjD5kSLF7ju7GrjRlhtYDH5hoDj3Z4bPcXiD+b5V
wxrevgiCfeV4N35bfG6FPinDZkTAOtOTG0jIDuCpl/M4jcIsPDiVKSmBt8FQLcgbRKFbXsSV60C2
ABEk77Oy4lbz9WqVRCaF2C8ahZVvrpxSVCzT4IHMjhomLJK/Q8LZu8MJEXmjM1O7F3ZSpGs+iykg
6URFFtVDGM1/oJp5mCIn7jWya5SklES0IBdOsOakZmyvbY+4WegBt/86IcqNsI9mu2LQ4tANPUSc
mEOLYRDJEFM4KwQEXiCF0qa5GT7tUETWCDUHMH9ECmXd6TbDjvOH0JT73mSkVWNWNa9BNIZa7m9i
uvfU+ffiqa6q/USuVeTIGWAxBVE2t+LcPCH+Z9PuSITAIPU8V3EFIGWcoZ3z72oYKKIM2k4LOHUU
QypKoqSvfsfW6AbbNd5srZmAN4zjz9I4gqLnLBxlDf++uhggkqYqH7j+3O1PpKx4DXoU5mQwPWI0
e44Jn95a/DjgMKgc1+DlMU/YKLnQA4ZVYlrbnUhLmm+X2IctyGr86OucQYQa8JRpS3iNl130zhjs
7UEevUAhQIv/llp+w0B96y2zMXaTU0/r/QwS3ui5jxdFvv8uE/7Jh0CBYmemwMk0bnwTKAmktiO9
lgxby4HLC4CKkSauPztU53CcKi8hWNFihrV6fRO2aVoj9vRMtSaN+I8V6C+rNBuJqOL4Lz4ScJyf
3eR2R589mM4vEC++/9CEU3rBNvsYFelLBJKme8O3d/e/T7H7DSwzVzL/MnNHNF1XFtSJAPLyCOsb
5uuZ1e9lnnM4sbOUrq9oFA0oJz58zEKydxS9Wbf8W/qv1wvDQ32AHBnVAG9p03kWXmtDeLalGk47
qmmoo3Tcscnsi6IFXD/ui/lNQA/q6VmbrFWGMthL6poxHqjufNGCFhLcP1NqiZ7+/3UfvX2aWMxv
GpUPefmgR21BLou6U1t1oZ9Eq3kFSA1Hk9BLdKERnKpqAWZijLyCAMx0yd5NbzCSUnyZIiYp3cBA
QsexYyz5lVi3uFGObPgjj/O1LHo1gInRBpznFES230qMsU3C+rPJhyNWX8zKUfXMkfdqQ6M11M16
SrBaINhHz9RdKoa33KGmaMMS0tOx6qm0WGm6yQVFJFSyI+6826mbvg3U/GmRqUdGmiVHzBWJV0Oq
VZsLELONCmtTdO19z/tb9W87oNsH19092LuO1HAYzJrKkWETxBeWEaVADrS7eFYDX0up5SsXTtoV
Xuljl1C54D0XPVoY4MO/yZtN69TqUNxKDYcc3OJKogx6w/RkzyaEDY1Hq6PD67DpwbMzz9UHkv/O
CNH7YD+2l4sFOMqKNb2U1l+3KHUrHr5qhfQgFX2ErZzJolFuJEUnghh7CpjkhSghgIKh5yOJcSgw
/WZAn3R7AD+WMEm49B5REvbh3tdgXOysWa6FEoCBTC3vYRs1TCvkGKLBkHHCBrijheEvlrjuiWg0
ozTZNa/QrBfqhREYo0yQCIo4bCYCc9aEpUcnBwkd1IJwqrrk9i+z7uDLWE+fa0pxTtytIxga1D2g
CwqiIspFwBgCcPYJ8F7YhNOjYeeSkqZoKCXnyn2pWaCDLo1/zE4JiQO863ZxhTvY+S/dSCzZD6hH
io+5oj1Gjomv6Rr9iexwu4Pd165V00KzCDA0HPwuYgt2lQBR0NLb+NIF5PusVr35HjKyDlDCH6bT
v8DNxxJ82ZZoXHnaBImbZUFiCrFew5SUpqcqnF6ZxsInlGdHdM9je4CYDVxceZ7oegIdR9k8wZdU
IVZxnw55Wlfc4e7We9r40mYp7l/uNmh/l405kfU+yXSNzU9BDOWnD0MKTCY1OzsafeuJXz6bOlWt
oO2QtV0EIT41jngQpMwM9l1LuFU8tL0JaaLGbhGkrI2LlE+iQUJyf2GpHbLD15rGve8blQY5SGQy
DUZyF5TigPwCRlEH4V9jJIl4UAUvzVa1+2oArfnSes9RITeeqdvZjkEuI+poDr/ah3YjonSOjh2H
QgN/NQdtceYLrNTRp+zuJhfI+h8I5RHroVGBh+T3ZIysdtdhlCsN1tpV4BBiEiviVbA7bbHtliDR
wmsttf3sAKIzkSgAruZKLhkSbxgGgjQmNinAWyRFbRKL1n6cYFho9Bei6szEvN4YnA5Cb7WED4oI
OJc2PU+VLzIzzDkmg39JHgvTN7pssCsZSc/kg1elPNBZ9txbgR4w2M71MRGTFTPG0pJ+gtP/94Hd
wKAakAK8sqP22/T5L+yAMrInLzAIguJjYfVpebt3Mrwkmy4a7aTB/3Bc9ZeMzTwxQexi9U6tT/eR
PHamKyJmq/AyfZ2uUSqKuvqIN9POPEq9BF9TDL8VLaoF0T6J/EmKZHO3eDw7uNJG+WyseqVchdtJ
o1PfPlsJu84Rqd0aWuXrg76Z11/U6+bIJ+E7pR9XV+6cEDIxVNajHw6kTw146E/KPhw5gIEMrQXb
yty3TZAA7lERoePJuov3LfxNsub4BkFrElAKL4NTc9O0n1I++UvUG71n2WjbzC7US4LRL29thq4v
ApM3qxtTc1cneBaXLSYrCU1RbkhfVrmLd5wnyVg6iNg6OgfuvnBylfR7WvNyLbscb2HIqGDkUzDb
Zmxqx9Hjl0nDxvp0c0IwtxDuuhLQKhUY8MbbjxIYlZBoZY73urrMvOY7mvykbZCH02hXO6EjBTw4
T+7vZdGxjbkH16eM7gaBtL6olJ6E7+BnXvc82sWDnBFghYVWEZHV0XO4v5n9OX9i5ozPmeX9w3Hb
PjsuTQVXcUgOpP8w92HkCAQopMY+zORkaccWbyyLl+n8uQAsdx0FnO/9q6u0VfX9pqz89KuP5/mC
MLjRC4FrhG6W4yN++H8N2Nb/anIXxtOzSNqvV3LltLXsDm3YELaUIGpzH5Q9XW6h2c8f1Fr+fbvA
u4n9Gm7xu4xRSAdb4JxNi9qRzgDr9Nj4Xe5OaqCIC9axDyJQvG3T2pDfjj38+G2WsjgbeNpXzI1R
/2HggeoxXuECw1iZSnNvrjPB8Eg0nIgrAUwmoFf0JHq1OXagaOeSwtUbNxB9my75BuQgXHjvUPVO
tQ1vfzlHZRFayTclDI5o/njx15RIE2cXQa/QqN8a90+ttuZnjY1fmPCilIh3b4RA4/CgaDy34lwy
iG+MNhraAodmjZ80SMHRbh9ZKacauoE/1tYE5DkOBA6yzd8Rcc55Ce/ahdc3IGnNTxMukuy5DRb4
0jbUDXkYnGpHNYhW390UvWifONf8V8EM1nEzJj9Wzbs3zP1UlLFhvLERCY0DN6DkyjQlGls5m6jF
9Gp/Ra8fD3Yj9fQMa4gokoDNE6PoffGeWS+9BMRnx27pzD+vHO97NMLGdxQBNKtFRAulZmYQVaC5
/MtDynK0wXpX9+g8Wh6sDTIsCL3hsVR/o216KEmdEmzjcaVQfTJqubdXOlJi5k6LKUP6dqHv5A8k
FC88ONXNC+oodffTUcLWHGv9gJwwRoFuk5MHYjfMAIoG7afOP3JBtpceul8+rIIwoWHOLfeVJh+V
f10+eQGihOhM3sfifBhBbPOv12TAN/ZcVyfjaK5PSAimg173Q+roLOjSVn1cvFttLamakfo1fslg
6BWrsM+zIhPzsUlMDGomsRfQ9iEkvcakeSSXWJCpQehhkGC15pYdrquDuIA7ShzQCVgmulGvGqam
IEpNH41zwjMAZMmrjPHQWkdcIj3HzRhDF4rnsF9BPbFw4MqmEwmuOMwr/s8sbnxNFTevZEFuutMx
d7oeupabIqBH0lDKbWTimDs680lnD2uLGpzZbPDy1i2nSPL0kMDlly/MMulKSKsYu6rumuH82MJd
uwH9dd3vIdK7hUfvPu4LYNZC7gP75pZivj5eh7tvtMxdBbkn3N6D+CICf/9QFGVGngymk+hedzJ7
Bhs0VzeB+AmgY/gdmBeyGAmGrBYGnZXnxWk+06e3d6vPH2vxPgR1Jm67VCWGziUX/9oDiRy6XNl7
P7U3bEioyl3HRAg66+OD73HeC2yBYFx1G3YbR+bolkyWRpf/TBxYnZAz2AUqI5UD6PkrzwEyBu30
pzRYwiUmGGj2OW7XzzFPkPkaD2aEbP6kAxopfGCGVgotgZaCLryj/s8m9hCrLIN/ODWWTOt6qEN5
WB+7F0361pm5Z9aCjDmGLhUsq7YTAAlTrzkBd7b6duhiuaEKZQQQYdP71AJVzO8IPYgnGcDhnF8F
BIT2GFjBXIjZGcxS2DEYf45t3WBphP+URZHuum4gb6Sb5dHQAtUGIZtNdVSfXloYxsLmM50Uf1EL
DDtmJK5ix6S5dQCE03fCQHPju+OsyrJvghqTw/F0a78QQz3gWbgqh1qf28N+tb/Yxlwr0Y6nZLl0
cGRsRgAnfglYXckqB9xZ3+Rdt/Cr1h55r303qX5YUCXc6hMGJ/jH5XxVu9twv2+laQcGUELPU7eg
YdUIPrZA8pKGpnXOaqrGWjRZrP4kNR/iNqrr4itRxwORzjCtdgNI7FiIr8lX52l9g17LQ+uzSuqy
gL7TL3uoboS+A1Xhyn3Cuyxj9P5Xp9o+Me4P8WlP8XCwgV80OFoxV7aImaWq0wDzbDh84ecq2A7c
uctcE5qQ/tcsA2XRJ4xD1gtq4bjKcfO067GFriLTAw7Q34pV3SNQJf60XglqvP8kMqOdCeQCPz7F
wBgooR19OogSP97J84rQFgxzjeq3C8+uBzPyWAFwtxu5nIlkXIN7X5Pr7jTo4x6h8WfBTQvc77Ui
BwoMQIELXWRyp8NGz4JjvY9k9HmfyU/RahWJtvt4NAJda6xCjIEsmeuZkagpLbMru8DlZlmDrXoo
dyjWzVhmCnvFGSPQyLClg2bIm9YpS4Fm6M6t2Zpb/ROhxvCRfMvNLcZI7DLtGwnLgACL0Sp4jhro
fN6eJpXfPfnzzWxoLL3+HjMxIwfr1n9mmIdo9tIH2Vn1G7JIZS4jgCDt+LHMHcIwKDK+wSWU+5IN
3J9L/JmFhZsq7OuaQXucP7W1YqmAKAG2b9gslroAoVY1jJDgcMmkhTvTwkWlH9oppqkHYmAgOpid
ML+wSIOiQUu5Et9wPuAD0M5mhFWbOE7tW30DQwV6Gd4SHqLuA7dO8kEgYQuSI00837Z3V4h/KmAs
P2r116AC3Pxe4vRbR5anb2PCc+2g4jkoFcKla6RYXWsph1Nxl1aXIXp2QMEF+WgwH9v24lgme0/O
Cm/44Re6F8NI2yiEJyKN/cfjve1v2dZJaRBZlj6b8jW97BHYByHpTN0rzZARSp/NReG0du1Lwwbj
AGS4aRG2UQM4yzVilE9MAdF2KTHhR15MCyDwFCoyynP576TrcJuptUOc3zqs8Us9UM+0WHJp7bb0
JS6rN/JlWaHf5+AWuzj6vnVY+g6vyDYFooCZmVn7GXhmet3cUm9S1FIETBpMo48Dk5r9AVTUar9K
y7YDuEueP/Oli8myCdaRR4mo0oCMeCnmv2EmkMvPOcK6SEqZ9z8hP1yBdJd9IVkl9ie1gYUPbftt
J+huHbKxqL/uVmu693uEzXPKyH35LFANpvIptHfgguMc1unlitf/3Uje6zawSr0JfJnRd9HzbEGy
rhs19SmNvbfB0+1ahrFI52aZdxZ64AgbgitZwC1Zohm7pwXApXOLR83+k5L6GL7fFrHlEa6e4OTi
pjoI0BEDnVn1HSJTiieZZlYWpqlOVUDwRrJ7uCczIfeLaoUeTAO97ECrqX1UJjzk3hHOluQi0Ogm
Ofn4kyGZLfFxztOk80j9V3q2VYHSRAgZCfhUapTj/cJx1Ibyj928+qLXjjq5qQ4Nu1wqnmTjXmoA
iB3bFuDH8CZ6VZ1inT0KCMpEl9V7RJtCDMCqvUm8vcblF9Mdf2g+tft81wu1ffg3H9iLuaawRXLu
81rDZdLEtJxcJINZ5m3n6WbCd0gXgbRUBag0JQ2VTCu6520X1lNeIoTcUZaQyctOnYk+E/oy+OQI
T0GfS62Q2BffMJn/weKODnby17I8cgmMxPQRWoh8fwmLuMCdsKwa1qhVx02F22rx8Po+l6HvWF05
MiXoBsyk5UMFWfS6Ei5BBMn1q0PQ4qNEXhNLEZD1g/vcYGyRwJOnVbTpxr5MLyelmZkwksnYYJWZ
86HvUXMNf2pm7v1sg3KNG0SDEwhAOVULAhVzQutrh/wxprVoeARzR8dQnhsmEmQcCl9zpvgFVtgO
z51/AkK15nlC+EfWW4llNRRFXM3XXR7xWQEclS+DpyudpTfi8Dw2AVTwl9H6VDc5omtlsPqZJXaU
jUDIlc4coym3k4I0MrB1urYNODU3NrD6pfQ30PSMdJlttLiH0/HbQMNE/+wBAkOk9xQnJm3EBJH+
yODfPUWnuuSF96bVL4terFy5W1f4LqfvgJFOk1Uw/bLdwFf1RBkycKkkOmul1HT/slp2Cf34KJL8
h/+F9m+MFWLvEGEkmNHKP4jNOKUzdG/bqs+riXcjU89AJ/k5ZZjeO3FT4g9W+fHGU9j9LGZ2sDs7
GnatHmSxKREvNG1XCRGuNZOgXPrKZYJk1bTOT+t0sI8wHdRc81i6RWKnpV2Ejh7QUiYWHIJLKsDO
BJpBdplBpaA0wO7qx6lzbChHPMDgsKNWurJ17ZD4MmFJiUuqp0l6yH3uynyWvG0tSXSoS7LedIGw
YdbYIHKYUjjWLM6m7QP2isZLTLOlYG+1C0lCndX0qwXpWpkV8l2+1brbfcFyWnoIn+JXbq5gLA+f
XRVySTPDnAIF5G/BCfzmjKq/nw+zDgzDCxRDtxcL9APKfj5FFjZKCS9fdwIgLRWNfUTO2S9oYoZN
+D6WHp3T00wuTlFfP360KClCthGEfz0iqyPj3KUALSzpdrOpc4w4s2+9ABAufUSN9FNIbUIgz7Gk
QuRd7lVK5Gd1l1rK8uDkYjouuhkfZQ5lElMCW2Qx/L4HmddzSjXKl7wIS3l63dbQSwmD+UgCwPPo
OziK3MvA9id0+0bZ9K60H2PBDkjnGtsvSMCSyPfudo/EjIQVq41TER3zPpCNU/9xF5AlTHYbtj3i
tnmWZhSf7bDLiP0wqtNzNusiwsTbTfJAolTZH9bIvMWPGhq1+43vbXArVl/oHQED/58NLDd/TSZA
GuWIG5WAgsyo4OFoznaFTrF2RPzDncqwnNzukF1AXKRfMV5NCWp64xWCc+sjDXy3oECYJmVm84t/
QF47/p8ttwnOY4yJ7H97XTQ3+vFxjQldYCUNnp3WW2v4oO1zwxIW0hTB76Ap2gCtNtsWsh6T6PGj
wsddHemlv+Kxp4HAeC4G3SXaAH6t9g7jFjoyebjEeNye8V5JoszC1Lc7QeRe86o9CcT0IYw/q60F
gl/Rq5HzEW+D1q/jFW7DJFe14A0EDdMmgfz/5jiWhJ3ZUxIRnqogX7zgML8mXdxEHbNzvdek3c7n
Kr81IrLuwtY8DSkp6M8PShChBaGZWnKKR/cxHS8kbded6SYt3hgZuyjmMhPs81yaDT2MztBCHwHI
mh5dxXEmG3719raYeFkNVaCr6FbRjofmN4h7wbHkZHYZY+MsCVWhMkP947ArAl1Pp2EtOJ82BshW
S5H6not/sryk860SSYsAHWbDK5cZ40UVucK+GrcuKG7i8sOmqPids1HQx8T/5yfahg+WS9WdLVDN
1wjaA1YNsh0EPT4UYvxKgXJmEyMwN9lF+CVizzH+1n7fQOiFDasjg7nyqmzeya1VoY3YIhiiGDEg
kyi5doHcniYb5hu5NkWvtquaXJYcHAGy7dP9MlRjk2+nJPpeP1oPldGBsefsCaIv0RkmoxHygX7q
8uNr/GHICdg8iaEVD6j5SDGd9rSuc1hnlyxA0Q3t9bfhb9S+FFhf6Cnw0/MxIdpAo6EKs6p6PtAN
HchxLX8ApZ+XYY4pQJ9HlorDeX/RZ+yX3vLApJa+MQwxjBjK5luv+JEQ6B0mbmdk4+KiAv7F/JoS
e1e+WHuN/LQ+FG3vW4SGiPSkH+OOGHRdrSUdE0OhOd9SVy2pYP67u3YOxJOQEXy2Q8SwSvlm725r
PkOr1M3kmWWcinmSlnCmcCwiICtmEVYO0p7iwmKSPQuQK0W3xen2Zm87Io+jHgefsdXLRbUz5V1W
9ESyQT0avmOUJz8QvG3CW4BQHVCA0np8qZHE/GUKludZJAPNDTzbl48zFzQL5A7NV41lFrVD4YHq
WWT0D6qK38JViM5QTlM6/2IrQYw5uINU8wr17yaamFtReJsBsADEJq2h2NryVJdHLhLwkKiDXRFu
5bWdeI27ZKs52BAIyWKkWT+Go6nY04T2wkskGxDE8G4ViEBqWNXYXIynAI1pw+Qi90+VH01XLn52
UywLuyJbn4i2hc72M7epxFCWsY9hezsk0HYMBBJsYWgGVhP5PHqt1LT+e66xNq5CraL7kj0vke21
LEGDuMqxY6dwDpvFBORxD9xePbI36bdKhOX7Trtx8e/slKEPqjIqhKaV2O9nXgRZTPwUSbqwEcW8
6KKzzx+MOxlBgzt4uu2OGvTvYU+RKvOiDWxaF/k4SkMnr+y8rgttkuGpV+6bXJQ741wKTNbVWnCQ
cQs+EfY3GpIjk1QalwVRThEIiS6OywQ8JI73vzjDceZQolxjkv1jOVUiUcMS+xU+6pvCY0lmc8XG
/y4O08lEW/07vuXTA1BYPqPHSvy3i4dPbREr3K4sCTKk5UV1fuQI+weOmA39dho+rfVz8GGfD0ar
3harP3+MCPBBte7xdRUimrztucHtPxuUazywvrGcVBEOyDkX9EuDUQR13rsJxP8ZPWA0+cNkeXTz
C6gnOrtPzCxYKPzLyfQcdNbqY2ztPHVtk/61kzgZVqf0acr8eGtzStT5I68jmghesikMTEOafnCr
zlMd6skS0J5MIi8QZxafmM/hwissB5ZtOyTQlSsfaeZbtfyqNkLo2VvL3O9EfjPD9IPlg33eIR4p
QkY91lhHZtXCJgw9FCnseMuXCsXUmBT1+VegctK6EJ2tNXwRfvBfHykVNzhFhH78FIkuBDyB8RM9
GGQqU+HbJ05wS/S4YmVNIRXeDwgy6lAuYZLE8CXE6se5rFecaFOorAE2pmsTVK1Gm2aVm4LM6DRA
nOg9Xu6qgsMnA+MSvUdRJRvRZcAE4vDLrYR7ipq+dcyZlYarn4FmPzu/1HijjWerboV3cGl5j8du
UeypI8X/A9D6I9v+GGqTC+VHiU6UU7Vtpc2MrzcIsNcRrPdHkWMD8ZGarefD9B6AGvdOvoYWSnCU
zSQGGZrexvuCihSvVHItfKbkZwEb7bPh8QD42tgRTtAWl5N/fsoA0xi0mrkLllZTsroGz0LNuGVN
DygdJ/QUrJAkAMxGZmdboMi3KnTvGmY/3NnNa1D14qA3jQ6T6xXA5JAKjF6McQbgKx/js9QK0cAo
hvngvq+tszkMbdx/a6iI7N2e3it5oYVuz1IEImoSqb/s0ejGNf3COpFzeEevoqwjRBJGd5/W6z9P
qgnogJL28PdgxJo64DftwxxYP31zNoUdsyD1ZycLlQLe7SORWD9/y52Vb1VwFxYJexxfRZgocviO
oSmeXjFusMOUTInxShKhUedy5KUK4Sa2C2SB2rIler+bMZTem1a7yCUndXKhvhxGahyL1LlgNGvS
DSf6TbqTY1SYpDdcxEyAnr5FJYw0PVrKaErTBgdS6oBktv669od+O87A/lWOuuIcunSH393HOwPI
9JXKCNaHFykGDc1dNbFGRyLBvKtAxwK8wmlhdyltGse8AXihNnG4e6pYkLeyvpeJWaHVjTu/wqk+
n9g5AUVFmHPfMyxBk7NCKmHLvbYiDf4N3H/Zq/etRVFVtWWXzHu7KpMt2+PMnL22ChH6BySyxUNX
pLvwFD3Tt+oIg6YAeEblP7dEue7+GHrVoSg3CBooYZFKdUFhCUZwUsQddZi/WpNaYZoErDNmfSrt
0KCSTvKAHe/Z+jJp/K55UxwzLbM9TLkI4QrO0WgB7XLRUIaKHrf3I9LCJcICzTaMQpx7YJ5iQiN3
T8x7zepfMjgrIb3+slEJzY1oi7WISaR6t5wulsZv9JGDRrheDDuItcEvgdCCly13BPtVNH3YMPQx
oJbEVFrijSJzG2bAe/CanglWWzYc/1MmjVq1n6L4UC8ntfJsWG6kSDjSw491dY8h4cS5a3mOBmei
dXeHpv/kfhmwu7r1RuG+vBMVqZ7AiIhnhZ3sxPHJs5SZpykO5vae0nlaapd10bvluQYSUOBOka81
p0R0lN7egI9nVt1DWSLbhb//FQDXr+JMD4KEE3TE+68Ee6Dcq5887i+1WlWDAWCCeVN8aYM0VnN5
PBjKS/PnNi2hNFd0i9HeN+z4g4Rb21wbNZ/PrQVCwGFiWD2PNqG8hQoKIE3poCADvDa4pve87yLX
jcxmmgWb1lBdQsPlOVNroWGc0XCFVSDbHRU++k6dNSqsEFy94r2e97IgA8nrYt6fLalCFRxCMQyX
tIwGcV/93dOpyljNKGC5CZNlll6TSLOaapUx1N79fUVOfX4nZe62kd7E67fvIIswQqIafEM6VObk
rpd7qLzb7xpU3emVsGmmtZHMyurSRfRYtndyiDeQ8fQv8v2MEnUqDvY/VQ088p1GNHdZD+MR1Uge
WnKtla70DgUXUlMxT/HexxEY09RXQHCMjUXha7Fg7iJh8xNMop9kvQexIZnPKfLKCKSzKH8PHPIH
OIVOqWM329AOYW+tZDlf2jJ33vFnoU1t8K15RyQ3NyQbe6e+VFBJu0LpGeSPoqWZfUZ45vSlpd5X
HNePgySWKhUfTPewSyQ9o0xhbDMj0Z+DbXnvOgszfFPHuwNuDUSuvA/lf7GkYrqEw0zWsvMbHBAJ
mgyVOYp7kX5VbaWcpVMGyWZh89t19HibXbrNOhq61X+1aHhGuNLlUD2UQbLGIXZRIzXCbiVMkszQ
3sBI5urC7Fm+ps+ipB5RYCQZKphOrabsIe1OIwZg5YlnMPNRSVRwErtaxJAt+5zSlO4/P7hKndwH
SOkBgdVyivBPHkpk2/VCXkFxDVf1hhB6TaS52cgNbgOtAqUuhE6whF0/MXbDyn/wNr4MuuI/AhUj
x46q6LqNT0DFtUPLbtNed6aIUkUFg3sRZFC8isyJq7d+b9jc/iVRai1slsWRNygUyczrzJahG1mM
QzvDkqE7R2G9kjFN/70ExGdcE6XG4gJjdoKpuy7Om3KP+1A2XAuHC1MBWXOlH9mfwj2Eoo+lD6BM
FmRt2UimjBXFqR+80MKp8xN2DgPWUJopkUBWKnaryyXt15BaiM1UsonCDdiZcCGMi7Kse1TeqEAq
A18OnK76uai6F9UEO8f45+HSbJf49zH9V6eMP4MbzccR82JwIWF1Ra5gU3ohagqgT1jMpUZKbt5j
sNgXFYpj7ena+iMrOarxU00pE1eWe/8MFQMPqzlyZ65sK44MgFdW+pL/x7l/tYpP4ouV1IoJ6mcA
mlO52j50u7+MIGEvFihVsyvd1fgSETl/aURj6NUFJSrj3IO5HyPh8aE7bBgswRguk1l9RDbgOEmT
ZH2pSj0vtL9fxuY6P0for2Eiftg6qAEAYfQRfy8BNgX44f7/payyr3e14ZrvurupteuasWxnkLQP
x6XVMmDlBe924AF3srn6qqPlDYJ2gY7hNBhId8MwGIUY3f9T8FRXOXxCOaVcjweZZb/6bLQTA4T9
b9c/r1VDYmrSFh7lKrPeHR78oTE7wDmfxgZKrtFHskF9BwIhrO6xILdkEQi5vSFpfUo0TEjWOBdN
+FMZ//whltw9cgpXl5pESvyJM/OSKE+GiJGcE68MV11Jj8QfPb+mE094ljx/u/zLf1Bnr91WOtQK
o82JT4oxII/BtTR07kwC/3Okvh5RtCak1nuQxcqIiif1N3FaTMhKVY4r4RQg1wSF4sJ8HPIDTKs5
m2gzpN5E6hZvvA8gl5Or+dBiHF23FhVpGdTlzMb09M+HScxwd7VT6fs8ciDiblS2YpJ5FuiAJ0fY
KXZf5kfPzkS6+THY74DBwUpq20EdqKuZI/NQD7woaepaiNYtZ+iIXXGzIfjyQQGyjhlMHKaQ75iy
zXQF3wtiD0FustJZqWRDjYSKXsDZZuQYlzPktyn9+PGSzHcfaEREySiHUXKp/1ADXbANP/4o052r
eI3OaVb131s1Gbdw67NIPm/Dnq1HKTO5ngi40vtUBzUBxUvwtctqVeyrtjEZ6DWpQGL+HZVGK6FO
YMWeUHNLupiK/ewnpw+mJxp9T7NAX5VpbxNE2ziiiOrhpBW4Out6LCWSY5S+NignVwOTbvJviOfO
aYNA0DYg3R3pXQ0m3j0vUwHRwaysMLHmSa8nlzf3RmY+id4SD1FKrhUDWprgTP+txSunmIBK7Mx+
o5nZvIVQHJXxejkW37vdPYVCLc3/qh6/cKDttfWWzTlx5akIw+al72mNsea1l0TYhGhx3jrgaDMD
IkvbWfGwS6Qm54pLNrDv8Yn78yO9TBujTZPHK89QaXHdPqLZEdYsDc4IxmQXnUz6xAHxIV5lNu+u
i7M0INSajc33/euZ4FYOxFAIIg17cbHsnngO/K1bcfbaGIiD2LlKB7PpCHKeJfd1S6pVMFoY5Tt0
ggI0V7R8yYvJZqqM8P8bn79GHqjEUHjRUrTu70O+NWWRH+DVALUjj9q3hRRjZvdAXiikHs97lmyG
217bDKAXLzksldTVzNdn7vuwRvWfruxKiuQqc3x6z9VYrxqQVhEy3+/8brt7i4cYrG4aE/dbsd9F
J+CkoOnOutBeRei7LopdJY4CyVdXfYOYk4xXTMpURDRnRrnRBp0g5qqHS1e4qGZDyIwhdmObO/AB
CPb+O0qfX62v+TUlqSUvI6Gst3OcrJBWpQEnaqZHTsGDzecHV+/nTc9NIimSFF0PtuVow8mX7lgX
djf0oXVmFFX/tHxpYI9Q/14dbZTamdpO6n4mFf78taFFOCr/ohM6oQuSNq5j8xjrpgZFRPekKptw
U/6knktc26aj0TWfVXXNQmNp/rVcqZUZGX6cERaW69+AN9MrsWz1PP1WC3nX+MnJ9woWTooslivY
QJDtfo84uINpjm+ZgNc3u1GLtXvE0q1wg8sEnhlK0YJYaizaEPDJESyecRCpCyu4JHXOpDDEZiu6
dbfX4pMtTnL+/esE2aQcFSXwacbFTn5ChW7E8uAxK6VKdve2mlQe0LNS3tYbWfParjp72HLo8kLJ
uFMaainSZ/ZS5UVhEuJnB0Ir/A4N990JYA8INRw3keHKpAs/xB3CoRcJ4kjpBfz0CtV86QiRHRM+
uIyzOx/Zy4AF0L+F7MtSFsTQgQyYbXaOWv58qv0RpsmCsu3Z2pZAADU/LzRxwU/+ESGehCFFCS1h
5i0gz7g1sPeR5bTLtKw+jHjfYoRQfBIViczMRL/klUsb+9MGQdbX8gNF974nR2UbZKQsMXLdE43o
X74JPTATmG4KlAxBeqdxWO4BuZRpaU5q+BRKFzFpYdhuzrb63TqPMYNQkoGFzdJ4QFdQ53nXX1y5
0ycIfwr6v7qG+NHGHne3MfP801UFogh/N89Pb6z9WnPhw4bhV0hx/up6cAT1CioGfdp90yBDwwWH
iaHl97f0/fbU0hk5E0soyYX+zer1RyWVRMedMRbaE090LOD4qVBK9Qe/HqmnkBzAK/0D++J7Mz6/
TB8ckicQCVACWIUWu8WWAZU8lz3exekgv5/UpLWzlHRHOQjv4oX8WrLI0/eT2w/osrGYWw+cHZmg
55HdeECwdsFyE1KIS7zQnbl8XhiM/9a40O2UadLYg/Qhdpo5ArNQ836XfEPAIPDTJIPEP+KThnB4
PltQJN9IFL+exAONnTJq/2NA/XDa+J7ZNWpW2Bjm6nyo+AaMT75i/NdW6wXKzr6w97hk96FTvpLI
Udza359JhtS5LfsxEMrBtpst6axVpp8YS5km5WB5NQiY5tC9I9JljykmZbIAnt4uGbsGn/VydxFK
SJZkTnxH8rsyXL3HTkfEGp7wDsQqJ1CbK9oT6jAc2UX14yDfBbusbw9JMcTKUNGWarHHk2CfdipB
KhGwIUkYordT/w16ancJpUgPAQdlnDoppvf1tJV+k+yZRxhTWa8wgAhLugarrinKBjRwM3NfzqdS
q8CLI2/5LZ3Ujh/ag53KHmkiX7/nEozZK69oO+gn9vNrwS8vG8SPzHzF2efYf8t+9Vl2ikIJRuEE
SvwnAcQewcYos1k+wc6dXVN/yhbaZIHO5KEOZ8GAv0QfUTtJ+HQXuLeQ8cnJxjMJoIraSka5JL4y
h1fHS9GFa2N0bkkDEPL6LohbnO5NmVPRXz4IlD/RHPV8waOCXsVgYF6S2lixqSGlBnvnFsiwVMji
XA2iO7O8Qd5cD3Y/4tZ5zH0VoexRJyvsR98PtZDLX5JducHhlL3PrBhmov0VL0827LJ2MnEBz2wx
cnYxFaslvCzIGaMrkdZMRkq7DKUZO59vEV6Op77mpqoQ7FMdnvLtTkaXGnoj/9iptqOpP1pRL74j
vgB1c2shYg+IzedxezJJszByXo04DwOJnaNuVRzgTt15S/BEG44VsqOmWFK8hNnXm6+9xgFJIFIM
a7gtC8PsLVqG88/lTtRzqIIL1dfw0yOa0AI6POniowj6/rZHNUZYT+NXJrNV/6PJzdnvHp3IgPHk
zyZdGbL1u/R27HvsQbor7yK17YJd5cxmA2pnm844xJCuUkYsX9VrqiegKcnNCop+QozC9z99Iiwx
JdqKxSTd1tXiJg7mvoBT4RTcr64V2OLEUU5obalc/Ng9ZmqPUZsvELfWtlLGmWicNF7o0j/VchzP
i2Z4Zpd7TjS6U+NiyevjmWygQYBV1OsWQ14D49T2mIs8ly92PGRYCcxa8bQanBfBxwtKGclYfPPl
0KgRAAz2zIipJm+7KvV83XKpUfDGVpZbloAzWRAUN17rGKBNr8WcED+qz/I0fdLsHMAlXJmn8suD
F6jWwWy7vKtEwZT0NHge0CltIkOROZZoonjVIdlo7UtH8WfQaAAPfJeEIeLlazzxGZmcl4+SHNpM
fx35y9eSRDrJPOEOprPrQ2XGndnejx1kBr8B7yhkI2Bqmwc5YJgFCClNFcyzbf+WceyNEIAbsxDj
gaqh7MAp6OiRRdELPxuYkg0aI1m1nqH1BTgmTs35RY01hgTLXE6q3tLRIKSDE4p2ZrDQkNlLl9vb
/iPLqP1R46hkP0jAfL2JOsfwisEN5kt1lFpmfbnTvGLFyfRTRdf0dBsXlMM9qsIiLcNK0lh3qZd5
2S6QaZg2tL0TtbWvtWipVXJVGLGv2+Bsvz8EXjZ8KmQ2M5kep0UmChlPp9Qyt5dtzFdtBunWFmv3
XpgKbfJYSDauMfcWtiroCAVaUkjXM6p7ZkcISk/ijcx9Rv74xaPGINUcCjGAR5UhCvXZ6L5+6QIn
NZdgEe+4f3r61LmAuMAu7jYwdFhH9iB5Vya7cg8BrBxRkMQGP+c692/cuVOWygPVZmThe6iGKIYp
srMJ69EHRbjVk9s0SxUTmIs4zgwjQzAY971FNn84fpsg74hgqqqp8p0aHtm39ZNtRSm7GOd6pz38
h7jf/zWJMJ8tu3PdnoS+mJqZYyVUn/gFAlON6u++iQF0hdlcfLylaxmBg/sLF7NHgWXJPT4hYXX9
adMQl0+lq5bpQUyuPbs6/hySXP755BNF+b/xLnHYr5ZElDQjPUFl6X6NPq4M5IfD2DKN+w/nGzg3
bQcK6QgrBFy5Ujca9hxGKYWb5dR1Osb/GHH/kht9LNRbdyEuEzY9Z4yJL3uHxKwlQSIn1hOsSpTB
ifHNe/nWb+dkvCT+t7Qwwfc0v36No7L57GmpL429E26dw1Gi3KjH7kWQZykpWu46agGecn18U4yn
I0sJQWzvQDWS1FhGvFafj3ggZ31GG1j4mcD4emYbRkGowN76afDSkakOtBvogbqPJ2TLdFje5G4H
SPmJ3IuzwWtVIB9iMwJTBtWCughzy3SNvXc5+I9vlWlBxqqHoVOaSPKFWEyoDflVbx9ZzWn20mUh
zZRnLAnWKmLAKfuDYK4DIaHamo7qdBKwQcXvFy2tIlCTuJlGeK/dInLkvykK5HGwVGzfRqmjglEc
k0ouavj9F7v9zGpKOjAYAF/kGrBbgPbLYveRYRgyQHczLEjl6hkkDGx10G3byqNY96LFQph0dzqx
OzPPygGAbIlLdcgzujikS+lywvmUaBBDGIRdvSEelx1Gx7NNp3Y5hM5HDMAwx6HdDRdoR1i0Sgkg
AlLGgYO4ud1VujhC00qjgzq8SZgO9jA5EtSyLF6KOXjNsoEDJQvmo4t2k5AUZA98YyuDADrQJmih
nkijzBuZ+jXkfA+P3ZOc95229ydwJ2ZMRXlkK74Cfh9TgOyLPgR5Oohun4IaELvj9T7reBgKNZJp
VpgHb/mJt1ChUiZUEYFCYSwwOaIciYwk0ESzXpDq3eRU9Sbp/RGksLAYbLyQVhWhVWG4SSJPa6Xm
Y7PULsTPQez0bc3z0qoyYYpv+etM06A3kA1HnmyowTNQ3VWlkX+1SFP/uU4W9GunbKXloZtoVTZK
tdeq1c4mmAwHYpdJqCjy6OiM10+VxC6Zwj1UUEjz/F7/S0QreZGlj7sG8bZ1N6+5e48apssCY6QB
49QvJZlej+uks/Qbp0OqQWPS0nCWKKFU9TczQ1bkBmvIS65SWfL69WA0MCDoJbrUNtBytt3/bUJm
LUoQ2VFFw+8COA73Iyr/5KW0oo2VtlrMmwkcSDds818hlu6zh1uzmfJUZ8kw95qNz/O2UDcPvdSg
1KzuAExLkpYAkAqwYXQnio13IfPTz/JBHwyJ7I0NJRswFKPGoeb8dSMdB3vX0hhR2tKzings9/ho
EctHr6v02tXza9Jx5cIrF3C4MW2hRCq5WVkxSgSt/8OZV/OyNdHu++Z9bdncS6bWKvtR2uCxrTNq
R2NZJVkpU+n88O80WgNeuhbEzLiB593C11h1XkQx31jpTUF+m1w7a84WjmGrmw+NarnIy2et4ltm
JxIAEZNuTStn8ol2DcPAD2Z0XIdR8uH3iswEoqlsdAwHYGTGiQKDzuMqrk7ZrSGd4KA9pA5al8iX
KfwpjoYjYIIoAFd0/4aoTiLOheW4cPpHRaHJ7Ol7SNoyQjgCeadz/E4P/YKiixfbwrFYdHDXBVne
cP2aI/9FwPB8zTS31ORKxmzf4ngMyhTmdr1kpL8dzVguO1AG/XKPt7i/x0NXjdqD33YQNgPMNh9z
fXrnCweZTGKtwzfltEglTJIRbDN4lOWfR5ofzs5mBkZb9kZ0s9AW4Uf3HOY5g3P8zErx2UWQQDo/
yVFZ34EyT9ejXMhpOYFKxpXG0x2zok3K/CBq6E44O6KrfXtEKYi0ol2PP3mFj24UDDpoef/h6bv0
NwTCTqTdBhGH668VpiIiDJxC3R6dV6PI5QUaSiDJ0evVctb2a0xoQRcSqLg8XVv1OPfZeZm8Kxw7
ySUcdKljq7diLzc2JkshV/lIduNQURVgMrMXbXf3eKBTDjnn68lMs2iAp3nmBw1i8AtxJEQ8j3jm
t1F0lNhJ6halLYOKchmq5hFZDtsPSyw7iRCEcfBoxYlpzdljcXQJaroDksJiW3bhkhvNfVu/xpJE
CUAeWtDbtACOMR9qN9NMsOWlVJ+GAFVf9mKhUHTJI3kck6FVYeXWrM9+fXjoan6EycfWBO1vQRLI
iOnnqysTADKvefuUYKS0CgffNEVBXQdI5kP73Brwn4pXfr2SWUpDZSrC+FdQkSS26YRAn5EbavCT
SIM0Q7P9EyqTF01l1Ruz9cr21OisEy0VWHoD9GNFkTNNEjr7/abLpF+H6ASDqTsGfGVTfmj1yHS/
P8NsX+rICaljS+O1m08v+0TN9fATIar2wriOGcFJ8cdNWg75fCMEG3UgYehzizZcSauv9dGbAcuX
2R9eyafJ0JAdmMIoCL95/VfcoJcv+AE87fD+Jsei2KRuhu8HIcSNQUOaNNmazX3ndRDYLDsYDMRo
AFplaiKVy/y1tkwNeiklqrkjJxcSF3i2iaSNpEv6y7UJaH/jwb3pniugTlyLAkWKic5fKe3rwK9w
Bortw2nWnrD1sDiH7seBh2YIj9Q6/mnjyBs95xaQuhxhe6RwX3upw2wcSsLUjTY9xQOFn61Y4MBG
3cD3Dgr8UN2/vepmUB6UPZ/Suymnq8vaT4BobJNImeYiHcVMJK+QBlcty7h+gstE/FSs+DtzQRv8
hC4vhU/89tVZAKtuJOXeygHjcOSgkD+xRWEhIGyiT36yl/7CJGUukS3AZLlXwSPmdRBJqtOSV1yY
0iNHWKUa9+b0EFJB+xnOf3+jdRW+o66R015dNgI7UMZE1AMJRTHV8RAcC5Qf+JO4Wnkw0P8llOlj
wUWSSm9P2FFcGFgWp6kHQtevgSmxlGdR4K9HYBOjWdc+EzY+uwcIsqDvYAkXbmd2C1wmn8szgu5L
h4Pxt/GXf+tDetDPw53OGzPvReT8Ky0QMcsRRHf4pcnbFR3R4AgBfseJJ8IDQvMh4fRsYOiweSYb
byNuBPKh3B2Lx8z7nkBhXDJoDJG+RQ+WGwX1dusD3yzYdI7nXq+QeyFvwYWV1mGJfY494h42xWgZ
Dv6OOE4XNfW/k4Pmjkuwdd0R2i+UgXGTWhJ8A4DkH3jS7OGxmIY68TJPWy3xImsKQgxu+YCj9Eoy
ZFRqSPMSzJgsE9rGfUutPe2SUunhK6qV73pNkFaIjmfm8tThQZXbEtgpNH+gR5qoZZEVGGdYwg9z
54G5YvIyTIhZWrq12+/Q2fWELlVL690Ieqbs2lslwntfqoKigXsePZO3NlfCHRhDivXKEcEjPokF
tpv2crd/gx7zScnAxhQbef8mbUA8qe4shJ5b/+KuX2TXLu3KPDMLvr41e0WHa3pHYimZZ2AhiJzK
XECrZFwHe6aPo/3HjOJR43IWuantQ99Is7doXnlDPLGhewvnpdXxJW2iASn+YhknbbVoLu3xLg3I
5SZms6vUH5Z7ErJNC+CvhsNy2arHL3fXwfP2ikRRX/KAFXEdd+jSDYIZQgAltVCF5NkAPexCunnG
IEzxGoEsjYtiQXZd0mV/rXw2/QAByLWV8CLp8S8XCU6UbE86KQNgRhjURCeiIcwHr9vuGOKJL83w
tO4urBm57st9e4o1w/sn8ohcWVZNsZqFe53heMLQdRpUQLIC+s2qgzRhxf2RdmO1W/4X0SwDuEW0
USyGP+DtvvrnaZpMddyyk2mdl1vbuDMu+mF+h0z3ctAXDM4sV7q+IllM825/KqTLuDD2/addovBB
kQEpyMDVkHCLyCzJkLw7JQcJIALZ55z626dd8+zgGwAQU2O3e2/+U++u0yCuFp6nwmT2Y7td+H8d
xJkrdcY7aKvmlhTqa+AQGMnlEPk/78wmGYw1eGbK8s/L0/gCfaRjQ++i94dNJwyZr/psCc7JbNTm
RCtVaIavjfmE+udusj68aKW0ZGa3UDhtQELWrv5JexjCvlinBHetgk0qdn3cD8jWPvV/Kd2CQTD8
tnWfdNRgx/H1fKFsYOvnswGfk68cJDcH5Us0/mrnvaTSjOcidj9E0OqEr9bBsPjp/i/DjVO7p0dT
T/F1ihHkPc56vxfw1MWH2kg3Q5zGvBr6wEyAkDrq7eKs929zVRPFIK+lioIzH2AALAWGHXm7uBcy
BhOlbyAAgvjnbEgFWcubo3mCMmPoinGvBXCf3/oms71PIJA+McsyCgsQ+RPdRwrhsFyZbp8UgUgb
fVZ3H4y6NGDLJEuzVWjYfRiekXbGWyqAkXN165vsS+6FPonV1R/SA3Qy9tLzrtbQj965r+sgmEPW
SMOLRcLT5sehKI4V0NyWyeJ/4KQSlEkqTs+zQQ4hho5JbB04a0wceNwjtnPM5Lk4eiDnIxWxGIXQ
kkJpGbiyBtIYl0/OrEyKXi5sxMcPo7OuctFwthsrY96KIJqrr/lgeaE+qeVTeFFcecZbfRT5gO3E
TIc7wOvK5Tgw9TtVqcZBtFcJHNSpDTzAaEMpJLrtLM8mTM6/z8ftUlTxPSoCRjXnVBMoxHPUPUFe
Zw1YoRxGpD8rkSrqd9EOoiBYFrZbN0C4QMs5vJHhohoNs04wDxgFFzZQs7lMl68f7/7AiNA4TH+r
3GXGxrGpS87wu2HuQPhsjJ5AEj9gfhOQd+6hQftvw1i0J7XluOiDsRID0svmxeYDIpja3NLwGvJF
iLVlvRxQ7jZiGpC4uoi5fzyKwWvRQeb2/WcaqxAx7j0odRP7xaXOwaFr3fCPh1mdzsW/GOaapW/o
GzdsAhmvdeiiS5L/7I8mcd14aYBjubtfmM7bntWWFZyU3ecC7Gotzz/QZOysd4Cg5cSJlT9syjY+
04QOOCV55NwVETHeTqF88PuDuGzSrwosRZAKXUi0rektocHu/8RujoLZ7zRHDC4GZE1yodGNNxCp
amOQ9B7SsfkcPc4FsY5sQ28FY9K9AIeGIkY4gtpDZDQxkNgoG8rYjydtd4N6HnIxF8PnA+RokMYx
dFwZryFr8sjVyR+GLbeOnVp8OMj/d2GOrd1hPv+siIZJx/9bHp82JwPV7Kp9d1LhEveiZgxUhChu
SgL1rr6cZaRFEqCQQfr0EqAdn3YlNclYkbqLvv9+v00VCPZ8Idt11hcz2HRiseFw8qF1LcZ16zgh
o0g5Writ8c+Jtn7oEu5KAn1j+zA+tU9ryb4Upzkw4mlmpsI9CtrVmS+9j1l6Q9tuE8Ql/WHUp665
a4G/ML0q/LVB9jIrEHxcfMYwrguwPhMN31fDXmOQTDf50qw8rSwLYsSUA6uCCc+Rlvkme2wbDSW0
88rRNwCAFWwxDCrttTmLs5+xslmR/jvfnWWf4HcdT+OFckoY/qFZ10Sv4NWlnUdA2JBqYTYtXCgu
HG+/Y+bVv3NXWOrKBqYn8OM4oqMdNLGClr0uSuuF/WHlisNhbPgXrBdmR5jpLwdaY51fE0z6XYP4
1YJdBMeMH/a8sMjRuRB48yZFro/ZHxCC1I+NFDiOpoW6deF7BcAvoZ+US5NTMUO7TBXO27nO3xm3
HPgq3kv45TX0HZcwTuxJ8ign5ixif/3L5rwAVA3jLZ0rpPtbqQPGnxlNuvzp9Yi7szX2J//jtnDS
2YIPwH8E6VeWoKS7+3zcAClgugQZwXMbXszpy/IqRWRWi8wycEItNOFLINvJbpyczJ5sSB80EQjy
OiFSQH8O50t9U1YfKSxIGTFUz2/cYFgBvtH7AA+wdCDsKuJ8wIwIoXq5zXTM34eb/hNtwQFc0A8P
g9mLvXKdxyEe1QGftsfHDPSAbCBMnF1hTN+GGu6e0pZRIPWGLmNY1bdesnPd1GqMlBa4MXpq0AKN
au1hpXtYOKYdErNXucCa9QQvDgLHp82Qf04LIpeuDTU8yuRTLBjyoeYnUS+N4Ed0tueCPtuhdkMa
U6NhGJDvrHWEGNceNgziwmkfWv6DN9hz2+sVnapaTiexMapN9a8OqREHrhhBzzOuJ1jSJq3KfS32
nuPNur4f9cEvY0MLkRB6zBEGODXGDjb86T/8YjMNhadi3+/Z/zEUo+tiIa+MZhXNj/vIuVDzcwwv
yhlW1GC2hVtdO0TvnBI8wOI0k8UOZcWdbs5BMc0kkddqlGncDA0D+hL2y2TyOJLkMyS6ixhEdbRg
NqnQ7YVwrNpfqT0pUa9fRVmgLgwaqh91JZkUPDqSq7vh8djfj9cbUvPkrG33Vl45bPi0JG2brL7q
dZTuUgmzLXR2S9Tuja/4GfgjkhgQBVc6fd1seQJDc3zvx1forloUTHfz7Bmurvz+OesRkZKYlE1v
cTIVTDZ0sjcGkaPzyK5NBxfECR8H6sWkgaidYObiaEQ8JaGFgwowKhQqYVLWOdd4UHwTFdng+zCI
+ce7Zx6Du57rbMiKHT2/wLld9WviP0VZKDj/6YPL1f+fC8wuA+bAekzPKOy06KUXwYR/kL49mcP1
Ikc8Jy7ON3ChuBsj2Q8xOtcp0yQyfUEI8DAHdneaYkHHgYkR7jrgkEY4hiBdrLtyfPW4UnI8c9NY
OEnlx8DSOmiJOR0aJuW+TC75gMwW9pg04VKoButG1RehvKFroec/q0rjttpMdJP4PfWgE1dJ+mbj
+L8vzkB9dK0QBg/3P5NJ7ApMQBwxBi3E8e9YVOH91a+1YM5ZHpcfNPYePZ8gPDS6Mi1Ft4pa85nt
mZoySY7N/JXn3+Le5LSBfHtpHnVwu96WD7zmYgopxnA0JSTTwQptnF6EjRI4ltCnHRdgENQSB6f+
H1qKYsQMWY0DUqQbTzOmSMyEc/2yQOyuLAYfDtx+7sGF02C4J8fxs+5+bgJlpNnhmlP87aZY2XBb
Xr8yxkpxPP3dVvjICjf2sPe1Ap+NJ6MXsAldNmAdnhmjuUwtMry/Ptlbc/Mh967uebhgm3Y47Apz
68gUucmacB/akvuRhVXce3z1ChTNbbEGgdQiWe390RyucoHh8pxIHwhMKQcZOqbZroSyhB4zc+9b
W1I97JA1PD+pf9H+N8WeX9dA+ZmwqGBPwi+HyIXIRAe8yb71djXyatqsTsUbCP2J/V1/Rb4Pbvp0
vNExeXOJ0H1HVxR+ER2nhbrzteE6IK7JCucECYGm0wBrDA88/hNl5jj9Ijk1E+AkKM8BZImlBCwP
AI9wPsNKdJdSSXMKvK3YbOL+/OX2ZG00ZUvvvPELozXKQGKmNA8HJsKNs+QGykb8LrO9sTGV5k0K
XrahKPr1twtcN/QqrlR8AbSU5tyvUZN3OqG4GtkoRIkRe8kooQ3cHovlNApqNFhfPmCHQicdX1qX
DKRYG4e5BGVkTXdzC5e2cNCTxQbKLa0ah+rkl+CesY5/Y3cj5z93e1KINdZtemlZBJIEC5uhzxGv
iitzQrPmNiKqUJ8gNBP9s8U6bdondrvgs5RbfSDLiGosGQklT/wxyg/H4pXaJF0SjYxvYPQ2ymRG
XQiFqkM9pA1u4xENZl2XcxJ8MB+BodfnX+yp64eOQNeInkAXfP3GR0fnR5630ToTrGqNSxvkNeK2
ozdaTw1O57q61zSWsRi4RMWQ12qVYDpKpJzaUpsG3X2/6t0WR132p3EotN5abNCKnlXPuxKRq0DR
ARcWszSV8ijq3Vlz3V/UaOiLWLOPvH18aSl5S2IBoc6H2h12AD6jeCrR8Y4HY/BzGv7mHTB0x6Lb
BSklBR4Js+iDLVvd+cv6AqDMuTIMFZSomPyEHAOPkWvYvcVUMVlFcWClp294l20pK6iNywOtgAxh
we1A8GW2fqaWhORHXxJ1c1AO7PVGyD0qMiFM4bNPqdZzmXeAWWRcL6XWAmp4084wc2mJQjQU80gt
w1JGQ3Q7f93RyVHSikE98avbV6KMIi/iEjSqtgumK5NGEam4Vk5gj4Yyw2jawK9NbCZfX1wiB8AR
YUwHTXlZ52piHLL2UVDlcIPB+ztsBnqNBo0UfW7f5PTDiUgPZC8hLuB3z81uBW0tNb2fIoCGDtom
Dc0MgqruTQXi3JJ1LkppcYEzEr/MzGkzMC4zUn0r/HSGC3t5OsMqVwzv0W/jRRxtsa3Rc428+D+Y
7f2HFwzOZmAiDIT/IAbylopzdTDd5G1eLcIvzLym1IANyfX7rFuPcFFahFWu86djvBlOTGycLi+j
LiuScU4mDftgcmr/zEufqKa8bTNlVsiO5J9ZtIFnjiEzW+CGzDaCp+j/T4NodDhipebY8/oTGonr
iQU6e/HI5CTHmm1P4ZB3FUKtkd9UVvyS+2tpdgeIc/xBABu6hLDFZ4jjZtPK6RvkL1Jlw9kQeEGG
0tt4rIKo/WvsQMSKuvh1evfHWY7KMURxWd30bDfBjJGvQrfqamn8WFruUH7K+G6SZKFWrP82Scp0
gOpjopEHsBb4bZrmP6PDTyY3yPBO2lNirLvJhYhaiEex+9e1ly6R3RGICUEYyNu9BRIS18eL9i8V
/wbqpp4p8s3hICU7nWGr9fTKQM4Ylqmxa29IFYgV7OJ8decaWohaTs60N2iqmjq60dqRFx+VdqFk
onY0fp26iIJKUw5SUaTfgxnVhfC4EoQy+/CSydIl0unMA1D5mO4tw7EVjnWwnB9OY9f0nycp1l03
pxTR301QZ2xc1L7ek8wnS1VcB1db9zOs+YaE9Wy0vtvRLQHZ8i1Q1TYHG7UAdJt960cfC5Bdk38a
R5IOr+ibmc/oSL5sYY37IziRDvgYzAopUhXL1XWglg+fEuSGWNbIWjRTz+TTL51i8TxNxB1aaUfB
9Q4lwlxPtoWqrhWRrkjtTvTZUJBZhLKrTA+4LeHtziIIIKUbUTcSYxH12zRa8H8ABNeEvGFQbOud
61JAjfHPvGTIwaimwh6RxYvUJyjaJQ1rGZ3AHYc4YOQazglwlrTuooXGg3Av1VSKDUxFAAVsAbB/
1ZTOwXRkKcdRvWAnF8yjskXZ3wPXqQEpGuYBYnA17Zf56SNyIkUwdu95XdpsHkuhkbpIkqXw34jk
xEUUy4dTx5yqqpWRgVZVg3USyN7mySyEHUbrZwINcJZfgCEMpvBRqt6bcrGpcY1cG0E4RqD89mr8
eSFhOUvCimMGBy16GaYZ8jFyY0iBODF7n8lv9skJY0t7n8RDEQZU3kMS0uSX/5sfZ5bRwkOW5gm9
O1mmpE2YIabdc6jqqmWH0Iu+wi6GfI9WgOxyH1JYJ791jQT7/8/aI/Al5+nTIPWczUqTklmu97Yj
HcnSvvht5/DdkanyNsK25xDqR6lUYAsGtERrV96JlYoBtJn4p9GJgshoWOtJXnglBAj2ETwWqn4p
R+k2xVS7HtdbT/oENUq+DDtVYPm9chL8KM6aM3wpfXlgO+EMEe7aTUKqo7XrikyDyx/kLcPo1KWU
10K/VazCgPumxxfquFrOV472GM+d7NWJGCjyoApTjPzm4YvqQ/7HQ3gNNKOCjksoYBKAiaJ0aIly
Lqv8WCt7YbYd05+ozU9ZMCvBoEI65fxDpUvixesrvrFbrZfFo4uiD9EDougDweUFvE5/jCKzARWK
UMwIFLQMud3NUJ2ypS2IcDQpPB1T+6+vaiEG3ChF6iVfxO/cehlbGPJeeEQdYSssHp2o+8+d/Woh
hwRziWtTzdu+TK08VMbrm6SUA2e+ZWdcy1YyGaSNVDkoBj6egbyDY6BeTPNHe3uuBigtjVMxHnu6
ZP1Ow5TmLc+62DVeqEwGIyHXdYlxbKhoXaFt82aRY6VIULYIyHABomgl+IM3ePB3dB17ADNwKJVi
YMnfT8blpeRdBKLz6YvXfGimBStLWmPQpoWj682gtJ6FcLyHb+JuWjIB2WsNJwufmkEjlUCoiaWb
tWid8b5Ia7PxQZ/HbymVhsQWhKNaCV6rDauCikaIm/Tf90c1Bu0Jhg89WAq0LPFblYFngE+yHfvk
toRiBV6550MIuSj9FQWa2LozbTYhfMynclopyHqgz7d6GAFNhfWHrFToJv/LxXWfaKGDpOyk5FZ6
mhjfCXZGjmFG8hJ7ijObSMI/zUZ44RjGk25GEvB7QpnKdfQ6Dasgx3zY104sVXeS5knDQaT4QBl5
aTiZx3Twwl1upMkSv9fYWbXb8zVvWi5p/p7vtu1OlxiGBOW4nDVKHVXI9zLf15iB4i/TYVj5+NiB
gFN70PSPQWZ4QGIznCUAkmdYH8nF7q18CLlgwdC0m9DBZqWy3wBEULNKroa57tC9OHBsSRUdo9yw
OqOL3INqZTHHNlad1Mm+O08INjuYuPN9+gmghQ5IwmguwSLzknOOXu8tX9PaRVuA1BCDFlQCBPaJ
FphkKPcOjUXO7SNBT7Qv3VnuErvHDR0Zh4xwSqKV86fk2d5Gt/ovAnhBnQJPMMC8q0golY+UkB06
L8GixjGFh00cA8NIblH/LYao/JtLLuhRkplZLOp1OB/znka5WcVzM/GaqeRGa/CvXWQ9Rbm2t2Tg
zqPj7Oo1cT3TnW9pmvbcF/8vmjnPds+yd4Jn6PG58uFRI4EywFJ3Cm2LPAqhAGnIlHqEC9Sa5xt1
xgI3Fdv1/Hy2ur1aPtAQMiF62jGlVa+qflZjcGZxMZxxEq3XmaNd3zOLjOoC1yK/+UjbGRg/EWgE
1fKyOE6HndH/LXWAdCgT7+WRfIBSheRoxf4TeAusVz3uqqCnBdefKfECr6vuUFL8rXH4F/43Qu/Z
s99QZi1xWRF46dgsRBwJ7czH4t4hmjplFLjQFyiSI0/+VPo5iCKyeYoyrud+BqE3BiQYiCe6AOR9
niQ8EhOkWmBwoPT3xOcRZBjeT3vUAdkiHthRsuajgZhOls5tnFvN1fwzkLbzDcDxqYGV5jHckx9K
lTx9Wzs3kLa5BdSgZzLysLnc3b7PUOUMhHdjA90ha/A5hpPpEhWCe/F8dDkbWEr5T+WPgUiKQ8jm
/VmZlGdRKOhCZ8F5ECxvVo3SFEFj+mYvexk7Oh3YbNV8MmPn98O8CvAE3NjlIMfL7N+E6RCZjAod
epka0jjxhjbYzvMyZfgZ3mnKv+ju+geuIxDdSw+Ns6jtVPQEOcHGXkieb/+Mhj4U3fKbgWTQf+H7
Vrj9EH9RObWub2HAsq3Uz+ucchCLq0Moj/lEvcwBwkPkQG3o+twiqt9SVx8j71TJ78Rx6JjAOH/t
sdOMt9/k/o0dsXCOXm74Uy2xtITeqTewdW236Vdlf2NhbvvTS96SCGEV/H7yBE0VoCosKiXMNV4B
SaC8LOsdBjdUdHM9DppyOAxf4sFDMNWM2gE+qG048R2jS1BvpXpakkqkv9rtj4Zqgpf6xZlvvlIa
511TJXOmVkw7+gSwJyssmm/uwPaMcAVpVlonKAgTpAWeP7KIHN9dUQ3cBnd7Z64SYbwoXvWuGC94
uO33CDXtUOhi5yYd19X4B4NjWJ3JeV4IVT0a+5cZzCL9uJmuoPDwrBl8d+aJEfV7O2jeGu6dfYSL
Yz2yRIRJBp14VikXT4QJDF2DHJzx7MWBP2vfN3RvhFDKAOt4sUXCrz3CT3786ClWBCvXqXkXlByK
KUV3m5RYgRy+YH8jRU2OIj2Pnvl+tQ/1fLWuX0/3ETecaHQaohi/zENWliNN8lm4RlApCV1209sa
ovq7sZc/YHBvVjPBH87pRLrSXz/j0tXeDi2/QP7qqMH/uxjVNIuTgeWnFmEuOL9xULKkn2fggl9G
p0DyMion17YQnlEJxzNxVK3gT+r+TwDprZm3iL1nddVC71FXXLOiJEShFHvMxsXyHsIVGq4jAbEj
t6XvVxXZWZkLISTtxLDJRVDQwcyrOR8TBiMfzkQWFWyt+fE+rz0GD+Ea4VleTd8w3mZvr0SYL3We
apbCKanWUfH8dZUJ0JGveGqk22238cFA7FrHhzjQeJalq/nMNwp4taEbcpn6rRhunPBWj7IPXXFN
YX01IjqgeFlzRggii+29IwHr+dgsurwSLiJ0E4B2qgz1Pg1FK75kglWzS3nYflXj+ARmNtzaqjXi
3+zcOwv5uQLwIfPAGynGgowBHvobVB0hrgIMaPpUXax5dpbhxbx2HpavTZC6ga3WE0H+W+KIalWX
ayqRW/aiROS4RqrpwrtAr5cBNybNJrGmwvTi+BNcsg/SpElYGej/dxK9gC3RmGiEsJyT/kHrsJoj
2O6dKxOPgcTaKBADbHPtYh/gKveDYl4nzI2xwY3pGXdUSQWiD8zLDthCUPTrDahOGT42JM+z3UKC
qe0jpQXHfi7eID8mHIJsUkmqq+ernUMCrE5zdfYIRZk3jGE5bDrBSjBSclXq3JXtcbNLVZhS78cb
DUod2oPV4g8bsdiYA2jlvMlkhTjjFoUdVEroBhpx41jM8SIyv/O0rsJ2oI2xHmXyJkovT7No9xKs
PS7EPOP1vk6ZTo6ZfxdZHHj84F9d89O+wrNzwfENxPjAht8yOW1D5Kd8yrxx+YCZlZ8WX2AqdK7E
VR5z9N25iHBn9hNvo430PoOfGVvtBviaNLQ5c7ytQaO88pUOL8i5BhAmbgE0YlzSZdcksr7mS+jA
PsgepkvyWJTQl02XXghlnSmfXH8MH2bDJHEjdON50LGon64IaO8FaN0qXEwiBnphx5+D2LMQRb3q
/6zaFlemdlX88KtoY0/vreaNJ/5WgXWoUW9UK4Q2wruxao6n6s/LurQXbnUEcYlKQsGebiszedpe
xVwporXQoXnfLVGeEN0OpVgFySbGt21K1fF6vWroDO8EE/IA/y5fTMMGlaxFydgGej6g7iRIX36R
9jMdHXDdRvUqLX36FoPXRcmHx6D/sFxbDezBSHHb8N3lnjVC2IzXVpiORoAzEQPBQPLdKAly+S21
k4nyYqC0lbx1N1xTCVgoWL7lOCV+Gt2diAJ5GHOn5irQ0IuP1u8jXbsRHmoLNZCAdnMq8pE7ihSE
gf/NWVrrZqjfaHs6Vwt1kjEA7mHO9Ru7hMqyF2aTBFHyuJXSaFnFsx5rhtqT+bxDuFw4G/BkuERD
DvYE5BcHfOdo1AIJwzsUrmCfeusq9p1t+C5SKm6nkyN2mD6a+PTZ1u0pca+JQUvNK6PJVlDxKPDP
y0P3Mv5gJd5HOLmI3WhD86hFp/+Vlm8vznaPUc+ps1eY2/2gdfT+qQB0f3+DkWrDD45QopmLTwqL
LOwXLuZj7mA4eR/sWdGlS7SDSMU5wrxn8OP2G/8fGSLmGMVcyfZVIJmZ0B7M1T5sQK9+eVx++dJw
c2GFF57dcsuPTW//Rhzw9AZsW1e68WgZnVj75ifmrJTieM2cHnkJmMMRwCJGBzHr0PxSMOWw8KfF
DLFOm2XdZenqKdYC//iIFaEPfkyKhYlffHsZ31RdgQaMJk4agF1Le0TXOhobdxalq9QSG5BDPfJp
jefd/dZed/n+hGrTUpe1obxXrGNZ5YD7JGnAdCLYLhkAyKk/6ycoVfRNlcRiB1fwKo44Ou6YrOFk
BmAQbnADdFPyzmciM0okKsKfqyHVWnwlBxMX1elWp/NruysTK1BAZOfotqI58QSky3Au/5JYTtWY
9kDGWEo6aOuOt6IIHHR2iCgV/CLwT6m7jm93SwnaG/DI1tZXWVgRd8GZ/VjmvLRWVx8aktd7Lqs/
t4yqZanKzKie+4FjOO0RjLL8i/KOD8sNjm9IfnzaDe8YjytbYtXweKCHvRuMnlqsjoUFCECp7ws5
5n7sdl0YDgS4CMrRAeblRMNGXcXblMK7NlpSyX1wfbv0DMbY298iNNYnNzNUIon3Hb3JAzCpWWy4
6BOA2ZqibKsRybe8peI1ArhQzsw8M2zytZWDw3J/mimyD8c6YYpr+m1TLyoJ+DF1aUcS1vSYhSBp
LIAZB/62+Ln8hPAH2JvCCkLPEG632jIG4gkR6Qo8yQRZsPxQnVVIzpwmgn6seHbYTAmJfgMSCMPn
WS0cgRTW8ePio+MT1EWX9J7efLfQ+F8ny+VH5FK0SHLcKipACWXHvqZ/6XAS7CaMhwy5Jh9JY1cZ
Isv91OgzQ8yvHajCLICBQSswgSlhWvFpQwE1TTvZprBkJbzy7piS7RUbd7la4Dx74FrDil0NFMu5
vcYNd7O1TgSKp8OLt+XFkraMKUz6rHDYbjAeQ8NVDUqLHr7ZpwQr6TFfz3FShn4wCvoI1ZC7fkxZ
HN3nmcOpAaGbjlwPC41OxfTLgXE1BlkvboQgRdnycuWjlUyCr9LUxNGRM9Zl+3gIBLqSyN62XveR
OcDiUHY4a1Nw4X3YEPSP4Y1THCebA1MMXdrsB+ymeHTbBJMLhIzz0zvGyhM0aM7AD0fEPX8u/AiT
bStxV0ih43JyQDBl96xtZglR1N1p17CJYmCcWxE8t44XNj69ZQetMwODJuTMm3jBtltGXKdMAOjY
BN040w+sRjoctthwTiGEyiFlVlRa74XnEDbwuS4qVjBOy4n3YR6ZBnrOCAFx256HOcvygMnIr5RA
r/OInZ9kSe02lpnI3z4ZCEe+XZgH/wdBrKAjRyuYk3i9Oq+MCJ8/dpRzTGIZ1z4HoxRPsAcoZ008
bI6XfQJCwryJD0rQ2dvv7PsQfUz+WqAvk7LSYmsvWEVwS5OVbe/WDc3AWlEcrUZ9rYoLz7bK5su0
qd4NkqFrYL9hhP5+Hlo2NR4tUDDxYDhxAQNphhtSuq64s9ef730UxpUvnnMbSN7tQx7mLLesEYtH
pBbmnQPOaN4Ix+fllQzTW+4nSS7375F+biwHkjhZ7H+MIqx0HigxhE77ZChC0knIIw4B1OYaQo+v
l6hztXKnElA47kmufkyinpiW+iyx2dT12+jqf0ZRqAngKppD/tzEMpiKB7JsFfna3whlpHDLZgnB
nXADs5CESizoJaF/tKdjRfYjQ3GA7POczYpkWyTssOlByGcxR/pAl2oieO5M7sYpLszwkAiW9KVB
OxVyb5cB16A9Xz5fvm+Wbri3SwTWOOQgqqoSV5/DxBcnB752JS9XmP8Tc3LJbJhLW2tUBfI6H3Sg
JSJsJ7byK4weI6PSqoV/Mng8rb8oxhatF/tZ+Bt+0mHi9yaT9E8MD759d6qQYQIjgj2DKLpdHw+X
wvg6510gbc0sO+6hA232qMf/6N+Mzfq4LjD2uY97xeUN9vKCG81N0RH4Png4lPpCCTmsickjOsVH
gy0T+mpwuCRofHg7e6UjwrnqRLPERAabD3spjpm3uopoeJR6bpYd+TFKWjlTNnm3Fn7b6AGzWkZ9
HwHwnHMNSV+vBvajAjfJ+Iy1NexHnOMANGYPqvLhWF2QA603Gdf2+nJdGx/DR1IEL4W2xtQ54k1n
c3xs//ptq5DydqWIICzwEPl7IIj4KLfA8iSHt6nuDgZG/98y8SyNjKM654V3GUN2GLYtM5SkPB/t
S9J4bOfIrGuhPaAWDd1AgN+hmL0I3lDt7Us2zQuGirpMCTV+7qWFYS1tswF5nFGKKSVCq8HgJ76n
d62EX751eJ2XYKdpIp9/KB7CXQtsaWuJnI6mtxgrDBnwnbK/LEMFN1ZSFs9vYKiOnF/2Fxr7pnNZ
6ae5hA2rwGbK0Xt7xsqxu5O/D5ij7dj0tgYaP0t0F9fi7XFYh/7JyoyZWSSopdK5AyJopYaRW3OS
7fLVSob/C3CL0kqq3LSfT2RVT+oa7e6W3zsvR66nV7U959ofmeQhofs3o1ZIX4XxARSYwYtKsrRG
OnBSvYgwP7bQTCXCDiYdeSAISrERGIodG/b8Yq0p2RB8tduFDYZ29eO2ie1F9KhUeHX56gg00zgU
130BF3BkzojVAtVOKaH+WniJo9S5VwdFpCZZqsh/fLYztkAlbNOk8XEqPl00LVPlDku8ecSkYC0i
D+4e9sTXJhsksvlauJv6cXna6Z9A7Y15MqUXC7Z/J2Wh4eVL172HvBHJueHI+NcGsD8Ib0qGaaOO
oGd2GEqsDQZgB7Wd0bPjOrE7Sb6d+odrABstt4TO8r37cwZNeeHkjZP0FcxMsjEmzHt8yewF4Puk
Dx7DO5CF2tMmWI66LZj6y9YeoscmGuYOpkdIkwqmG1+UxWK7pROJj0D6hsUwtX087QT42frPG+WW
L68lUJgjNTbNYFZzFnTu0FKYDmYTslgWDJcopI3CcREdTBir5mLOLZ2K9Eat8SUP9HNlUqyMtUFx
PTWNZcwoAQHVUb1SYaZZgQfk5T85FKg1YK91ORarr3IT4WyeDEGilbGJFOcQA9BJPe7yiL09kA5+
HL2mN81DTbGLVR/m4VdFQX03kh0Sk7ZIWw0kjZtOumSYFgz+YhCMPAJmhh2nZNoTSDp3UwFFTx9M
r5W6HCMmEYGXpV5u87VY2wE6j+uZj14wDgyxFNMm7Z0M9mgLBezOEMpNxUlGFcFX0pSPD5zL84C5
QUBNVVFekbRW9SoTIucoMjcVQPDgKspGgAasIbpJXyXRsEc2Vq9PcY31RzARYOjf5bCejL5OmSrH
zIxyoH1KAR+dGFZogc5uqVJ+oVTtONF9YfHQTv3CW/qkfROug+mOWR7wHKoyyO76vTkYRT6s5Xmb
3dwdIvjCd6qgJ7KhK0VhNj9TmOLn9OpP80Fh1h9pujeR2Gw+hfUf/iGIatretCuOxnICfrK5KAJe
8pdpqVtEVz9ljcSaJlqXIFw5FSAv0ydpGlB9wtX6R1frkLrebOc/+y2yvOlNEUH8rK02PQ2S7j/l
D3lUXKpz9kue05gGo+c65do4rWzjr5rrMfqNrtLsdPgdttYDIKuJh3F1cly3h1XcwGD8dgZKpUfQ
tg0brzuUBlGLnsTBSGx00jnDzOpxphyEMDdpGcB8l8sbW8GpsVEwB7Oyl7naQpPMYowQFzotv+nL
dwe3I4aL3hOknUZxpDAlVVwRonIiQ/6AIjMNv+WBuXC10Feu1NM2tXHHv3gJcjPKwi2IUCvYz+YQ
pfqrn2z36AvcXElZvGeFsLjWzlH2q2y3jR413RzM9ux2TYEJHTp+tiIl74fEx7hk3157isqVRTT+
8CV2hjdNVKmCwGr4HPP9/8iEmB+mBDlS4q8//SUn2dvfvfjpHoymkETqEJUSx0CCUGoxJSkN0I36
l6qBy4QkdoYaur1kmidpcNUWQj7B8sK5W3YxncIomIzgySeKeA6sYCg/4quHxiO8lEx6qHKX1RuI
9xmA9VPJ9g912PXFeV6LKTd/hiieDl82vEc/1G2UiIQ6K1q+z+J3CUpOBAYZmN2j1+GK75ilxecE
dy9GQ6jtzeBhRwymm+JYuluHTPlTzrHehVMyGFzSyJJSF8C0OotTMULyb9aQR1o5Ogkf/I+PIai+
aLUP4BXxlo1ueG04XI9hivAJZwb3Lm4h3V13Y9bM3RL06lQvNjYIc0AT76dtak/c0lbMx6DP9+d3
93wmAG65SbzRL9r6t5EIPLWmcXqtWUsaP4MRX8wKW5lZ5n6o5xm9wnDVzgV7hlOyG1ECKjDr+hX2
2ALN3ZdOrXuBShU7ALRF0MVxPrBzFzm9ywsjB9Bvn7kKaTx/GTf7EDV/+dw1IHmie+dEAPtqz6Ro
pNsZDS58No31rDtw3lIMKlb5ygvxB+yWtqruou3UFhkfUYO+r9/fJYcY0aXvx/z195VXyUSxafqd
GEwhE803frMDDf3NFzspP6aDh1sjVmcoz4nM+gz0A5R221HjsUVukF6zOQdUBP8+/nGhGqLSWQh9
iFKRgez+5MoQjkpNCk7F0RQFJ44eknxqbL8Ukn/VKmC4up19jTvynNjeuTKEVuu5U+NlRe88bk29
wP759yLGkXJk/WHUgza0SAT+ChpPw4KIzsoZ5eGXMhg/MpexZuNVP+poHwP8QS1ja0EzuIvsPaKd
IlXF4VClwmkgP2L7+3mTdYb8JTJjCdtd6hR6TcVDccY7NmFb+lTeoIUzlB2XJ1JtwDZ7oWc6HPAj
nUJC3sDG0QQuNMdyIJA3vZ2QI5JxhrihQkSUHRf50Fi3vUm4xgoTF57AYqAre4JMcsonGjss8oA0
8wy4pqSFr4Gvn4LwE814waSPIarXXxgZCCQn/7/zFB9O7oaXfEtdvt6hnsfiG9so3os+YKJCUr3i
UdgdF+rBM6FOIFyneCNtr79htYN5WrJNvWvxe/8NgT4HyAZPU62IJWQJMmEJr26T+j55Qnoeu0g6
+daiwT4EHaP2Rw0mslRFXrzDAmk4xj6Ae9JbSkLIG0HGuKk6npvYtRZIGDiUUtLijiRBMBgFEP45
9wyv8Yn8A2rxy5L0MvHRj8EDRkQsnUhbBx+y22F3xZZ7uELLrO052B/4pzPSiuVLLWzSxpAFCbvY
sylz2TKYa9iDq09YHiH4t7EnJH4Y7OjynZL33gshFTOi2pCnezECO8XBYttCsx8jrnAP+SyjRb8Q
ZWzfjEXkCghS3LhAWaYTcT7y4JvRWUQ02lNZARu8nJUMmUEMZ6Ucz+t0JtxgkzhkyJffU3NJ2irs
MqlrsHqThTQEyE0+tKRhMolLJmrSasdDa21p9gY9ufv1FFlNQJXEsNfG8/P0KM8i+T5CXqK9NmQ1
d0pftq83jljNsLQ/Yk0Qlt6nX3fF4osJlfBQe3OMfVWh51+eQ8wti3L7zS1ROdvMqqYB9C5srFah
+3NbxklUICe0segUlCnPEfer0gT/uVJ0cv9TyOQcBBNEZ+uHp1bRmVpRf0FfJ/TeRp3OVS7WcU+8
2r+JhWeZb+CgtcpDtEUJWqX9Hbq8XS2tfQqhEEgAlEHDd8sAGaN97l3J5WE5M0T7fkNNd4toyaJQ
Q0UJURsBrB+yHHocF2jNKt4X3k8DQxdkiTwzh6AXOCE97tQC/5qX+pceFknrA31MQYLczBZTEvy6
adsOvk3+K2/nxnshmbSdAbBpXfxuQub6AuxRtrFnkZbBtyz4LmwXSr6Bp7zLWEeNTGDMVzAj+Iky
NNdDlOuiSDNrXnH/peKNG+gXga0ia4kM/WC8wmNfL6fbVvOVHV4WdjlrsWlT5MF3+00OSnKH9u4n
YMkefmp7X/llO9BxsjzF2ZUxbV6kxuOdseq299NWmank2kTt9fpNzn1kZ/ww6BYiynCUGSRK8pOQ
s0yHsbc3SvUzZPdu4ToqrjVGSD8l8BYhXubB0rrS2twiAgtzqOKWS3+qbCBRI1bcBjtPrLxAf3Ch
Kc6Bm8zE/SiwwZWpwMDm2EZH7ah/HZ4zh4Rdx4Tpu10hT8T2kRXA8rQoS2gL92zgCQ66t0YJ3Dko
3rLyArQqYKTvx7uasfUUKZOewJ9/ix8Gmm0c6sI/Kf5Yd1kWl2mYC69HQGnLOXZIyT2ssBt3mgqW
5GB2YO+Uz07BOiEe3jCk1D3aKsw/1TkXk4SlUdKFN9UZmqoTYIsEV0aGFJxvS0Q/UzaiGsRSUvAx
rdCe7baYIprDJ/KR4w/8ic77EWGh8f6L4EpYVQALUwM0I29JjEYiJoEEgxwTtDwLem1Wd40MhPbp
uW63hvHBVpulb0//U/a0WsLLXyfWHEXSlFQQGbnL4WkKF3SUwHAc6T6c8kY3TpfQEr7BQFBFTjJ7
TFY3JiYQOKh9sgiGHFI7J/q6+/K4bkRL3jQrX/uWECr3wrcEIwX3tzuSJGgoFu2mqkDu8Df0NmtG
q+IWtTkwoduu7m2gokVqsI6hzpkRqHKDM75hP3oeHGsmypk6EeFPp4GzljoPInvx69FZCBA5hkFv
oQ9ulu+bSxDYE/Ny0EIAoBkXzRAVdBWxT9NvHx1SVLrjqh2TMVz5HlUZ49Ml8v0F+2T5yE1nYhrl
4ICY/gIWBK2YizR8VxE4BO6R7+nR1jLHAKZLzS0if9GBV1W4gRrN3XsgnYVEWfLZV1Q8+79WGLzN
yYmPyC9So3RAGOd1R8NCxtwYpWuNiHmh65g/6x/k0jP2FmjZWpiEe+Y3U7K0WMHIonanBVUucvIt
J6yolunLHky0RrdjkHxw7idQGvgPpn8rd4aeRon0f+qDhsi3WsqnZ/bd0C0XeTrqlFSkkHMPMLVP
5WWAsJCts2nlDnW9TDxRLccIL3S/m0GEapMtqkMjmZsJbGfVrwAA6kMdyY9WoaRWDvrt222sGN6O
E4vHt9n1CyWg6WWeGdRO7Iy/eKerHVpXXQT8jEj+rUOyFlKD/cC/sgb/r2cxJBSjrZE6ec3gE5ar
qc/HGpRuRWG/yF5XvTE6YE8diE8q8qtB7siDRD+jZKM6udOpfU0ba9Z05KEo0PhImOODjQ8khMIQ
6/knRuBd/WZC6q+bZkOHOvlpk6lP1/JpQI+jRoDzGMTKvVa+axp0UbGnv3RT8V9I1gQWFELKuKVP
1hCB2z74sf96uscBl7IYFmxwqLUa8fQT9EbhxYhyaboSCE6xAH7h6uhCKGwI6BH10hgDZO088jVa
RXFLJZUa0TkwbL4MVzRGdNvhq/opfDyJbRF+Ty0Qzu6ffFjpf3tSqaUUdmXegw73t/l2/BWzEM+x
jPVaAZ/zHfyaUoJGXD1AlchZmfbuSrWGgJCd9yAAyNo4DQejMGYsisrPgOGTWy4UFdw4uC5uwmfG
DJp/xybeJSZNK0lUV4InRCSCSKjuG2Nh8LzY93jsCAoenpRIKKwMUfsyyGUFP7XPA6q/EICx6e1X
F16lyi7jRysq+7lrFCkhALnlEP+wqXzauGU5+j7TsXUaUeqytdsi+VlUI3+QfHJ8MvIHS85cjyHh
kqJcRaWWqc0iXrg36EACYIfn6Q9Gp9TnXtLxz/tUMN5jxqBDrLUhr6ASNSErgpoz4Cptn33XgAHA
p2Gp2VVidnZ1DN+UQ2Dxf0/MymVH/U8ClusDrteCTsQ3CmV7YzMTQZEAQDREnQ9nUoWvOJydI/zt
SgUrHJEDRwZvFuE6w47Vqx4yQi/JydWyUpf+EvHQ9IWoUWOpNslTwLXnhB2vE0g6V0PvmkLz5BZB
sDPdIvMnRS2Oj+/PEbHiwivLDU8eMFdCPH9pIl4q5suRT6iTbQ7ytdczYFfKJzabDDXx6iFW+n6I
6P4gBcxEn7GOMSIov5FUJs0pZh/FMEo+AuBgoLnJHr40/Eg+ErXpY0/NcdRhaIdf5DifBVUfaV9c
I3JEJosy8PrXHS1gndzl7qPtNlmMSYaGxYClL41yel+uNVotffsZNkgbe0xDJV5pHmMqWkT85cmU
GlpRqvzK2e4oyHmDBN7HQV9sYJx/Bk07UTAlkXAv1ul2O6tuYjVh12ptABEGNWxvxZ8kXcU/AIvc
lMq/6QmHTszE31gb0cFO7u+mLkH+FOisQQoHCj6HcesIrC070Qweb4B7ZQHRIt2On0N3T0pSl9un
CE1ZRhncyfu+PVOMoRFlH4IuI8eKSFFkuJ8vWL67RQPE8wLupRtk/nRnQHWIqiKJ+wjg9y5EIY6Y
Q/A2DfVA7bTSbYdXJS0jXU9QFooHqnikezDGgpkFE0n4eeRnxMeckRh0o2I/7Zu2RiRsFbjozZSO
rJDKzevhUZ/kVi1+3euOmS9YLzRxF47SDLtTLRXiPsOsg8d0F/9nD0YQqsCcynTPrlgpWPYXhNMD
L5yC3gEgzsnQtaOuIg325Ei4GZ0WeSxv7ckFRZPm6OvHSc8wUEiWFhoOv2S1hJrsNNSveXK6VQGA
CooxxOY7Vw1GHqhTnso7mrm1XrtCXjT9JVNXs6mGoMnVZsd2QwmvRNsqa/ODf2Ac/QwCehPFRc0r
hBvtfiKpaM4LZMDIK0AdYv2P8mxpWccIPseTGdM44HAOuyAyadQOkEdbAQzYiwsi3QDb/miHSt4G
keLtARUKILjuXjMgWf4N7iovzqWbKaapoXYBkIzaQ+EmrtIQywbt+UXjPdPK0D3YK1Zyplr9jwus
GUsZj3S5ZhQFkSaP0qt1sJlH6UztMqXASfmkoKjCycJd+bIqY+ytrQQl5k8AsLUrsE/jw+WFoqB3
mWeKf3sd+Ly9KL8NQPYA3AcnfUX2FGB41b2lBnlqyZPFH+XdEmYSyhtV3QenO7AlPq+fbo08XcPe
89JAWt9mF0G8j3HBFvU2odih5iJYnMD8WSKH3iPJ6Ay8w2HUVqNKMzDNc1KzqfdT1Nx/BHfukHwJ
IBBGEQzbSr46qBf5f7VP+XJVDrTnAIy2tqp76j2IdDVmkW/5zjhFYoFSVujkqvnnwtwZKzw2kOq3
yvcENDUI/eO5G4CQgPLQaEOlDBbX6a/gKeKn7lD2upCG19lZe6n2N+wAJN4Udi6w91SCr9yKuHn9
gCKqNWE3lVjgQuJyqookUvj4R/DCSSIgE3dunf3Vkp4cbFt/OU6VoZrBMWU3s2C9gLzzGGQJb4PO
Lcc6khLfrYK4Qjcn5hZbw7TfvYU47mpl7Eb61n8iR6U6TD2mUK9LypPXFZb78GnJOFqjO3bCzWGt
ZfGlPbHTvY0AfIg88J7LuiTorOz3/Nmulvd+Zi+wTl5lte3aMaA1P3EnNswDRo+/Bubl7LAVdWRq
177+IhVcIwpa12ht0bXiOEo/LZb/yFopjw9I5GL32Knr59sN7XhP4LXmiEQJdlQITSIw4vobB/wo
dfVI8I4iw4H4Mn6fLhshx7ezmLArj+akq/oCPy7lepp6KobVvV1Vsr0mqxXpRo1/DIyuhsrV/GHH
DwjkGrTi/9lcCwYwgEdiaPSp/OxB4B5F94eWohUubc3vLyDdQ6i6fQoG3vbSeTSUAxFI240ds4oM
/0NjYWqIK1oTVqY1bqXgg+7f0QSRsqyGoDF1+bjPtYJGVkE74ufPOUDIvWw9XtVa7z1DsiwTTm0l
+4FJfaWvmntr4mP4VRjrr4NV9blKhd6BaoA0eG5vlvKC/s042JsxhAHyXDIJ0n9qUtDmCP7wroMA
FH3Gp7c9jMkgvrdKUUkD5OZn6xRYBHn0URpdy2YOoZ/SQKU6Ro5xqr0JbZIb+AVatUymN41EyCdh
7uN4HlL/UHVId3BwZSW5v2GvMDYkqMALHWkP+0NplZwgeoiZhGT73XQx3Y6bnmUuYfS6M5lPQhi8
BR4Ah8cNKdCGCrkWbz8G5gWENQdWAPJP/kJE8j2MtRg+f6s93WqYLy0G6xK16FH7DkAVpA8p/TjV
tn7BDmwzqM0XGV1eIQG7LCOvtcaAHBl/IScuweiO7Z+AFG8uH3iqoDYCtOSxxLNH7Lx2iWUkLa1D
zaTs5SnwZIioO4/iTAZxiF1gUeuaNW5oxH+k34MIAAT1nK9dINGktnWVT3L+C56BKrT6rRyHB54T
fHgB0x07tAI8HFhAh9GmH6L3ULwV+EheCfHejHD20jDqMnMHmRqIWx0JwPCV60F7rMhvvWrXn/mM
wBLQz5SfnYsBPIf0UwGtgkVkUiAwSl8G/ThkU+sexcMteFc6+z1JegEkMimLUpUAU2VKUnHK7j4j
j0GpaFSLtRaDkjmQZYWRJazx/vdhMn10yP26yC21zOigaz5K5gwO/rVTbajCnftbTKI9rkbqA9Ov
+cp3rDU3okDUd+rGrzDhcNzW2qnywO+fdhvDnogfZuRZGxbioAgqCRElHCoBqmJapDaNvpYRozUt
/rBIEiRF4SNtaz2Kr7Rcvl6+PRTEPeWC3+kmaAyMt79OLPgSDJJZb3TwtJJnG2Y10LQxIsNQCiyB
u0UcZi1fDwF9rsZPQG0rQYerE/B9F1ssuDXGMQgmjUwjvH98z7hvPtyGu6r7bR6wcTCywWaGodDL
aIo4Wr564sDE3dHNYURScDhA+GLVjQMDqaf+wo9j8RWP2tWgOOlKF9jEVG9wfVxZD4ODhhNEmvLt
anjv6nORgJnMHyum2QaiPqYPcKKPNngZ+w8HIIscHVmkug1dAcfXq9HI6THU9MfWkQmlBw8Pof49
Atit9oyUtlRdHeCUyS/RsrGdpvTtQuoyVqoPWrHWErr5dJZfvxrjinAwqx5o8kiZ1eds23QIJMHh
7PgckorQmhfazVVB4GdZ5Gob/TcRIFR26F5E1hPWoR8LI0lhC9s7/bj2DfsnWcbb4W9vBnZjCRW4
lJAH09T8sVrN/WnWvsAj6k5UYAtZj0QgmxQRdoJ42ETQ44f6H/i7wfG75LIW4920MLl2FKb6xZ92
NBUHArgTY/CMVmQkAswa6RofL5MZ/BJSwg1ZAnxAqWGrgzXP5VQi10JBbIkeVRhpjQxWUA/XmLrG
EoyCkN2O+puzmcjFcDC9L3hu7DolJ6tI/7yUVBBa7F3eYgMOctJPXux+U/NmlryPTjH2KteFtJJk
GOSd12yDRqAYae005beGd42IQ6069purgk1f4IJeHUVJe2lGo24tft4Qmef4f9hdtQq8Kqyis4VY
QneVcBRqB/EaU5n0/0CzQNb5Q30kuWyy5yMYqEVfHN51hzl2miBtyCfO94skEv83qkyE+rcDb3vR
oyCg4lg7q+6oZUrDe+8kbnk1xWD5PGtppVQPqlSRcrzDIKQy7cCTqKzLhZ93Iw4y0kUi4w1pslcC
Q7JjJJqqBXzzGOSt7MqclFtx+iqvA45HdHWp6R4nvv6Zj8+7Wi3RpWXfPlpjTpJ+nr4vThZfcpjs
uC9lFlQ/z4AElmyYZ0S3Aq8Q+X+u0OfbDpco/KRWDfy07HYzDYxDcco55JFDXb+310BgE+jp/XP0
1bbmBILg3DYdWsPCCsOtv+bx2iX6x/rWa53mOOFvwg00kFw93huOBJTXhXAeMvZQsbH0jJFBr0R/
1VSaqk3s3u/iQOAlEfSx0Fej3dKAjvtPxp64cNlJDfjmLdC/7JFJasGmX/JeEw6h2cphbdxC52lh
RlrdHfRV/afu6vP2540dUn8Q7PsFEweQdJNBriI4XvVdK+v9G8nZDffWCDLJbFk+06CfJkmYmxD2
cXpsULXjXNn/jLxl9wkJ/+CogR4v7s9orGHbaPJBOimrxdhI60KiJynkIjcVY/kN3aehFjfzS+93
zHYmFGFtxhPT6aPTc7ly36xqPwsaCO/ZrG1YOiZsZqJPzi7m5Zg5yNaYH7jY78iyjEvbsLQ4v/2Y
mx5nKsJ/IW14ecrWA2TroPdfNtcOi/2O4btEAUWfJ5dvFIZIENHcws2ICYbXDFH020lUZSj5k0r1
DJg9LtPZirCY+5selrvR5VnL3r9X7Z9A7uWZpvkZN9+wHrkUqHvYKFOn6VqBNMfjR5RcNog2PVV5
99Cue9Q6f3sZ9Tw1435ueC1lnYKjA41AsZfqXD9r4G4Q7rWXL2tywJF1HuITobDwhWJho2e3ftK6
yB8OY4DyYKfPGpGwZXIKRqdvYQEULmoN4lxLksM4l4Aw2a4UsALgIB0JeA86521Haf87c1cjB+c4
vdr1iis1WbS9txAdlz4yOb+N0gihipvwQNG1V/RDOeLktN631dzgxKHMFe4T/wkhGc4xdar30HKE
ses5QWABGesIU0lQjDz6tMm1HjOTfVIhtz9Qe6BTYBS3ZD54iy0JUZiwC3h3ukJRfW9D7AqGO22z
GIcTPeyElBL7BxyMZE9wNEZoiR/K/gzB/T2Z2kr44UJo2Oz70yX2CcNTbbr04ngNvlCdy+QV1QKE
YrhaqABSbeyl8KsLocP37vRkpAbMpSJY4iC5rlpiSNRlanHWYYsHOOVf5VLpAouNTlkiNrsF+6E7
ATSzY9c7ZzJTGcdXKIkoAWDTR6XkjEz5ErtwM+fSUEyo6GNDs0fsklmD48G2xekOktRHNcqgHfp+
OW0r+RFJwAEHAstoVKliKVOk1FQjOb4H8PNuFjG6r6nG8srUkjdtaHKkjZgz36AnVoNTtWjO7qg9
OadHalQ1NYZZLSyh3omTBRWwVR0ta9YdRcX3GFy29JuWubfkHudqYp+KFz2y74BOgGuKzszv/NBS
Ty2fQ9UyoJuYW83ErInn2krDgBfGJQIParUfqAN/EZ6eivXfXT6EFSMYIcZc2jH58H7nQWOZxYic
XymgyKI7kB9eQjanAZsvCjR42FykBOYzBmRBAXjAhOdsLrEQrLYm3vksBFeTpT90Rb/j/uH4SkfB
KLSjAB6JP+4yC1XumOlRK6IGGgsT6gqmDt3zAKZeE69aah4ziQBmWh/mGmp08FtmfKqlHOv+Y1TS
XXU7rLPMkSoVRSHDtE1GN72kOdVWFT6LpuuZAduffgr3ZldhoNnfVeC4o/0Zvy2W8l8IhshtNHLr
4G8bUehfYixYJXqSe7RYJcNwuPKvg4/rY3e6VWNAdJkAnrM7VYtGWK1Lyx1G7D7D1EjCpf6/YQIb
vml+oTR/GDh5uQnif0FgXuC5VY9soZ6zx3aeD7F2JWODZU8ZePEIsdp2cHemtYZPD9RLno/g+tbv
rK+9sIdu5ww8hl0H4iwNdJ48hELIIACRdeSCvMCJl81NUs0wvmV7bB0CUHOZZPYCASPOwF2stlIf
uXkS9RtXtq2Babl9Jjyv+qqbQk+8kGqiN055scYRID2w3iQoTjb6UgjkZEyzRujQgaDCv4px1NF6
McKfrK+CPCrbzBZbIcq4y83uEThSlu9dSd3bmktWSuxBWERJR+wbGuWHOtbBwp9jPsKPtUG3nHVv
buTHrVleUiDqo1Abh2l8OO1AVRhlpPyINDK6aLPvgVSiG8D8Ze7jo/EY4CIsOfHZs6uToMSmHNJu
0pTeDY3oZesaI8fPkSBbYFe+O3yLx02i95XBhJ1z4MBYUvwRjA/EJludWTdUCLCMhGoF8zVqYJZD
u6wG+ldZh0FvtFPhHuo0JeK62huuTkAuj0g0IMTP0bVd/Ypg6GjclUj8fpl+LvQh78sUcEGizCOJ
lDJmbaHWGNsyD5XzmM4WdN3+mAq79ywxAHO3bOty8W5MMlHx2BJDgyh0GgcRh6VMk1OEgIMBQ483
lyDsW4xBHh6RxPAf4hmUdjh4H8cnmu5GZtk4iQHTiCU07UqGGKbERamzw7Np7aDm9CiBXsQYbF0J
B28iwehrI/g/gm+2ZW1kKRQ6ZfhPiGsiVI6LEn6AmUCD749q+vANr0j23WAePUo6VEuBgxsGBBDW
XXdL+Nar+xXw48YhsR5Gz6ryVdyYexO6J3t+Nj6mlesCaAF8VyQbFdnUufPg+UW3FIOFbS7YzA7n
DRST5a88J+slD9qXMq0I587NqyRqZ370eYQRMyP2FSrWgZ1BillTZlac6/9BoT1P2nkYZgx3ZjD8
SjKj6iigNEiTPNE0zv8bsILpFu/f+wAU5rD+2JazY/MsquUcw9mxWQa47IHUSuj55xqFqou0bm1W
IZgzFBrdK6Yv51rhqRzix83EY3BX5SidSVYja65x6w1WFsiLNdUJaFSEMPn0c6VJwUxSiB/V2knJ
0YczxAQO4xYHt46op5GmYthGHDI7hlJgsYhfS1qfUTRJ62jWqYJ30lcCuIgpih162PDFuf9FdEI1
7sQ341pwST8LP00N2TntJ245LJdkWJar1J7ONo7jzpkm1b5nFdquVo3HORcRK2Q7J4oOeHVYxyx+
CshsG5mIeDFCk9ZcfpwaPuCT6iRc+6gSbChss+0mX30oM5SUWmtC771oRUzmodU04hOD/1WWc9+G
pFfCzQKVTcOm17H4L4Mgh5spa0d6ZZuTggyV+ReqMTFpuDzR0ZynpA7/+UoBieHriD7y4G1/nVoN
6OHWXnCVD6by6TEQCVd8vo6A9gVaJvR9dMetfrb7fbcNCR6BJhH9BeXp8yyBilqnktpVwk1AxFDj
bjWXUyOv3Ie0xdtXepKgm0U5Bjhu6eOvKrnQdT9TDb49/GJUeu1KYMAVKpjL8FaO/FGfy9MYYiP4
QRXxwSbK2qPINfX9XBVHvh7PMaPl3/OtK+GDZcC5+NruAjTBY9+tq9iq/dJ9sVKzgvrbCbdIn+aE
pDKQotoLkggwWT3WimTHSB9DEm6bOHxlgyBQt6Wcsja0G7im5DN66lDw5GKJepNWT7W+xKtBEKtI
gr7rFAPLGzJvWnhqIlrOsOdYjiIOViPuFfFedNAAFPjKjauS1YCTWbFvLNy3a5KvAVOTBQCKQGL9
Z+uxL8cf/Ij469Hyd9FlR9UdiJZT1wYC62L7JMSF8v57v/e9kuuYBpROGbVn3UNUtha57lvzUmXs
3oRsPj+OFK77Hq7BDqcv4hmCS/pQ9EBulRdR/MLG1RGmAsECPbRPXCAXqtjL9kkW2b+GlapREYHN
wRWQLUt3KRs0AWgW3zPUfqKBj2xhw+HNsoVH5rbbD0dHlOXxmCllrqxAroyIkBPa/hdiZRoKhroj
IYjGBVV5c7YpsPp0Sf3TuN/fCgSten+v5y14QiHkP47RlkMPGvz0mTcy5XSt4YZWdhJdW4ASNPTD
5vxZzz+mYZWfKWUJavsA9EzRuciv0Jc2HXeLF18frxOoR1UXzvqMemY4D/P+kN2Ve12zzBAMNECx
mno5hclpnBVtdfkvlJqajtbIa/o4eoMPyw5L1eOZ+XdbfdiAA80GDlUElaG/EGKHn+Inear1j8E7
CDsy/7L8qjMlodHtY3GdgoxET7yGPkGf0PiuwRNkmTcQGnup3ICxj8ze//sCKaZHLe3D2x/FCX9n
1fD74gOfB5Wj/yfLsKlIOyMWFqC1oOMaT3J0iDVQy15QrCsTkzcyGTvM8XIO/r2/0f4Gejn+dnqf
c4remhu/AO8BO6Ejs95qCBoin4PcGNguNlP/MYbDFzjKcgdnTwe6Wi46iNsLULtOcqabvP3wV7Jp
ztb2byP1/wwwB43v9Mr8qoOKnCFyK51yn8OfBrux5pQXOs7/SJERYEf3hwUu5EyN8xHgmzQTa/Kc
j4nmyzXCy1KYHiEYH/kn6DlUNRauWJ+KAKqDzZD975PAZ+u4pJEfUahRxWiYlfYx+kVG19W6zeXr
R/YCwqz2mUoS0JAqVL24U4Xg+ayVw0WxnmACCgWMmlJur/5Kw6KlvRlIuj9Fjd+vclw+e6JpX402
z75Zl15yZwfsEGZK+1xHJCWY6liZCL5zwWqDqI1SCw3WpceP8lcmd8RiHkT6JyCBO24MUyARsgot
OWqHM3oFHFDhMmuuVt3jgjBFkO3ruRJydl39mRl3gRvPhFdHHEiuBtH/8KXyMy2dmmNytNDMXsVA
Q1o8sR3qzVCyGqc2sylXpU3j6vlJU4cB5qA/06rWgqUb5V+olq+VJmruBpTaq4wHOKkJxEmTBYPr
HYg5pt71eXnLaWr45mEWD4UAELdewVhB7pP9r+rOmXWvAY0jizgnY/T7Gmpx1kTmJ+pV/aQ/Zc+B
8MkQNxRl+vVK7pZg2BtoagCoOSPI7RMBOxViHI6qGdGHnmac4TZJcZU3Bx2LtnfxXR7fkzTv/jTe
XPXj8kk21gV+FRU9tL+39vDu56VPAdz74qiTSNcFeNM588I7nBsi2OXK1dm+R+jYTpEBfkMxbqmg
F8Rh1EqIbeI6wkzJPZThfsLDjcsHr9XRZoMBHmVjVnenMQP0wxmvD/Ayc4dcE8a61chmozokBtxf
kaPMPvb1GEHysRHzqjAD8/Hxu4T66zIuzZ9xVA6nsUy2dwyulYj+mOsJ0Ih4E56Q9o02ej87bteb
1FHFnJ2gHSpyY/iBLrI5ZpwvVOAfMzEMRx5i/qdyRIuobWWMgScL21x8cZBamPOraNT5KBxyjIZo
sArO182jB7yYXsq6YbZdoqAPKy4WpMlqaBaLSAB/xfUly+1MXXvJ0jNrmVD11cMu5ayPR9//pWHE
TcA9bla5TSROgjJhz2chU1ii4EBFpCWyDTmb61xltWqlam/oLL5ilRP5fWWuUe4DLRB+CJz9TZJf
kM/IvawnzRGA3mtxmKBOamgSXWC/XZ/vXMRrom5xi+bEXPMFy47nVsg26TNGiIggha1chT9NdtN7
agRFn00cO0i0MqBotYP7M3x4qMBgX05OTrWAH0y8mNNPtceC0BLGMEoduKhG210hBUaDCieSgcK6
7fdOALyWvkBkgyPhq7/0e89J2eaL+ZPsa3GZGwswxK3jYpanX3SwQNT/S7fAT3KY7hOQgFGywW5J
iatf86cjNH593on8L4I8Whx8ckw01CPPROrQThkeQv5Dkzl2qlpDTrpo8/tL5PJ1LinR7DINZVX3
ylue06K7wO+V6+KMGPtAU1mWIMnMh1EoWEsAfsCj9ZHXIUA64uZESIGHgsgYusDFosldW1xAwRkG
MMxAv2jap/YM3I4CVMDWHAx75ITqGYjnyit8D3K26I085PxJw8khSOxyTQIi3dJ95wT+KtX/dArE
DT34jw5VeK+o/Q+trcz91A10szwynRHPOl/uZ2p1xnPY+DvsW5iRzJ8fq7r9GbR/v6P/gaNtzo7m
N5D0y/yK80jFqLi5OFFTula9avVU5AuYFTXKJwQpXJRPx5VXC+f36zSk6vm0GYs4/EK1918WofTy
sRYdtyPIWmFsJmIBZ/9h6SDhj0P5R7kbjFr+oXnB2iFkPO7KbYax2exryBq3NsK+OXG5v1lyP2Pp
K1XA58p+IFm3KAlzi6xhpslNLrlXi40zZnfEVWnEyISNVlxurngG2jL9D/JPGlsjY7JSXwsMkJ4g
7c28mX1ZEefIP8HpqO3SSLhQrzask0fY8zIlXVDhq54Q9xHF7/UAZHtCADt03B8r0vkeRwIOpsHg
zLNCM75slfO+3h+bVu/iGVzPn9UVhflGQKeaHyi4p6t0Acb4vBlqujHpOXC6ac/91UNRSDbeEpcK
lAKEen3p61mJVjLOPaO+CXTQrvrk9dn/tapPiDVwkRWzsvU+btm/ND3TWBJgAaBiyTZuiHygrmQG
/GaeKiSivr5O3P+VluNhicnAatyAebi///dymt5YgVqB1QyQNP3ax4y7+ht7Sakd0zTQUnvAuH+E
+gFI6EDdX6FdQ6fqPy+5dDpF8DKsxhTt2TR2rY+Zrt6jpbG5vFVF98OyWri3zNyXMpcdak0rq7/g
st4h/bdpI3Yd9kxZi5VtS1zKGovb9BDXU91ECiYGnpiSGTmRqBorEj+BETlE7qHhxBI2k1JHaz3Q
H7KELunFxZcDSwiQ8gtz6axoF2eeJrsV9wAebRRQtoeqrBUI/qkCvZ2GHFMMnhcbJ8Nbx/eHEKpH
vEGT/9FjCCq1gxH+cNp4lEkmYlJ9AXn6oijZWle4cA+Q1bidpteI6rujUsmr23qxQ7rBPwOmDA6v
9iDSt+a4OXugfZnvSk9RpPLoR6fRe5KsSLeSaYGEL2tBwP0/5OeFu+hmDJUg7Tpk6pxQ5IlJQoul
jgEzDgB0Jg/zvICpPzfxYP4Bc4fw4WGwVqW782HWBSlSAL/Xi2dmoXKrYIgfdepLhnJfBbq8eEp4
u0Ph9vakOxkVw1jUIFg/txPgAGTLZR9XEp86PMTxvrGt+2cYC0SrbyX84iE2NnZGpdRWKG7mYDf7
VeXcbOFoZjDnfyFXDYjiM1FUX+PIxcv1T/VzXKG62IkCii+/rKyRmlUu8o9OPPAhaIhede5sMlos
Xt1pS5/bQbDTlKF3ejs35TKGKfe/noK8oNyJR21vHU1gEcQJAxRKE9jIVWQZO9OwRpzGpVHICnSE
QT7KldIS4xYWYcfdgNigqgF0P8S5G4DstZ9MqPHMRCsdIXcS9Bq08GQbdPfgWkDj/UfiqJLBHXwx
IXwv3RVEB7jkYBNvwbWDeIeqvpuDF1hjXTCglOtZ3Y2Kc6U6V8ZBvglf9e1F4JBi1IK88T4DeQEq
Tk2/8lz3ZWb7i0vEXbCxZCEw9vx208W355PYnrDwBJ71KdOHDBCj9pJ1kiLM/OhBVA8VObah2bKS
yjgbsLTk1/0SxgMgUZ+Dg/8YbCeUzcAbPV8UvWqfCFHA8NlWQ9nHTGHm7Yvgo5uroFmXbsa6lEoi
yyvvqvWPGdvwMYR0Km9G/mRk5nzSw2sr3SHn7LTa4jY3aWXpsLKBOLdoDjvNiau2jYgwd1fCqU+w
G0WrFsm/3VWMIvorBYxhO42xXMKIpTq2eOeDPNi75B84On4bburnF8FBnrizR3+UgdhGwV+0H4x+
cpwU++9NOlTfheNrzVU0vE/4fAsfYCVcEyu1QtXNmT1V2wRp2OkuDS9OiO6AIvZ95M+EYWHH1pnV
jVWPsAjj85afTyblyO23UiSWHw6sXmhG1c62s1cwLUMVw67VUku7cVbROUSHiWVLUMvQPDQ/CWPK
ySYuuIt6Cd0kZCZjU7cYK9jGzAlAJG5xzOimmFwGajNsmgpxFILPMuqUolhLe8pSW1D7XLVHPKXv
P/u+/vfnlNZukZldZ7DQlqlbXBsZOLSP2NlzfhNt/3hYHzXfXqiMNlsFvEkGKE8eVrEcawwefJe+
wCK6QKwcnRxFRvEzOgGgxTQ20o/tQT6QMkUKI39mEum0U5n2VZMw/rizEkqTMDU5GUa4Ofxn7pnY
YSBCCgch+oWpoL4XsPaxMxBSJmrYZy3GINQ4pWC/8kTzOt8zm9wkXPksO8SwYblDcUJ7BGle24Q4
KA5+m43ET2g/4XAl9iMZEe03uTHUp85VM6wb4PVfWuXFI6cnWI7GJjIh9DQg6YRLjACWrpXDbcop
qd8EXHBunfXR0gVfHBKSrd9lu1uzp+lwgx/qoq53xSVNOrYLfLqpzosMrIdoRAW6hyUq0DKTeRxc
VQ0EqShDNmaN1Bbn+swc5OSzYLblC1UekQR2SLjmt6ZuxR7MFFUdkyeMgfDzMXWe5m1iLHbJG6SV
k3pyW6C5Zr4wUVgP4kOGuzovrY1ReCVsfOOo2RUtw/btTt9o3NQr69sonr0ZA9r41/u/Qbn0xLMm
97dygDMvlNiXl2Q31QmkudCfqnQz4hDwfKm58vi1q6RvBbKwVJQiwrShl/Pk0Yt4r6wke38ivbFM
LVY2BPe4H3kWqLYQ0p3huiXLrZyQS/5rKN3wTwn/7I/7Z696hpY6a7ymoLpZNRYd0l5Iu0jVhp/1
TdfwqnoZXBfa1atwk5dCUq45JKvEVJ4vY//NwW9GDK+BcOq1QNKR16tyaRXxvndgEY54D/QHmc/n
11Cw/PfJT7ppE6x0bOhXQFz2Uh/YmPGIusuZM8LKuTxZlXDcI6VARGCkq3XG+Jf/Wyt/f0oJH188
QmqHKWMqe/gX75ungEd8YdN1zt8h8k5SDQBT1jWJ0rFifH6eIFpmHlKZG9mN6rhTwNcHY2xt+DnM
IIuagxgmSbfP8KSZ1UP9w3TRQwzbkXs3ogYfz5pL1hlCNZ+kZzlA5znOR0axdWexwHDcb+mdAb+c
ZnIaV7r7IrcGmHfPhwk73eS3T9PnBwHwQTYFAtuJNwuvK3w9zvqsiqIKJeYKXQW6bVVUsf2FwqFc
TG+2ZOp1obmYeu0IwJHUOhmEsKO8Qy2H4V1QaJdgbCrzx3dZAMxT+IkCzyx4q3KUKpPdhXbwQXOA
cwgjMK8rPuCxhsLMeSdEt0o/lq6rHJecmHFN1X60WrlFOlB76yxLucLW1X1T7M37TTIgqML8mtPA
aWq06fUIwbIbGVlrC/2vMwvmUT7L89OFuqVr2HYfIyZ4LGDXyEPyTZl3PSIF17p0mFKckp0Y6DT7
1MOvx/OyrNQXtiPuA33qEbu8FdFKJfPKoT60L9zmBztjZ3TeICeIxdY9wa8j/VgdvcmV/sKMfDkn
l/h86DzDnItn0TUGIKzsTm0O30Nk24laIFlR0KrpIlDRYoYmYvORkgQtTdJR3xbvAlDBzbioD6r8
PjLJ613PGWTstHnUK3qJEh9lq7PzBHT8m00BbaY2gumK7vQJ2/wozrdXm7w6v+qu98zBArY4wFfk
14gZK5oDZkmsv6VPT5Rlm+M0RypsgTAyss0Yaij4G0OTVVHuToUncYES0X6k0o7AwsBvXUzb4zKG
SXcKqNNGcnZeNA3jpJiwp90EVqKmlV+HKczlRSOtuiT5uTvRkU73JlNuEheoYIiF/KIzTRqTXQM4
hdxOhLn0EfBnkePtaksDuroA0BAq3VjcDMCnAkxY4QSqocohV2ONABcmyDeuLDhlu096IkPNuIcK
0pfHLitLvDqUQTLtvJuPwWkpEe0zPQJ2J2PfEfSaRGjOaKKXNsF7Am834BBvyJeIWq+lXML10Nmf
kLx2KrSxHvPdEWALzTWC3t926umGLYs+UrJ98q9grmOsYrzHOiG+XKur09sV/2R4w4lo9VPnYJFB
9n3Ft2fBDeEHBip/mlsBlBMigcjbg+gZyJWQ2uZvgoRCS4J6tmMSST3ZMovz/Xkxf+N8taHwdzy3
ECPoVBfKUx0Jp9+cRpjHs+Qhg+cPoJp0VWsQlRJOQNVzkMKkt3lQmYflqozo7eC10jKytBeeDYTb
hhoKhq0rXWROdv9xH0w3xy8UCEtAMCkrReKzW0KYWYNbW/d0ydcCGn4Nic8l494/OM0Rt16Qzhmx
X2sKB2UBlP4r79hYKg2GBU37cj2xDQfQH6Yp5NoZcUqQs9B7J4tWYHJMwEx9ZA57yLvY3iZ3xqSx
DPpbL1ZopQV7Vcq82kU8ity5uJBpX5x0R7hM4JAZKuAItXN0y758rIlefoX9D7PwT4YyhV+meYM+
/v9Q1qaprlotf4Uhj2OcVXMdXK3zB05OkwzhoFyVrMn820kIQ+mbhTw0opizvjiRD8jmbQjq5mD1
jT0h3i4A8qr/qPcQH31M1qURL1o5t5NAEY0P183aNqhPQzK8hZRURkCKiDfZyf1d7vk1UrSUGBJp
Qzy94ttyTW8/D+/KRF28xtobSNnFenWPYiKwTgJBKTxe1/k1hq/+LQBUjmU5MD0RbOHBwxSMkCrj
u+Vteo4cEG7p9WrUgD7Vx3/33jAWtj+WfoALPwNLgxG4oBn+ZrfYYziHIR+lDC481CGeb2F9xgXN
xf3v3KrBW6gtxdcoT2icPXOkvmFBTSEIKzbfd2nGaquRXc2ph32PKtFrZlW5yf8YZdlyPr2EGZon
uXWg4nmeLSa1fWsJnEScJstucFpbcvCRejiISrRcGqYuagLBqr7NgUmY3UD9ajszFxIESboJV2Xm
asNvmVD5ub2xyqsicTCo+/Em+2QkxsU1uEfaeCyuWna8aiAwUXaTFLKAQs14dqYK7a1V1iiAXwmC
u1In1gArzvUlNZLH826SydMh88qkytoTec7Um8ZEpk7jeOzMC4yPjpF3u4aW7umaE9Wp6J8dPIU0
5ybliu4ryWbHKQexfQE5U6wAx5yzZMbSkDHtl9VUxXBZ6Ntc9KfDKkktw6eyUcFzBEGU6M12ReWV
k8fW9atiAASW7RdHylbMkFBXeJqheYrFJOZgnqjJSVwkkKbuHnv3FVoHSWCwtq5D9PVFKhIgVk3o
IS3HRtXeAM1DIxkiV0R34mECaMGNeE9+vixPYfAUiqS8sQE5IlwJ1ODIypmEt1bC1cmEue1nJ1y7
sIq98vlZ2njuyuWyhomjJ2Z9THYc5jXqUo7Tt91ecu+KGOhLIXBm8ejyLpy4PHGKAQxeJohPTErJ
9r3yWapCXa4yZwzlE+s9e4XvVSDdz0cAC7UUaprLC8gzHKcSCvgnhQLQqm0Oovvok23P+9KI6wyq
Kxwz8/NsrVh/RC8U2GhdlzZ9fuGzRnr9acZx70JStEg//fBMkpTG6tRiMMP3rhQ1fUeLppHRopO1
Tmf9YMHyzGbEAU9kcbnJtc7RhkFZRvibOrB6hexit3duTMGbYxzIPEi7/DqKxcrAhqao1DP27Ayq
qWmH2SS4Xrkkvr+uIJtwF0XIg2DGdUCp+V3kWBJhup4TFPnDTxzORXThAfJyI6v0BkvhKxR7hHfj
E5A2yFpptyhqVO91vLs5Fo3ZYAEF2M56LBpZ0R5gwzLCWPToNiP8mxYLNMohZZVh6V6hHd9qkrD6
iiHf+BtN/A287JdwPxD6I/ZYZqiMXgUUi8TIJ39q56PKTI13PWSxMJIn+wb8Ztu+sJRVU//mddFb
hA26TbifTwKeeClq/DXZ93wGydR3J+5C3bQKFjHdPicO9QKQ0yYxGAsY5wNQnB5FH/5q6G16vpF0
lMCHu95QMuQ/xKthkJX/wcXGki6Hv1tyW5Q1QeoO4Mrg4axDCBzfS97gfAa9ZMvGQLmflPomaBR/
6RkfdTJCRxpfYHLJBQXAtrUKp7W1uEsWgWX9DM56v4lRiDpT6knTVBn7GmTfsWz5H5VF12LfO1gS
wLj/fWjSTQKPIlaodk9oK/avaqhtWrI7KyZrB96N5e69cjHkaqbcN+KCuoKSl+prg2VJZnDuOf7E
Pi+k9lHFCkRI9WctEilkt03KNn7IKx1W8jkaSE4b0KYBeol9Ky5dFN1ehBoiz2biLs34d+dNUFTO
kou4ux9gPeedeGf3TKKoTnfu19SjmyTk4l/zuTIp3bcaBJGxK3i5gTaj44DLg37OYGmoZMC6529f
bPHoLOBmNj5E1NFALPn+Xb+wqELNL9tXaC37PsYX18DmwD40MKP+m+kEVgVvYsqAJNdm9mca30BP
fmUG5gyK3UKEVTZk2HS3ivZI8WosCRFgT8zYc1/PhypX9MB2pD3YF4ufy9RvvV1OrnX+disoDdgf
6xsWzm+1Ggc9TlvdgJP3EbBXt41nw8VCyV+slcIb5rOrv/T1kETjmDTrBskYi/dmiyhHR3UXbjW+
Ecseue9Y3OV5EEvXugpB0QJfk9AXamfYg4juQ4TZ5OUZk7p3ASGUyrryrhP3xCszN0IYAbnpwlvE
2va9arUvnHYd3pTld3cNbjrBdSc3HR7WS43WcBMjO66ACzdtQUyMzunwUg7zsrCPw8B4TNtEHV4D
ePa28yoWwnCVb5AHfIThCxiAi8ASmrl1atCqAglgN2LjpD2q9gRpUr5dXWlqBCrh8Td4gwfyqXar
D5XhN/Udk+1qatXuIQRRKWfPX1RlFIb5VGc9yUihYxscJeggcpr66EFC/uLASk4XanlKXaGrXrrl
BDvalxN4G542mvufiH8RC7MfhZP2QaSnMJkuuZLuFfc1RLmP4fSxAR8k+5Q+72I7qtUM3Fo35eHv
01BfhX48JhPaeNAM0Y7OsJLi01phvmCIfz9CYfmhyKMynpXaPkyPpU2SCWwsiqN/DALc5hcNtgmA
XyaZrtIBzBEQx5MXO5kBneaLs0eNKe7K7naXGzgdQHKT4IejnNLHzbYUGzxw6AIFhPW633xP9+r9
y765nW9OVx264OE4g+gYITpNdc0jSFIJqFvzOw9Hzing2q8bBQvpTEUWUwE9gT1rxvQNUf1Wzeya
5JnFIo3DYz5aQLR3gQjogxysYp5ovhSOvkXoLDWLOFwi/sBe9tYqBXlOuAJnma1xi+II2rPvUOG9
BwP9iV5W0yPIA6f2QCqNa/bI9BXSTxrMY6ESGJIrJt8cQtBizn2LGbies+BhsT5dxNh0gogVae/+
BWQ/EcKSUywl63bRDZuRohQAIPTTt7ApGFyPZmamAKukEv2nV5agzlBdk9F+7hHnzNqwrzN4fgkT
CPGS42MYr/RXN2gfj15QWsEUH/ebA/YGPNQob3PQI9H/2TByfyaMywGSawBn7tU3NdN/n0ZK6Wq7
tJsabH3YRPMfrC+HfmJusGoXJtJISz6Gj+S7wG7vryD/6Z4Vi4zgY9r+ogQT2PgaPHsomYrypAPe
Ds6o1fKXHZLZ+qZUzT9hV3reyXoqgc9ZZlHobnUxRED8unbT1OZqaZSBf7jVMmfRK36sAOCZdlXx
8OBZwzAKEhrGJ+YIyeNo7dJ3lPDWEV33c3mzNu3O+mjABsTZ3ahdfgzezf3Hz1uENem97Jqi34Yj
7B9ZQ7f39ablTxMk+xCLq7NXkAghViTw8pjyCuiYVVkECR/YheRf+aHXvyL8HR6XnhbTmnwn97Rs
/WxRk9wgRO0dSySsEDTYlMpI6rYoSkOad11pTH7HYYPqwwWLISIOIZTsnxnuZZFt3pqRABj8+znB
8AEZlc3C3M/mlx7bzzGN9Xc4dWYjXHbLats1ojibkL6u8059LJv8s+yE+JdOOcafH3k6OjQIAunq
eOMSUH620q7ogeOTKZ9dQVr+MBx26kFb3/E3JbYABul1sR+NdW+mnxz9wsojeSmE0oV4WCoQpmcV
eKKJW80HGKGWhsFmL6p212J3Z2pFSxLKaYEaDQEDIGXocm5oL3ebbuSU/nbQ4xEDNwX5WjhEVkfE
A4CJKqwkP0rR3nidege1rq+mICw6rBRRjRwd8P+hcpTyzMqz0rNOg7tNHtqnztTEoH8Tx/nBORPS
olPtm7E2Jw8xxjt2PlqJkY6EX6MJUTzOzslJa6Jwv2KysrTBf4BMwuXx1+XNrOUVi45q6Lnqk7kH
CWKu6VqmTHNErRMYP7g6/LqnQwsjS+5X4TIpv8pmp7XR2dMQApG0eWi+LAwFVj74XoGiHRE8RhKf
03N1hQvKFSePGdMMKix222uLJH3BouWQK5DYFynX22H+0CQS1/Dv1nj6dZorYrb0Ya9O6RaGq8Ef
GV4V7RNHCqDWyjwYGfl6+WBm6Afv91sIEx9NcWmzdTE0D9VKOtTtQg5GPwSGriwUZsxyx2dS9UJB
9sPCng9vUXXoqrQQ1BIqMlZH0XmLn0sNoVYNxeaM04RyxHs/K494YNAxRjBR9Pvk2wj0uIOZwg/M
LBVQKNh6gPA3iD0R/SukV+8mKP5txh970J7HVHs9OseTc6IcXVnc2M/Zi4nzfEb3r2inlEcm0mI2
S3lY/S+EuU3Jq5GxoWhohZO2hvhu526m+O9y8JAjgw28Ty8zU+10q3rXZDz6kTjq1c4cSUIUrnRH
J0IBesOyl9AMyS3fueAuJi/HJKkgx1nddcIx6dkjjT6AN9L2RFJGMMkWALyVLNczftGkBLpkABWe
/rWaUfL90T6XnRLEz4wvy5LMNcZOZ2s90HT7AQya+Qm7gajDV3LmNQ6jvQnK0YErzudxmeEZhxZ5
SX5bNGl5TAlMTFV3FiEzYguz5iCFLtIwUtEt86REhKGHSYQEBUWJY961q+wJorWyG+y8GqgeTVVT
+BdM/EDzgII95HshoqPePTDi6z4YUNJ408LrRHckOGPHyt5C+dKj6jxd1WblD6EpaijQ6hLpWCY0
/NDHDDezN43H4k8anb0cHp/wzKl5saEjIglnyL6KeiVHjL1gU23PVz1iRFRy4PqAC7oM9WxqkZIQ
lc5XBW+dktCWLmREG9FlJDhE7VQkWRJ2xcFASbksbd1VX7Hva9DosCfEN8XBmZP4ZbTe+37QUdWk
NSr3d/warL+lEViEEyCz+gzWLqJntyTurIeoYb2l0vUS4J9q5Cj0o5sGGuPE1l7clhkVrRAF+DG1
ln0IntCpqzhCt7lTb5uIC/mbjKCkDOzDADVsq3XfmTrIWRbMgEbKffLZvKuuvZfvnOpspG38D1ai
9Pe1gECm6gfBgHaRE011j6UWQipEATAVFqnwRnOko/Ox6FdVkyeA/i/iy1k3nS1cPXWIcJU76y9M
vpPqoqDG6zRdx+Ct1j2QtO8iCzkPWa7tdxgMu0YsC6KYIIGxX0OP5XtLm5wKYazFlTvKs3reVKiC
B6YVwt4pHr0yC/IYtEGBxVajGrLVVXyVNZaz0Zkgd4t4TGRaPd2nLDtmMCjCVaujoABc6WSRskFj
A81XZg1o4ziKoCt4HNRnjCooH2L+DkhU18ABKjWqi6y+JLmvOrwW8yoppVeZUJHrgbC8BLtfeyja
jv/uSXYUyA/EH/VyhP8CQrHhyR4fcM5rU8fwBYCHd3J4KvyC7Q7RectS0LRyk/a5w+JJI54F7xbH
535Iw1TWKkM2o9qq33ZyDVOwqSvJQDLSQsQGKYmcwYlsaxLnBmf3phnEtAofQ5ynLDi6W5y9CHmx
C5GEGlcQ2GDNGcwvXhEKAlCucFbhiBFPYQebdinRD95GVj9N8d44Zr+TAJSHGMdx/ORpdSEZ+36c
ZYliTs7fU27KJK6RTbwKzMk8cgnYwV8QiOWuuF5JXzCSpbJg5Xj1kTjnobTcSe8cj65LkAL4dqbR
1D40214iGeFJzo7A5qpFnHHd+r6YIISPLRBtQkjCuN5Jy6ih+E+LupAGOngoymIqH4W9FeNZliu+
dr8KA0Jl9di6q/zTl5yxM7xHFEwa1JWRrEU8+NapcGhT5KOOWJdk+obHiy5CiIDEuObTTvIeXspB
3kSp69yM/uFtjKgUPrw/vqTmEm+MMwrr9KQdd3RiqSzFEsuyIYs1zojuZsEho4FDFdGLqJdCI2Il
KwCuocE+YkUerz320k8iQi9BjoSFfzq+VcYDE3QdBOWXcsbgNJ34w9HZPfRmxa11IPAeeErrz2Cv
AiC0ASWsb6f0T/3RJbSdmU0OVMlL1GFCq0UVhoiEtA1tziRnxNSgWBO0ZuoAsEfSeCRgRCdUWqCh
Lu9qknbUR8c01qrsYDqDrG/zUehxTHzNHdYjMf9YMds/R1QsPU3RC4CsgSvmpQdjvWroOpADecm1
shVnJm2TDeCpEJsT5QwVRHdmBntJVQEB1FbTNAe1QIh2N9b3nFndjGMcdyo3RAtZU+HGLzHec1zT
umFWMUKvP/Q/CEG0Ib0Jg0fCE5uTv+j0h+tJWHgXCXdSYiG4Yqu5YdVH/VXOqeCgq3Y/82hL2KRs
os0XcIz7MO529OJWyWD/G/hMugg1TIDQzDFbuEiwAffLoDq00i/mHpR5okYOZ6O3MU0/RTfW8zSs
YHuxbpP9a5cXI85erW3T9Ip06lp94YRPMEjMIP2FLOMk/erVl3afO7et8RBaNdShk2aE7EMwaZfD
TaCPI1aNDnZXk4BYHMStjLp+iAXPdhEx3GktSlTKBi33DrMamyxUC266gBhrhKOLxtF1dau98S2n
OP1qQVq869zqCzHvg9y9gJDx0b1WDW5KKw0vbD/TPLXcsJQwaCM14IJ70OEqhxe+4S9vkTlE+m1x
Y8oSzbmAgIIIWLVju5zJ00fKkOkicE9iZmo9JGTKUnTfqC4YyxUxnnvoNRYUtwoqA/mjLCcOfiI3
/ykm27UpWNHTDhAY44bPRGU4wvaNTSiHDcp3G0S6Gmgrs9PY3Zqknqcc+eN5pHJKTxyJQgKm6kAW
xzGVJEfsZjc/AVRZNFWhT2GXWHU4MMkmgRuWtT2XjbDK5Gtf6Ne5x8Bfub11iwVgnxTe/CDnMqSs
1m5TcWxTq5+5/Ow7CEokIdYLYIoTANd+mTRvWL1AbZuIcwQMKaFevY9Ehp090Q2h974ndqEejfsW
3D6nY1oZZ6s+Fm9kMemmY8+cHn0JasiHMoRprZ4Dbwnmu2TC1TEkie8nusGRvznu4zHDHjf7ReL2
2sxu0Ek0Im2eeEi/gdYbhwGq/zdC0dMVG3QYp+0+AXv0VWcU1N5fjLuqwMXYgW3iWQ3rd9xdx1M4
llSYm8V997DBPw01ZtsJwgKWgOz3Oiv4TY5bdyCrIoICyr9+vh9ccKhFsm+FHh09sh6BqplNzcye
QmGmyeczaWrN7mQ2W5N3syz1nMjWEf9iyusx4mgg2C1iC7x1ml2AZzHZ2xa5fFWC4fuBxYJXbBh4
A1vuPEk7+xoT+iS4hX6UChWidtBG9vLuvI+tucuWRYy0lyI3/PHiTeztPamAsdJO0NY0QWrxuxm3
+pAp31uO5SMjpS9MoV6mnyg7Ihe5TYCphqeanakOD6iHRRRaDR4ltWeDi/Y050CLWUDRG58doUs3
e+jD0zbhZhRjE0QM3jwqezmlF/3jNLY4zoN3SoF/FJg4g2YHKBkpglDZ903VW1T54k1Wx0T5Mc5s
sGGEKJu08RO4w7hyB0wr5lSMa/9uhW3DmuIupBKfFjaoFpYLdFckCEh/yxJXTO/2jLknlReRTWxd
1zYIgE3WEOUxfyLQiWW3dC04bjURJXaQQ+L6mXSBWP/Tj+UDMywkQW7gJqYZZJoUycltyEWM+EPH
ZYdUI/yMZ5TSObEePJjieOyoUSfOK+3l9e+/k6zpOCKaN77z/xMWLLNB22pQnSz4gUiuax7TH7ux
/92WSFcP9xx5L2MzmHAW1pz7X+O61Vx1J1S6X6+f72UzLjPWILjjhHx8IBts01EOfIkjcXx0OldR
OEdObaP3foThT3GwjkInVg1hnLskPJeXWMRMCeCXhIc9dIqQPZpaYOR+/jnLNQrZYSD0kLGgrO6e
wn0ZiOEw8m0HgLZZ76kdiZjUu/3avpXE/HzJW90DQetgmWOnGi16BVfscDpqr036VXzasXDZ9Jzy
9d5VT7WAsnRtpi/gtyrSXE6CMtXeY6Y1N5DNFikuhFL3sNHCM9rM14XtK4l5zw0IB8EgB7EhA92m
JUkJoJoU3jsrApXjbgOAvBC6I1Ds9k0vPwo7rrLXCl4bArnk2DjbhtXVVTTS9zNz3wItJW0evfQN
h57//6Vtm13Lxo+ckuSJKi0Lyg71LoSnvHBdRFuKLv7PrDqENSrk1Dum8Aa/oCSWDVWUvFUudPd7
gxdQvmP4XDgZsUoadzAPnMOAoBqBDdJ2DIvZ5CeHZnYRAeop1TGvBx+B2areu3ejT1pYwgTvtHxY
L6cd1T5njOOEzxFqT4DLHx+OEhoYniGiuiEkBXsP4Pmp6Yp+NtnVN+LV0w4HltwXJo88SsZt8zjP
iXhai41ss1jC7lSD/A6wM7eg2SKy26We85EK/bc5wjxqjcix6igfjShp5YoLbouvMvUfYL4coQBI
ORYbCtkrudOmZm641mcx2+Mayp5LIlXOMEEg6J8Elr06AjWcZSNolWMc6ALkIQypuY/PCu0GmdH4
x67oQGlMh2dFz7wY3/E6xpOMvQGC0lzBwYtdwpvUwL8ciS+sA52EFAvhfY9wBxj1Xwm6TTAcpQXk
nZtKeFKphyiGlsrKJ0t05KivM29BjxF25ZoSw/PeQBeDhqvUsU0exsnNwTPohGICSorfp7HFS32H
JEXEyEL2+mklNDY8CU9ovEhYAWI1woHfImtIvPbsENSyuYEmTRh1Zglz6ULllFYq+3sCoY5rUgFd
k/eqO4rBMJldg5SUhd/KYKudJ1crl1/PGlFmw/U1gxQPtatlowrAiWGSNqr2cCKpLNcgHM+ED3QV
cXTK7JE8+Hf89sf3LJbTpKXWIbWBDk8Xecd+qJ0UX4ljcX1EGtgHTjNA9UeWiLlliA32oEF8jN7H
O6lGLqCqZUOOSwL8WyKhvbbbh2epCZiQc3CDDWXVjPgg6hI+DbQv3DzrCkyKyIstwgzcjXyIzNWF
chdLcG1gg4DcxDzxzcgx4Hoddo0LM0PrWEdAP6uSrR1VM5Y39soXbE3J+3h0R5qrJSWsyP8i15+B
a09OJ9hGHQ+CRmpEHq6XRIjnmeHlGz3zTNc0+ebDu/haOMWC/Fm9YzPCmIrV5kUxWU7i8UEuLfsE
3M+dqSlK1CkmQTGxox6W6ym9TNmiy8W265LZuExBD+dmOHz7h4jzha/uiudmvP4+jInDlCByAK15
0RInbLprU9F5l0dM5/jNLBjHUtHZSIjPbOrrwAC62cr0tC5Q2eZaQC8Wh5HsEaKZklMwlv52pS4b
DhU/MCKU1v6V6Nf7tRCSz4kARR+TVIK9nfByRSQhFqayHkyK9ssOZChHalVII/3Qa6JzCLe7kkTu
D02gA4bZnnhCL3sRm4zPm/g2pNdnYRBFqY4+cuco43PPZCR9BN1/tSegpYWTPTZisNAho5pPTLzq
rhrxSY+C0yt/K3mgU9EMR0scTIts8Bc1+W66DNn1aa5lIviUEm8TgLMDGwiq7/OkuYfPJIcAIIEs
RQNoqnkkBDRXEydojV0FwMlSYbxIRIcxSiIuzKHnN35miymF2Os8pgNIyKtuwwOhvj3xeD+Ev5iy
DeypcEt4T6cbiWBc3B8C2a34fWjMzcAjgbNHeCdk9BtGHSiNpvW0x/x+ldqHsqHuFOBeZw6iMXdf
765RZjK5q9YLFXP7GJ60K3eMD3k+UpzEOfTAjQq+htSWzOUGjnag8o1GSAzfLFfLlD1wyvt0q4Rc
db8bw42GaIvgB++EbDh543893fcKmhjm5+YzKNmgVTKYGnMskihHPIZvlRlfRXi4xysjsJXaSivV
o65W2dZctLg8ac72Tan2NcE2IzAfEwtmhhGhWWJBQAOlbhw3HU0kxhWFpwVnyeKzJpxYNfF+ojh2
3beqSWqgx7Jfj01nChW60ZLPmhX9xLvySKHnep3hY++ERsHT1nx/weouLsemgCd3VZZvMYJ7pmKa
cOqBwKL28+7hPvakn09XKtUdxK36lpSaQtlhkmipriT37o/2bbl/Wh3qLe3nV0xMuD0hXVYg6qt4
VuH1R31dKmykjTT+h+jrH93wROV80g30tXlO+WM+IUsih3AvwNa/MNZjrGG6/6W2GEwoIgeLhnHD
qBUb/85lIZNxaeiKDjL4sKg32NWeiEyY/ZEdVeLvgrI9FNyl0dUHVTTzu8czxzv88ME3f9AovAmt
JOtOEVzwTe3D0hywA9666EjZfstWtmPpYWhrwiw9jXph03q6sFU1WXQlb45rlaMNdK5mXTQnyOEu
4BUNcp4at3h8IEDFTPp0d+qvKCvw4JDELHAatwM0vpPCT9x4US/Dig83boFfB9Vn/MGBoSp66d/m
Zp0lQuXvLcxpEPipEI89SiNEj9bk0cOJXcKp2fEv4HjfaOQ9DwufE9OQSyq5UkxsmHjCikxPC7NR
bVVIsmGgOCqCznbjqmxWyh1U9/eA9vZEXKJ4U1F+ZBfDMkBoafgXVMwny5S/qe3JvgFRz/ivrNtA
4+sshARuTRU+45Vew9n/AOWJQA+rDjyw+j30fvzZDROiRxW7gOe5ZUiqm0FMBzUdC6qwZia6QIwn
eKmzW7KTBOc31zuQDdG4SvYqYuKc5NjLUrjcR5EdVE8gMEHEQ9cy1AK6kSPu4TfvEkd8t5WbBElO
xqQGKedj7w+yVvhha6GsRgEqTX2gZ76Z5LY5IFXzxuck0SViWWD2ZMJip6MGCXkuUY5YRZ58ICLE
3O9AyPvEoeCb9pcs9VbhI/ikpmwDqQlvhINVEY2vCkEux26xXMbLv4diNzbdrcIXb/gUD7U6qDS6
tyl+6muTTLRZUEFfz2ooM3gRy3aMMOFD9zx/6ihr54Y3K6F8V3ZQC6TApZK08nN7BPFIQQ1DDCpE
kWmfqlKa4Pktv8I35K/eiLdf14Q3/umeciM7ycvwQinfvx7l1zu2PT2GnyYQak+FcbVCBf4a2QR2
N9s+mJidt3RYWdI6uMdrseWLmLWsA9zej8JBFNL0Gef38Jfwh8ZsUUH5kIiJmWPnZqE3101KZUjp
+Tdr1/H2MEavIyKQZKMfZfgFGJsHlNVh1OZORrb+BfE0spL4I5F/lZD3kskVR/UDBRxjf76HCSUP
1uscmWxxQPyF/GtjbEQnwEXIHAaLV9loyK9s72Q/bl5g2o20AN8P2yb0l4cxs0MBEZu8gotSXaRB
D8lOR98ynq/m5XXU28hFQosuGHmdEkvbMu7CsXdQW74tNKQVqoOzGZX6X1J1/guajFFNlDW+3Iiw
PWMoWNKhlVFacWI9o00nBcvI/i3+Ss4nsXt/PrTEKI1KI6coFBDnEArmMhBoyXyxXeMTFDHVoS1Z
nZcPablE2cJjXgsiN9LSmOCCAJy3TUrpCu5vM10tQCWZ54UnmuF6e0DzaLL9h6HU6q0D3a79Qo3p
QrzRtTgpAGSFTteqPcOjzZu5QkMTyM4jHcrWlK28pOCeKEXQgb0LRKVJFQEYe2W89drSsAePEkV9
fjoJYrChG3QKZUYIhmuJzRghxtmx9apu/hL9rL+/SB8AliHLKewKTq29CrWzZI8seObN9q00VQ/L
Xo6mD0ujlvwlpLncEJsaZgYn7fvGBDZnfQQabHdf7AmGCdfTALQPMaCnCzEKHpE5fysPiDSyPGc/
CwvqKvG2r6YYtkfZbVC6Er4iyTvgMoyQnBv2B/8PrWIa839yRb8O13qCZ93hZsDrn/dsZWKafShI
JaiX73c/U5FyUaXlplSiO6MaXdbTn0euA+rX9PYjVAnc9AnlrZtsNk1swIjFRRoe9FuwKOK+C4YG
Mt0r5uk5o+l/AyLcNnaN3HKDyOVTJS2mtlsDGo9fj5XWDvxhKamn9OtehE7sCLqq7pSwA0bMlXHX
AG5PJfsVa3H6L9sF5Kj2R4qPegIcuWBlB0th6q00Cp8T4SDe3//KhzPH9C25PjPj6Ct29HPtSJ0f
gzwO4bWe+a4yg++MGcpr8CR2UJ9d+H7VlSiWzoNO1q6EorOdZUUAfGuvVTdG+jGgQtqpmMl23zay
rX5Lz83PuSfSJWBm8FxvdH6QcP6VoqsmMdyfDWcE33Dr63TKR5FeaYt1oTUCX+Kxhcpr+Dg33+YZ
UCQd5rolGc7WK8KoxAN9HDXb3m+PM5izViGLGskBTHRaerC/r9+BMtzG4mn2+3A+e+7wtdwMS+2S
62xve7OEJejfsWlCKsXRZfFj6MIWiWHhIEFTkiwZxNfxZ1OgES1oPP4E1I5pAyvk9kWXZfvKpQ9W
1zw+d0sl+48ZP0TmGMBMGSj8Wc4A1utFvsF+NNeR5YXGE5SewwLja8narQ++Kiz7NlU02kCkTWEZ
HfNKbDM8vRRbOFhlT8NiNH+yriYT0PyRWgdFzeenTKfeEvEbsr/1zO41Q6MfLivtaXcI4sOct6Pi
wnMel6koeCF7bi2/R6f9u0NJkX/AFYTLGJaHdftjuhFqWFDhW6U1xLguS2Wb1rz0U4P6/X9AIP1w
DHhmVKXs+skQiTvASPwDbODAENYQF/D1o5n+Kom5aWyoHK/EmhugZJtinFxcPHOKK50w4fuk/uL6
3JIpDHR5A7krr2MUMUseMSXhSeBLHjBFuO3UD8c87ofIZ4a2sifVoW852ZgJmzfrk9FLJpg1oPOs
XWzgB5T+3uCbDEPmxUPuqa+iN6d2D+iUxgpKwIDsbbbrsBAoaZoOcuQgH+ow7GtKkNbOYCqojpLO
UimbUTM7WpgnNIKBQuYluZRd0AW3l93D9gyGYbxw+jzlWtLlJ3oa9StBmtSwMbw48C6bBky7t+Ev
Avg5Y0in2IPPiJZlg7SeAMV5ZN0+YJFE2gxQTnSyEq34Uz6lB+wfQ26JUrhO1YJVkSJkdg1oErVZ
CYO/VB/j/Ffu/ANDmHt9zN6anISFbRqqt6g4dp3yJSCRVJf/b7fhUQZTIqh32FBK6gz+VN7HPadt
R1HmrUOsLHcxiZjmGFoZUF1LLuQgO8BhQrdsl3WIGfKXo5lD0TcHXWjkkHACqX+cPsdrgffdYBUA
ZtPLYQc7umDty0abTq1QlZvyp+ONQCopqUpcp8QK1ezvCwa78DS18W9ByI44q6nNPCJ65XC1WVxI
glg3UVoGh5a0r8n0Lv6beKL75EQXiE2UFibhnFmAS8FpfgxRW0Gat/ubvhTzYOFRTf3Lu0R+z39N
Fov0X82En37kpGc/bar6ujl5bdtZ5LBxXyJ9P2FPO+YsaWQzEvxd399MzubezQ+hDizUJCJeOlQu
OvxCEJyTLD90UYFakt7dJEbFByTw6z0/2AXX/tPbX9iT09oDKNoLAGaH2a6v+qZnPR3oG1aq+KY/
KdtQwqcBVRqUKHxyNEnUsVtUX91QupW3RjegwsUbRkM2JqnzWDa0gjLxC2xKLbHVuGWIh/Dmwzsv
ZBSDEKzvClmX1Z5MQhennscwS4eiKtn61Q6pb/9GqVj4fU0M+pN7+yDgB16LKyB4lLenZ5OgYy6v
I6boF9++xkn2IivejI2eYezTDsHbIGDrczRjzjP0iw9xlfkPOTvBWAwtuMAK4RcSgzcQ+t1vOH6r
pQwRvL60iY+K4h0At6rrWbfgt8h52SsAzhMC6JKIODp9Mr9y6Xr1YqKI/5DUlSuVuhueDIscVA1m
uFdM2ER6kIpVNwC9K8ukA6DT3m1PT2MrWUYIkmVuvgpsk5xQVQ9oa3nADNhASq1R1LX4cyh3hAiG
9/7HHdgZ4bIcvCEjfOrDNHIxGTjNp/1+LY3fNK1xcLk9emdjN7LqBlkwFUPw53Nv1yPe2EQaRaxp
VhS2uAwocZmHNFbueAGeuoyVtVPVuei8WBt7pCmC5foaAZg0COhRA09jn+hU+j1irqLICk7oATBd
MufuhoeVMzPTO9kp7y0FwbHkJiMSUDWQfZO7KXHP2NE1109YB5aDloo+c0wrwS9gWg4sAKRpxqQu
qEP/diDMjyBAinbfeX8lWZU+mCjCk8F1SMSAKu8sU/9pPzkELdaIMRPjrKXKbAJM0B6DTv0ajADd
fJdrsfrZScwZ+RjC3dRjCkFRABkPX2Er6xHtZHOMv/e4XuWLVmwpzX47vJDh8OCWWuF8Lvn+nqyV
w8vcP+DiBa5SyiIYbj3pAYLvMESIA3NxXc42HGonOKyFLR/ILVtaZi3TwnLcSt1yFSvMz453hXsM
eGTGdWL2CtNC1Krwik0tXKjgQUidoOPfndnjqmYSFk8GnJOpFAO36Bei4i4+hL9pbc0tvVT38YWN
GUqAynL4e2gSWt8LupbUetFTrXqj/15EXmm/x9HU4AfrvsCWL7Ch3BhkB84ZB0ccyOrwMt07yODX
LPOEns+GjHwBqZAl9ksZUodIi68PGph7ZJs+SIUFBocFF7zZHRj8ogy5sbieEY4Q+9v0BaeSe150
8AYrbDvo5btwLIdd4ZbXTvvkfoXIJaQuZYA5xcfl1JUkRK1CD44qwo69L3pmay+qmS46JTZm9PFB
d0iyROzXjydQDrkSBZmmXLZmYb2BAIXCl//iayOYGjfuXAyrdlvS1ABXuuEAHo5WHiocd7pKmgn+
0qplyONInVvN2ItHBHFcPoeSp89DgHkBg7Roa1Q6bNTRgQJ+mf1q95o8rtFlM/2NKD1e9iwA3SR6
1FMGr2JejXP2LoRvcMuYyLDcnGlOnbjlaa022p/VbcCt/F8mEgfcnkwPIKRamQvck7yH8JRSn4+E
27sqGKFM5BhcmvOblXqg5FphIs0nOVQxzjnQ7iriaFCOnTBg2HUurL3OawiiHx6VoN2o2xWLf1eP
pXRx6iz4Z8yfHN2dJOk4J3LAmdkDZeEPluCsFGbsJhevKcetzu4sE0wOb97M9/KZgVwcTqG0lNny
RB9PFASQUwd9sdC6VQp+4g1NdItCVeI8CceRCFg4A/JY6hUh1L1Y+CQxGqc8gzVcbYR6grLEN6Wh
5YlVpjZ3+3fr3pYOWR1jNriUuFA6VSJ1vmfRotRQ9FVMoTlTovPG46rsgzIDepTr+qto2YW8+LJG
47UKwUvvocMNhNhMk07rPT6l9WPp8+5yWPinFyd1y1ydyF3P2JcTeso4c1J9zal7h+piG3gzdgfT
RS9zAYJsjjhJx6qZjIeTrDYq8iXEsT+6NihQmrSmWi0XnadpcBkafZMvlegrermqeD0FK7HpAPq7
9ySM6IWZfBKF/eqmFUUzl/xw0BoY+1/a4DxrPH1nEqQVTSIjoj0cfn8HZeaG8kOqzsfddQhIC0ok
94sPyGJSdaHi6GZUWkneYtKaDcoVwN/8QCsOxR4R46Pc+uQjECvzZcGNB+aJaQEJm7Tio5491aMc
15B9APCNW+784YbtQfjw/OjEbXNcZinNrn9CTANBB+ur8ZxGg48Ph7mbJKK5i9/sZS1PDTz1Kws8
+Y7XoEWhQFAQtM2M7bDXxUFFsLr2SqDVXHbcRgt//p9fm5Af3jq1o1UcMWyQNmZv1iO6WHgUmQJz
f1RU7KyEUxbdiqveg+7H1yLPUaQ9PKANYwJs5cD5hxCLBBPAnXLoipMKm6vEvsmNyMHk1GG8Rslw
CXcrd0zoeVcYwUaBp42kavcDWe0oTpMXEyOeNXymcxvufodYojscEnkhl3ClK1acjoiwx70qRhpB
HjHoYiM2A5RCpRB98+2p/dmO4J0W1MKF2ZgLkbXNF0f/7FOv0Zw9wqmsSThGq2IJ4belhWCgscSz
FQM0Txp5wCzzi238I7EhkEofu936VoWHkoBQhayF1VvD5ods1SDWDmRqOx3mhg4yiDrR3ZziFH/7
b6WRBuPjzNr8rB1IAtNN9V+6j8+NjhivbCsuIZaPePHwgVGT83yQQlEbNl9stZeZHTU2tx/6rFh2
UR/mqVUHtkQuop2lRMajzEdt8wQPGlCDR4N4oaVFd4CUbQ+SGfpsSnKAzbdGm0GahocY7JGSgQjr
KSRVMpgRvmkqK1w/yW5dPXUWxj8ccGJ7PeEl7SHaNIDtBFNMk40tjHtILYgvHFgomPNMVjlpih/b
edwiV88LL4RLxWS3G0Z9PuyAGjepsw5+9v208iyYvJedvx5bb2lsBbvPCjdzOYjo4HZPNqjUjspN
ZSyynPflGHSZS4qb1LqtXeFpvbkhz+mu08Htb2YSw8VPZLavRBT6SOnVss1/8+MvfJC1Mh6o6mZ0
GUAkrwsF4mFK7K6yEcjPp/7qSvkxl4gNx2lZDjQDp7uaSZk3N6UMfH5qfVo9VV/X0x0VjUbLBgG4
J9cpsRBUgX4HRn1kyEcIVcZORSciNhyDO6NAdg/E/+H2BZk65Dkfgjk9aEkHhNu1X8MheTwaxau2
6X2/nUES2/0pS+SUJYt4TZGv1ARLlNbJmwgLp3oCt/C446dKMWk1X8SMCQ2RZB1QlqAQ910K4z6Y
uo8Xunswxp4Ji/9ab0N/bFG8PwVBKcI3gJkQwJVn0VZkj1rPgo9myV8rTwN/YOsV041tyqkMv8uK
MR3NS2GrllU3gffk3CPviZ+6rTHEgF9iX5zFaBS2y34nM4c/9IYC2TrsGsbktcAbDI4OB/5szgnl
y1mrWaniX1/fKFjcoL6pW+qBcIeYBf5CEV9fxDwRZtTVXf7Feghs4ByKMLfZ5+rW5qB096Ed2lhB
fjBXJI3ylHFyhzZoV/Uwkxq/An4our18hbkdGJTX/kXshSwe8hF5KIbFvH0QZ0PXE5OyPjA3SzKG
mdWu4dJy8sXxjN9FVKJCKoNu9GB4W36ghhVstoK6zHw3627XjoE09X7RwWubwgyB0owXJT5kcjv1
nEkClnzmg427wQYwDnUrs/num9LxgQD7RyAdCsUiFNQ0wVbuayMq3Er4xifsVL01XLQXllz6Wcqe
qL6fuRy//XHs4hGiX1/JGrh9jrR1TLEQk9iilvam3Kz8eSgaywJLqFf47yHRj3vGGHwF2ir+fj7Q
MWesnJ784+haOI2NFsycSsWEsMi5QPtQMf4555Th9vcaUZ+vqAVTuTV89ZtmBQ5j7BGWLVoKk5pG
Y5DnQyfpvahcGEIr44pMy3AOhf5joTWlwik3YKZHDZZCoHCgGtKpOs7O7Zp1G/OonGkhj8Sbm2GZ
iDiNw//Mr4gsTrEaTp3IqrYxV2bPywFdRnPceozEW+xVt2qP9MttpCq3P9TObrBrZ7Xybs9e3LxN
OLnJkGEbttNLp2JbqFKowCn880G6dwWWNOYyj675aZhCL9JihJun6+pc0t4O5Wi3tHDdGy5P+aFk
uwm5hrIaPwXItFb4QDhhJ7Iuco6v74FG86PlFu5ExMGAn1BBkojvc5kcpMjZ7v0inIt54bBFXTjn
ch3CPp8ObcTTc7WZj3LrYyBmpB3hFVRkqsQld87CjCm1p10NbG4kU/eXgV8YlwbkckYAZu1QZGHb
aJLYYZGzmrYzkR/3KbqS+pL3wHNizSnBnBwLWesJiyZm11NW+eXilyAJKR4tSFpXheAoIhmrQTbx
1sEIlygsbEA8Zx2YYNMegZcE3pVBpDgutQqM6Z9fgspQPwzZSiGbIxYpLUwq50tLYc1qHEts1Rki
eltd1fLtFZyuwqWEVZVYTLo2lr+ZWmIRKKVtXIPvQNLCzGy9pdgL2YSozG/IyxXK815QT4CkLUoN
Fhx5CXElLJ3mCaZjHlnpeIe33TeMZQfquJu/hzLNffbXtcveLWm+kS23rMP58vJE7csJDiR3rBj+
9X/5FC1eNVCIKBMt+VVaZgb+u2FRZjINOUD58HUj4I7LWwEl7yfT6x3zhNbueLrJG4srXH/CQEzX
zTJ0FMX4gTcB+TYOSE57Z/h7onIZd0ue0C6QjNohtpD86r5xTYdqKIQtmM1NJi4YuJHNJfvf4Rxm
9A9X0/Yl5itqRFVcghmn2t0gzbiVf3qmuuqgTUOSyMRXU70c1eLurHKAzhtXzRM08TnuqGsLQVKM
uEVHtRcNoJWMjOJpJk7G7Qmlpc3nDVrNj+RiR4DEfgW+u3lYdV7U65Txo4oo+VV4XdjCfUBImAxk
XJLNJNLR0xaleyBcttbFJbCGEqBbD/GPI+P7uI+PU8tSZuz+fw57s5gtVtqyYb9u5E/FDGzw027+
tTFJoV5n+KfxSK4mZGWRtn4KwCPbXMGGTm3hz6jXQH7hiPUYSJshM7orRkmZFajwsuS7kLf9z52w
0b90BhDjJdP8X4FykUlq1b9xHXZdMR6qtwg9bR79Sk6bNaDM2GlDSGW3AqQR+jhI7McC6N7ZJrh1
LshsOZOis3oXLK13cgE6+RLu9Efa7okVNQq8vOzp8arDhUjHWOhnS1d47lRNLzBrgX7uNgEKUvxg
QnT5xqnesvkHOtAYYidMqc1VUUypmhWwAH7M5Ifie6MmSpV3sqKkFCimY0opSw3RcGwKl0/U2wcJ
UTWxrSc64opSpwFyXD606WSLpDCibHeYuRERXr9YGfvC0zecnRgF3aNdKVU/csUtSAxgjXg6k43x
o+g1d7q90wqwjnoKFCV2kuwzYkFckTu9P2nkUcSwOrOcSmZTQ+Tr7qV4ArhOGr0yQ+3Ch4sooXUa
yqi4Js6McHztVpIAAXfZDdTYYGnmMxCKRTI2wBZepygQ3H7c9DBr9hSNJoSPc2sndhS/zwVoFNrW
r5HlsrijpArJSeBB5wP3WYsI3eNMfmdcwVkxGgftSJNUzBI8VCPdd+btsv8sOCLDgrMAzeWgbgZD
uFCsYO8s/OqAK9WkKLwfrmqKtSFUf86FDvNXjloCgzB723+xlKLUDv5zZlqjfBweB77c82GiwQOv
vY69l3CEfDmJ2yCNmw2jfXVRUwWPDziI8mlsU1KAhF408NVLTziqx5hSVHj9neiOfHkMmC4Hugko
No4ovoBWEV4s/nBIm8rQu3dcOmLatVegKJt2sksQEa27gz9o0dfkAHUtiRinXwqT9n+LjWwtYSlE
tgjTpNYNOLtIeAn6GuiN8sEdRceonwgCGhhyP9i3N2jfjBiv41HSBGHldSMarceCH4SqTcbOvH0O
si44c/ukQ/5rxqjfGp/OqVg6f79++4wJMs0WrCpB69EiZyNLYumnkkJXb7AwEr850TcAufrlE4sv
vo60JnuLwFNqvKpZihem9LUPPVUMJINOvOIiSgg3eWwD2f/6zCSPZyhJhFHWLIJ9K7mjY7Lpr9Pl
9wNsNVJa3T7wKMA0ptDVWhU+0jOayJqMWdHD5Nx5ZVOE6DYbqd2yKBKay+8H6VaZpJaocUzrY8Wc
lcYdbsNGmFG7ERzAnidZkJHSaNpOxH1PmHh8wQ4jXOkNu42yWyMOpR3I+r2J3o5rcAxNBJucFDk+
hHlbSWwg0Vxo2wlZusBHD1vbJ6DeH75xh2hjBjUxdv46DUoXfOrVxFrhJ765e2NjBGkyp6EqR+si
F5jcXfCwRXiaF4ysumLQhrVu8MK7KbXBIFbubOBx4aWgdz6M+GbYpSUfJzk1BWsoh74iOjG/eGoS
MBGVSTK5TJWia1WXzZdvUhE97VYzMa8oEoRF0a8iF9WBV67BfNb1q84kk9h2pp8laXrgvGvxAiR9
x0wChgtYVttyYJwqrTnuM0xXp+eAxVFgB6naJCqw+CTCozc/bx1xlmiKUd2NLMmk1CKcsWUEgN1M
Gd6z8qAxEjY01KOovEllC4oi1n3kWB0lElMxDHMNcKe8XEp3Ca4JhawhS4aHDNhdm3eE7oIHBnUT
+j8I/TqR2H1DfuVwZcGGSt2huBatR/enScvFQAP3j95Nmw8KQE+RR9mD/4Da+LCmMudLjsg/MsF5
zeWvfT6UNjellE8mw0eWJ8kO0eslPtQ0nQQngaLFabxzrySqE2wU1XlhL6C0/4PuZNSbnCv4pauf
tCnTfkv+u5L0pGuI2UOp7+PlfCw1NDu6VKSdpZKEUfKWEq3M7Xj2pINiqRyF0iie0aj2/NpT5Txu
Ll6Qvz10Kgs669La0d74tj6cFITP/lp+L/Yme8QjRlw1lS2LROaYpeEA60reqvDxTwpHJ1HPgZ7s
Ccxz3fMhUPM6heVMNPEBPp1pJTBx6D51R/IVLPMXGqbrmbf4PylrM1Fs1VmzP+M+j5gwIF/+XdCk
1NuFit9cS61QUQUviaE61kl6QOGzpe8hlapZvl+5rmu6E/FAAEFSdfheIxgaYTvraoRheQ9fy26U
5rMrCEQ+lmxJnqApvXN19OfuPDRsyJ94EjTfEVzeRjmqX6xIjEWSKRfomWzFi8FozNKxEZ9Zvaz4
oBGav0lQMpq/QyZ+b9K5Bgj0LcZPje6eylJiVqS5tmIMsmClLZotc9fYbvzy/+52wilSfPtkWlhh
PVbPfg09L76uUhXcj0m0OJ0ACU7Bkw6cTqInHVxwIKoqTz7TY0SIRiTbECrOaThw8H9tdaM2hynV
zuKg/0N9Tx8dV2bh0AWDfJBBfk7xL0EJg8x47QzJP55aIXeelMUar8rIC3bAcUHN4BuJQR/mCTkV
ewGgUTFB3nuQTbVJKNjn4A0Ldu0+3eZMwO5LjVFpV/cfAlJ6oa8I3LWc5ypGONKlJIZ83+zK2Zkj
pG88E/tSU5jn7pFA/v61tXwJjD6hUV2iih5Kqut/ACpnVe6M3+cBWCMBGfiJdmxs1ZPpbDRFrC7m
N3JWSSkzkdhA+gj8yDFwUuY8H6JmXp90vMOUEO85fpSnoAqeBbDt22JT+RVyUjDAJjl7X5WXMpNm
y0owWexgWV0DKG6cL5iMN5SogpyOCqHLC/YSQ5AF3SxTRkIvdTpi/OxPFFyJBB2L4x74l95Ki486
sgtV3r652SsGU8/RqVGqgO6OQDiUTMX+6QtWvChNxqKPzMP7HAj7Teh7GrchMgRr+ekQKpnTZO7Z
nGI126L/RU/h/z7O/dgeuRWTyujDEbGh9zanHTHVZwbT8x+AwDi0WMM1vdhMBEgWuJgwVozItuqI
jFrV6TQPHUqDcXAZd17xgBHN1azrg1hCAxbYu1klQAeLHbEGffef0KCEaKqc1XcOaqYX5n30OVe9
hzMNP/Ejl/a55UBtdYQFzZNisOuw+cio1GIMzmQda/6eUS0eQ7AH6NUJ6ArotHmOqEGTg2ACMrwK
xQTnBb3hpD05tGWIojKpF/IYmJZac6GDaVHMi+2NU48W7nFU+TZttSmFXa5o6z/TcNB2FDcEjvGV
RzVffHzZpzRqdSn9gMggQdqFqxQNFTJIqxT5crcTtQFVmp36SyhAQR26aUV/r0cbX/Q7MRIHdH3c
nEX4GR3IO20fN3o1IQRtedym8yUFICfBrF3OzzqbFeKN+/tcz54OkRNaa7FKXZm6gpE/+r1tnUKU
0S3058sYxJ0wRMvRD5RIBETPI4s4YkWt5SojZDviP+we7JjYrj1zSl5ZeFltO/T1BJrFDia3Bvfz
JNCTPFuo+eddX+2U2aOoK0r9dtzf80CmaCISRcbSfE2w5KL/c69N4cjiXPtJJFdC6eBgOzpEPP5G
QQjYh3e9cgKxJM5+845UW3mQhSMHGuQWFhPpCC82FL2CYPfaRmO9yLmP2u/gidXjfWYZaOfw7rZF
KMm1nUPDOdOP8vbOuA6oAMwdeLFDEIf2UxvKjOiMqnoLpbgtbnyiXvowiVbm5Cp+fDgYGk/URH4+
un84q4qTTjfzV/4fB/i2Gkq/BgNIOUCbLJEiTz77Gp1NXQHxXAqK21rI0TrVhHOqqjClal5xG51P
98o4k6s30ljRlXQmhtbcobFTiU/1tk12aDxW26if0+1QPK2fgSvykho2ebZuj1ZbMwVapm+cVTy+
NLtaCb4jz6KoueY1QctgilOsvcwXK6/GMUkoF7qwDEMaNE/zd/KjNrNmEuF8U7LxGkmYo9HYWqnW
hLvgmtVzGbrFxF8rwJYFBwXo1h3qLthuJ1iLsSwwzvq552pGhoY4TnsBjKsFppPGKEdtwkCJqiAL
n3kFw3+M8rPSFEZSBpXDaoT68x/iqrxN8Rx6fHnewSI3pu7TVwN+kJfh+zAt7EAcxuJQClGy9+hQ
SHrtt+iKEkdXXSJuGeSqzJeiRv9wVr4ea6ps86F3dZeOi/2ZVoNbBA83EEqXb0WvumCzVg9gbyvf
oqSS6KLUQY7nfgXTElcWefIMAInIKBUVCRBU6tT6JrUrZOBm4fTlNmWPgLiewTboZS+no0krZ0ed
ehw/riopf2rwwcsv+7F0yXCNdAkTPxoYHoXaXLfjEfvJc/gRxIQyZAcEioCg2mE12sILiNIoLTPi
GXplDE6Hc3AcNYTEAxspbo2qZcS1foWxAA1P76CedPuahIeOO6XXY+sQw0ur2DiCbGL24rUf/I1t
pL56wyY26MEUBNRjOm83PJIfv+tqLCo0cPSl08EJ2HEFCEpjsdQij7vxI7qUZwFx3eC2HlzZcr/c
7AHCxt49iKSJsRS2MmRDdU/uKGKtQ/dS4ePNUZqGQHeSWDarN+rFQExdqZoPaMUwDBdvjn8YbTYg
PTr7/xJSwAFnzQk6mObrNy2NtgS5z/5cP2YSbyPykzELrJ6UbLPD9hACtmm8vp9pZROWY1phLk8N
t6QJmd4fe491+jzGRHT5cWLGVfrUF9wd2ftPkigQYhlbkRfu5/LW7YiKh4nFzPrEkMkb/ERmPKDr
w9Zv/T7JzSiz0kmoqN6SOav0WA6t20VP/alYu/t8nhIXiUWJ9Y6y7lUs4dXv73z8HibeeWs0qqF3
eA8ppn2XXO5LXx2UVhkDwn5n8/euXKt+x4IpSAix7eAoV9E4/WsTG5VyBq/TEVSY8F14GNHDgBxM
6dBynGTngOHxeLUT09yi93KNdOWw/sSQ1ttzdSdQHubGYtU6lI6OfG/iuPg2HdoCxUpDoBC/Jyy/
UgpeFzfcX4dR0RxzXXM06ObLXah/QImKIY3tTud3OnX7jMFcPbsvEo3I3MMgovrVLyxektGOACg0
BcFSxs13xQcxb095fD7/RsMVRhBHaJmyf8PYEv6r55sDZ8Ys787anJR8Xqw4Cn2CmLOGbPnibc4/
oudP98BxQL1DB9n3DILsrWae2Mf0xkM4VMLOX6pyFDvgDjYZ5+fdzpTM/Ucy0DU+jY70YnZope/y
h1VyoFcyvby7aRTnRpxV9w7lcQLZxBY9dWljRo3apQ5IbAINUWervAEyqQPW5f3anw3lOFpNkSXe
bmgVXobaVjSfZWkTmCxpdKvfLYPNv9szY0mGLlld51Ml/qwj2TTDIT7VnxMeyjQUloLZ64VTjBXU
uxtYOdwz9xuSMvfKTaxlcbCy84U/gwlRmVv+CctB9iJMOnKgYaA4TxIQfj+tQVsaIJTtjExTRyrn
R5KvjSp7I21iExnCQ7Pm1gFLcGigeF8UKZwyZk5GxYBqpydAkPEJpuI31INsCkNKE/syaeE/GnWo
BfNh8wpamMHnQVaNssfATN0guUS6+r/u4tRoAvLgDWek1TDmkl9n/jj2FVZ4cm4mg64kkmzvu5BZ
CWL3PtHGTk8Qkkz16Lu7bLXNxLjNUHLT04tyvQq4HBa/HdnEWdFMAEkx9hQRr5+AqTNi+QVro+GS
4QH0Ibq5MrgarO3Py7wemryMDc9obrjVp4ll6AASnJH1eoc5zy2UcwdsdamzFey4x1ZD9XdKfMf7
XCSr5+GYPN61ZZX1cuOi723IZHzGj4LzDIJnEpaGUEGxlm4YuhQdRs5xVaknvgdBlqQFyy74YXxC
gzqQ1yMUdfwkxtgHqkusbxzfAO6Lf0Y0cLDS7y5IfJ7LDrjourotWmRcJxuY6WBIwo/NGkq6ASHY
pAcr4gXfalIBgt7Jcu+KrmiK0RKj2sj9in33Ec8PeQ7C3jkVzGDL/fLQ+GC9xMjnEm8jZn7GopxE
/kKq5kVZicWFMz6zyptvoi0u0T+uw8qxWa/yQuQbmRVBB3uhwFtcx11F8qXh1/x4Pr0XxqIEwRkP
rC8B4/xtn2gsLcbBYiazZeqHRqtchRcBU2JlOH1VDiY1mjznkNMynubknRPBH7q8DaFf/rOToYHH
9z+XwbgsxGLQ8XqtVv78WYfaLNvPYeVsUgW54khM/t1P6L4mcicAXN6KlerNCaXyzXnJ7xe3HcGU
WlCpMmq4X+nPmOiTmXDCEUUKZUk8+EXqVdxxuUtWdBMBVZkT9DiVErGv8Nff+w6GMdhsUWDYaqJJ
1z91+yrgYH4QtgpBBq0RHEVLItRE7+Gz0+OQ/5rmBJd34Tqy8MhewEp2nvdYZ/W5joepXGDouZ41
q8QaTC0pFr44zz+4V5qoIiRNKTtGYLgikAw/MzqZspXaPn1iLXwkRklKbsI9qIl1TxNjX+CJx9mW
NSx42Obc1jmxP5vqtbk+9B7NES59NWx7ms7B/JgUlVIyDX8nN/wRjZStTU6Yu6NpeBjsPkVWaWW1
H/rhUYFfmArcVnql4R7K1s3LG7NIMnI9LaFrbhyklXrYBUU8T5JtUnMjcvguKNzv8Q61p9prrSs5
S8hmC6d2d4xEIGo9Chi6BGDJVu35XeDlNZwSwvWgMjpxPdVR4w4/AfTkpTeOoR1BZXxeJrXDNpR6
Ryj9oE3gurQ4VcCRGFuZD42lWci9fI9X52635lSgOlVkdNpz42jij8xnv9G8fEu0NzwtZ3Wy/RwI
DNx4w2YGGFmaIsb+rizYRgqoMaj1bo9qbrpytgIYR17YzYFeqtAK18vYmYfpWqUcz2uEW79pWSEe
uTqEAV++6E8hrhr+7ZzcK+YQ6xxziTlJoQifnJRmGhTelovr2lZxlYkLJxsgUw2jTSqmbWKL7Gwv
dy+Ui6wtpsjTzaRJqrydrb+Pr55OnJkWO0/oeJTfR7eIleUb32MqHX2lQSpIIoV2Ei/ysupIN22g
B980cXn8RfIium8LU+BKBCjW43zunRjG+invGkbmKg/IgMCV8nbxWbLcXmxkZ9M9zUyDhxqd6N/S
CqPxeH3pzDr+vkBYHnzI+QlIXNzURz3VdLH1aGeRd7nDQYiBPTzz8ZriFYMUsmFlgPFLKk3ugA9R
P72r0f0eq5Kpu6btOecocd35zNamtjqD0FT+CURTDMkmZx+0PDRW/zR82UCP8Pol7FiSu/xfdonN
vjNxH5QOOUr+cyjJ5k5L7GXicZebDg/u1dqgB2PfOyqmqYzFXVivU4K1yq+ge7SJjvlv5Ht1MoH4
W5LQrYFfyKR2kDMSVi5SBXw7q57AxB5F2E7JY+SfatCqDUOcvqsm+Jx6BL3Bz/oZ/QosGhjS249l
t4PbGmUxTMdFuRMD41VkKx4DKPxIlqQbTST4KUFSKnll6ie2ZS+pYbCsbVufue4SqBU1ZDgyQ2RR
OptyeKvjHWaBuQrTBlQTvrlSgDC4mgJfEoDklpmlE9j1dGymiGIunKMpgsgq6667WXL0KdFLdYnP
s0tegYgv9eBB6okkBaxIKbqhWafijLBpQvupnp6ZrEWpNNZTy9pk326Y97E0qOAfKdca8dHTOJQ4
jVonIxI96Z3IK+FmpAnShKokQYxtGL0g3EEEPbe9FVX7rdIs2D7zIuXiGyzUiN7cWmPUMyw6jaQh
ukF/9OSvx/b7sDWrsaWDydV8ikuH8eJ97RVLJKtrYZwOFFp2jwWGdrmVJJ2uXV+d+AOnEtFm2byE
0gRSCdl/at8MB9+fQIMDDpqDNNYgDg6FtWGRzjx+xrEJE47xOGYhAfaAhPaFgAoiqgfiJWizmhSO
wBJAPhQJXZdL1bx4s5XAF0MvDEKTS2/3SaROfYtRiMFcah9uUsxE5S8DrXUZ6zeyhDH8RmxMn2B8
Ik8hRggY2yKCgqVARqJyYFq5L0JNUIJTAzBepS+s93qdmksInoFy+LgzIRDPAT26c26oWQ6ehfBR
tkTPy7nI0ddozYn3U3x1kZ62IPQBfUDpb4xkdeAjixdXzqVenZz3rnB03ivwuTWWk8XfNPHxTGoW
6PT9gbL56QwishU8EqCqfBEL1u0hUzALnx+c2Vi7hBVrwQ7iArUYQHoHhmWUb8WqqOUVAOgW6b72
oed9ap0TWP15xgUQVv8M/0FZGLl2PekDxL7cmfO9Xd65vhSCf0R52aL1MsSSrcyrkQiH3ZPz4gAJ
RxpSu7XNozphhgrGRiFU5ootmEMTOjpznqyOFFS49obHU2oGrfpRX+1koYTblY0Vg4htnOwNeP/7
bfq5E90Yl3MW1TSSXk8wqv9XOVRmsZaE+q9AVtCQkuweC9eFFw3L9xkmHnq1TfDpejoSQZKpX8am
zHhwO5eCMQfUiuggSkYJ+VlgV0VrN2Le6fer/jrv+FwIIBHZDMLXAwCYN+o8doo8PfSmm/WN/oTk
3SR4vyoRIO/PXXuuo8mJQMpMwPxDG7H7obKJ526gs/DRSyjtBOmoWtKpzd9+fk5PuE1AvGECANEn
yKxpMd7KZSbF5niZJZgq5nwoVxUuBWLjzx9g8sUiFS5T5C0N3Sy4ye1Ex1wwweiJijkdkeGjVBVn
ttwqZ7LlXPfATP35LDp8FiB9LqUANu8CLobBy/kxJOIviYVllyERUyV4a5MsQuP5WqoHopUgrpAV
g44/4Qm9W+HmBof7FVcX863QMuP66jgu7f36Y3RP+E2u8bj43PKNkMcEmCxnfgz0EqmPGFQlT8zy
S+Q33FEw6aMf9TUcSjEnbGfkbexB0MboBBSseYQuqJ0CzVHXgfpW3ooM7byObPEnZGDpz+escLrP
xbOzuYo4oFVlljMA9DawNnzzMMV8XSUNDRV3WFHW6TJJYqEqKHbevZnr8/e7Ny6wD24FcrxTMQkO
FqXVNtmSy+dSK3HMPEx261pYZf9u3K6JisYd7wwyZVYnImIZJe8hJOHtzdOq9BfXPOY41lxGtCvF
ihXnccGYNM/VU52G7yAlLXizEeKfUyird6zUL2bwf64wNZ4diyG+cmCjsy/DBUhZK192l0VyzyPn
umAN96Dkp5PZltnsGtgeHVE0r8Q2RjOgUI7AtTZNqhqq6m62xr+lyUAZje0MKUL4XS/y67zmGuwB
DHH3xhPzp2v+F5BW0BYkhMUj7SY7AcjAm6XyW8ldnP8dbcn+08Ynpl+dIrQPF58/6ZHFa+CO0j8m
hnXJrQS54w/yU8E+CHu50a53w2gwdAHspQNpqndsZnO0gNHZGgogNQlyLoclEooUAGPNflpYMkp+
THm4TI055jZfBt+u/2A8L8BUg+ABAgS4WkV9buSDdm2Z0TMK/FF9IYcR49vfKqQekgazx5JPcMt6
H2UEqjETUUUfPMro3M6igHJ1eBj1osmCnkuumqW+EGHMVVFroNH2bQQN1xHTMM5m8rNTvjHyhWFA
8XHcIFrbQ4rIo7Fj1qV/1cY1zSjCGBAhSpxVKGsasB8/XFjskC2aZ3YiUWILNHDIvEAX0q3LO9x1
Nj477UVjhWE/LYo5lq/Fkp4vWacas92UhqIDCibTLQOhErRwaN1BBaGul1XeW3v7qsgspk6d9yC1
9F0kEcaaGgt9xsz/ZL7+B594J+K08LLPFGcKO2mZJR03K0qmYE8I384QjJsfSZDxBx0f0kxuT2sO
Vib11v1Ts4EC+FG0ccNz71epvh/A/i610k8bdX7Fmw1Ub5CD8MZnsz38v1/msW2jqOXv8NBRyp37
Pg9f3/0vs4XZioYJJMpVDO/RBHWdsD+qU+uI3j8/X9aWcIqoxKz6uryOZuRK8oX6XPh6zcfYH2hJ
dG3DPkDUAHTY4mGDcTT3tlXnspGmEk+tqZYCizWxSh9SqVpiLXnUtQ0/lSRdKC3Xvbxcsx/O53us
+9zgXSEHkVzvqWXr5SH/h+JkpK2XdD/a4BA1forADshVWrqHwHVboIG46pBUgL6MypHq/ZagtoEZ
A+C7NbFJFgaIjI/fxq9DxW42mtgyXu2t/Gj293MOJxNLQCcAqa14Do5XbJb93WVe8H3m1pyqCbc+
W5meFltek1re5uPVXNkN84jB6EAGKp3hkcq1iOlzt/SyiQPM9pDYSPApfGeHKoBjSuoOXE93Tl/4
ee9v5cFAHHhboNnIn912xCT2OdEvSdng9M4qDpXHYgCHCMliFLTBss7JiPTCag8Ppg4DpQBdy96u
14ROVadi6RFucQ5Xuc10Dd3OSp1uKI8XEEvC7poDKD73AIVt8uZAZSiZWLomKiAB9Mm5CLG7/WpQ
5PST73VlKn3+Glbf/2rh7oX166vZi2bsm6m8QVmYQV/1cnB1RdHnLLKnjLyDNc23UkLiJnuaFfqj
Coq279ALYAmKw4EiS58/LrXLqkloUTfSRfvJjfI0PpE5mcbCN5T5qEyZruJfzmtPNc85w8SOKZOl
WT53dl4iOx8qQXlugBAaZ4gsL0UkzS+LEPKEyRc5swpXFg1t999YUCIosWmgUEfApmrNE6EL5P1i
29wA3C6AWTT27XJL8vw4yigmdDG9MlylDuCatJxwh9nnR5t0Jwn8pWWC9tWF0VPgPj8v1YOm3Myq
w3QUf3WHzSpYKLZhfqlXtNTMJT+X4EqmZLvCxFnH7k+b0Ihnd/qAmwa/sQjx10e0S7yvk0rUqnZs
3uoU2FHrbK/6cVVnR/QgzlAADqqBOqB4kHej9LIXNl0UqwK2lKCu9icUcafIdGn7moh1mveyI40q
rMpCzVcU+WflY2LwkDNm9DtXiGjdjYWxlo1z98dRp3k+65rZviQxyNHtfGttyydMqm/HhHNbI1MA
jiKmC939lQOCJLyHS+wbHaapQA/Xz4PQydHaTqmv1cJ23xkF8tLr1GuQYZmcx9dNY9ZHBmDYYwoB
oOC8yXFKzjgbf8vCy16/rQIQ4qm/BffBtfibiTiFweNdc8yWpyIgKJr85cNMNk6yKYzI4AFYNn/K
zF4iOeZ3RPwLpZyx3fyZ41abN2Ms94IVjDnDB8jNtwfW/xhHtVdqU/Q+0b+jchD0OVS4SqAAQC2g
RqXdeFH3jT2UCw27TS7LrG2VkRDOIEL/Sr9sX0Qpik2kk76ZszzMRnsWce0W/xu3nAB0U47T8cQp
VHW2U7LIEnznA6woRIZyCajkFmnueskcH4A5jK+x00BEMbdN4yLFZiwWrOyROg9PetlN13A9rYzQ
Rpc+CX0k/VMEO+AeK1IhAoo7NcmLeMb9rsABkISqZeuE7seFM1PocDTmt/p7/uyLTxnGSssiuxZS
myFQiFNpbEBPnL7STXBBjma0mz3cZSfHfJJB05fKUr96ohlj8PWhgHpwvvYiW/2iFdWlUmIa/Ftl
p9wN6o5AbWFN2GcM/Gx/4GZr+Qt2Cknny5Kt+vaSTUPABDaAwzhgcvFI2ieoB5ZRtj27UQDkl95Y
+iU9j5TFQWf0pBEcHMyujGMcUyx/nsFj21xSNXQnOx2xAjLJ9oZasy18RRouOIESkhptCwcHaxSj
ZvQkFi8guh8yItr1ipFYyMqRfPaXDz0pTLTGXcZA06tYptwUm3DYJxDpZIm/w0HejXdyA64XzH06
u+30qWhHW0wSuh7ScWgAI4VaO29DHJodxZCtkNzgMsrJsWeDDWeT8SnEyifbWVbJR1lASXlSSSvF
4ARszRbtWBxubnB21+hk8YoOZPm0DzG/K3sw+BvSubMUtoDW1G7vK1EOXEpTVilQu5R6ZsHdjCOa
lzCc8eF6cML5MHVAkKTYZNGNDi3ilJH8nCYpq7d4h/iTfoX77sjhblWQzvnvWufAlXpg2dkIA7nO
DplrJb2wUiaFBOUhJxxTL15t6bIW9yPGkSgCoe8T6n0S0moK4YxIAlBXY/tXGAkojRVfRydjpsp6
9lDMAsclOY2ukK0vfpW6b+jCj24Ip7bh+zUvl/lLRaZa8uk64Fs9haBNzwdxi/qI+zbWDZePjPBw
FHoF3jxHzTY2v3ExFcS+DqaGgq72uXvmlhcc507FfICNmGPIRCPcOOvzzFApIdlvxhD0SMQW0gIo
X1MQufSCMWg/TPc9xzQ4U9Poh+vvjT2Co2Bo1DMxLn5hvURvsbIqY42XVKdnbP7Ke1pM1pCzAUdV
CdWVXEWA9HfwfEu41kJ2hYViy2vGZ010GqjdvF0djgWipUfdQ45vsxCORG/uP68sEIyJNPhW10LB
BnRZazjvUKUY2R/jC9rMIky9xc/jdHb+HHeQhU6fib4qLXCUA5+kNsF+5+GubjdEsOt/PfKRUB/9
l+yaO/b5QOp5RtgHOQ/pBn5g2cZya/Mos7BLclsizdbE9bLUR2xuAIfUcDMY+gjMX/hbm/i+m4H5
QDwUTIBoX6WAP+QAqM3krge8KjwkhyzHqs/ctts6/2rjIjfJBZkqJ/lD1VtPlDMGCdLPHKOyrxOI
mcIyKe2B9M+UFzAE/fGjAee1W7nlzUM6H4EudF00fK5MnwKk8xRsE7RIMh3+XBO6tbHEZOcM81VA
CWMYDb+5VmYgY2TjDOiRwQ6HhcBRHRMSsLRu4ZM5x75YNytDbcoKEkQtBy8vN9s4ZqDQa57OIoYF
+f+Aygh6qCD93qruRgv09nXCLVlWcQ0idtP5/CZRAiKEziowp91AdqdM0k/nIzl6HYLEK2bZbcHk
o2hcufzQ0ZDe37vbGbZFCv61Fu0zNFNGZya0X+pSpEsJcDdnGvPfIlzlGj0B+OYnaP6F81d/87iI
xx8AJfyCullgrVI2JUMHudgfA+lbc75Fjv7ZBCJdQzoDu0VHwkoRbkzuYI98ivsw0/s0FXo+zqV3
fcvFOfJAVAdEkIVNMgveKmETJFdebSnNEU/BbhP6MRseLjytiXf/y+oLHspehIVBO9RmYJ672dcD
74SdJPQxwU4TE9tu/kTI4QKxp5IItEQiDjnZaWclx72xyXfFIQRn1ACgmQAWCnCn7fY88s7+8qSo
KVjRelEUi4QK2VVHDavF44TFWxMW0e50cGJxoI2DFT2HlKwbxJuy1y6oTcrkwuh2fxEmeFQahvmQ
EQRQSYIBWSEdy/xEhad+cUytzIGj04kHO3T0tft0anISs9i+Jlm2qhLaFFeI5k9LtoqeUL4GuH87
T9vWWjB8FZQ580VNfo2E4i4W4EdGWnP8NtFQS4DoFWxUBf1UQcjAnKTfqYfOjYyfNkCStqld1u5P
B7lG9ZInc0UoHU1aZme6i4cf4L+R6G1mYtCfDXXBtbPho1Z01roQx18MY3hlO8cH0hcrvHBRw8Ic
PnSLY1Xr5OCjeHzJ39m+692L9Vrs/SOLNSVlPov6OWY2+ElE6kP2Kui02Bz18a07CaWLrwhIFBya
/5S5Wbj4xRc2OXkcEeylwTGji6Du4yY4Wgkj8qBP8tMG+NDdqFQaAtK46r9+aVEQDObYXbVUgm2m
8OLT5i8RuCebIXEdVtF+fGVDZQbtLQNQVol0/AL+ZjG5hbisCSWoPoHF4By7Q3lTSvTG0IskhKL2
BNMvAH0mAlANzTMkQHeBP6hXp46Qmyoto6WWKnloY8gQnHA+gni7aKXTv1mtU5GAyFdTKUIV8eRd
p4XDk3fd+farLAIzPlIZKqxLIGs7eEnYP4ngY5CXbYIRZPcGeCF9JGm7DnrjOqI/+GS0/Sw5LoM8
rG6RVsNSW7bS7BijYdZk2BZYjAcUj0qfAXsUx9Os02kBES41MwoJyTeeOWu+aIqxb/WRFHcGg1P6
EDDR+I4gi4+/kuo+Qaj1uM5OfALPK9ZVBE0rQ00g+oF958dvEEY+lnzpUxYQ9+A+9OgrXw74MPAd
wH0nwAYejrW51jGUa0Nn1Y+xIQwAFFo2F6znYJu+wwuO1Hh8V15XfHM7IalhFUUnN4Wn6xVXjap5
AC97yBkpl3u9t3/Pn52SuvFc3kV3oYAaXbtug3c8ccGQeCJTyFUOeTDoOCH0OBKKHwA5ptj7t2+x
3/Cvyo3gzAGnmNb/tQPTEHlElZplDSUTB4sA5Wg6a02QcomkOACQpKZcFc5v1gBlc7yIoz8TK7BQ
3MunZSDaE6aAwLVMxHrypDVZsf0ogAWPH3qXbEk/yeFHX7zysVAFlgpHNcNSSutlmQ7LheEfpmjP
QpNDLwXwz9flZqRrX6CEQDebJkHLnnALCi5lqRzVQ/kica5ANxqmDYUsLFKip4PQndwSbYGSm8Gu
MXVcIguTxy7Defv9Vnwf0/wfAyArGuZeScgpxl6+X81VWJFd84vwaL22HP0MxszDXa5CfzfBnFlg
eD6lQaj7c70xyjKVxtajungBU4fuGCEjToRazCmvnys5rxWN/30YTENgaO4o7Y2CM97sq0F9tHBj
kbEdhsOgW0k/TheG3A4sGTI+mq9kFGi37gqI203Yi8ecODoZRRZ5DBb/0POL0/DzeI3An4aVDp9Q
fo4q/iut21/fbQF64ycNp7hQQX4Xvz97mkVA5bDlkiNA96qqF+0csGLNyOWpbG3YuO+xJZPpdx1W
NqKDcRZLau5mTY3kCrAPeejXqohMGJXNLqK0wfT++meL9dIPEZTbjyONQ60sxEiZAmlJzoOgsQYt
JFik1ioO+EK5tGsvDNjnUufCB5I/j1/G9UwauwLDwCPEPorjF/nd7E7zT8Oca5ReAKRN4nnr5P8Q
a6gslPZocbH13ZKrIv7RFGrjZWWuZJ/ziArh9iIAQjihZmVoTcLJqvJs5JPqrZ6df3AoyIuNLUID
7Rj7x8+t0F/ogglQtbKN2NwupgAdSoheB8hFZw0N2S5NQAUNmCVsz2gbRJI/1egaqNzzs9WEY+Oi
cA9ugHFhchvuWcAlQSfhMlrAd9ylycl6Rj63dHMUSVvb2MZ5hoRFir12Yn4XNosnzEFkezeToCjW
/MUPbZ3urCvLz+h+UQidqPhMOTaCztqtSTrsWhIYnJ8omjyRCzlbcufpOAejSMteVgfOAfQAhEM5
BsUKui1O+om9ghm51zAgt4zf8H5oxghNuohDo/4MbTb9yNFcQsSuT3T4cIAGIjUf5E3SXqVGPGix
QIgCc+aA0F3TciRd5CxKfXEEqMKxu6/93nkozlKA0nHlCdmE2gszDubDxyjRWCV8Ge34hF7Aacty
1tvINegiVGFLdWMAGt/NGNOYcjiO2qN+A4f/YIDUdw3MwuBfKFkE4BUrZCuzducpLydRE5pDEcmg
kkKOgx8kNpFy1qyAWGtnX3pmg0HLxTVyJMOtIEz5oRioG1dGMcm/Y82Tja2QCi69PLXdNFrKikm+
mmb3+vP2i2wcK9p0JSAce2Y8iVbCvkdQPSvUuG3M8fHGvJuxYVNng0oBvveGm5lCIKYRTK8r/rvT
7HQ9KFK9Os3KDzj6iBh/Q+5MrANgNQ8fRaAaqNy/mzHPKsQMk7fOTfpQ7mTopa+pJ3KL+A6Lsm4i
Kdtwd+OGnICvshmnEi8dQ5xEuJp8cBRx95Pz+5q2r2YA36tvrcDiRFOylLWUFpG4zohlSlmtyy/V
RpVlDaYI/d+DmLJNu+vkp7ml5EHYY4iG02mnKFBlDiHbd33h7N+rIJZj8zxrRIzyC6/JIo7DiLDZ
MuVNTFOC3Kb9T8mbLThTzNYD8+c2v8NjpKcefKW5UhJxg232DEASa8S9R+eNW316O9yaZLUu6vie
haa2fN7LoLpG42p4L14a4+RVw+ozhrgKOhSX0UwaSTB/YEL/ZR2Jdm54KmZCkx18pVMcFBbHEpVn
Jb84wBNcuxRdLMJf8WjLwGEJFzqOsQ4iapuZV/6sRk4PLtxqrHap/pC43orNq4RNqLbv9NDW2ecB
/nqVMum7m/uaYWXVcTjJd8Zy+YX/TNo8PgfJ+V4YGa6w/XCyW8Z2pDTgg9ijKRzAAoGNPsuchUEu
lah95QNrAloogCNgh7ORreTIfTeTOiDFd6VsRIsMglLD8NiX9GOlJsIq4IFDLP+anOSD6FdDxT3k
JTyhv+gnkYffIsJmSKGo1CxmcbcTnIpCwBO4XnmFButfnERry1hX6rIuslD/8w01vRtoPY3H6e12
ZGY+5UrOqtHKCcLdwlyInuuLWdO+ltXWNUciolRZwtdBtHpVM15pNLzVx/NxlIZMUNuM80ROW5hK
ln64EDn2Wa5QxUm+j7VZ1Q6Pr85zL6VMFRgz5ZnYy1C86ZAjNiLpignfF1zLrGcAFXFy0hSd3chs
qpzwM5x8pKkabSdI54CE8wU7K/Th54ImvyhM3SXU5ylvZOjSmxtmshH8Wmsul8c4RjRreh3R+8BW
+W5+c2qcAwZrFcxYuC0Ml71RvHUKyhz/GcZL3mszyrvRkLX3INLcPX4Dww1OZibOM+VLnPumFkmC
DrrhYUOKTiIQby49+KRzvo/KtZzOdHFiZFTvPv5j2UVCWG+8reR+BgaHsllI5JcIiPuD7OZ7nxIj
v1iOvjhij2cwAxwfMv1j5EXuCv/fg9a6mt+FXteookLp9jTQpJs0Fk/L4ATj2U7pgkTsrvNUzfMt
TmLWz2MXBt4eAJ4RcvaGuSUndQoHjh/ig9J9TtgCX04mvdiNAhXf24WPdh3VSpTZQZYtwS0wGue4
rl2k0C2vqDWX2+VxOJEcwwIXOi5h/+bXFULJGHrbj+0vp+rRnQA14LBM/tIVPNe1X2dWvZhX+S04
stZ/fgT2N+oJMd9k6Hc8HG5j/jb5sXyz+E5V2+GL0jcGpEVtnHS8W/EEuIKDT0QCUjcvY7GlC/u7
8BKt79qq2jh8pXp2Uxnklwt9YmARZBoKl22gxKt7wBTJvZtVBUI2/qeYpSLz+eynrR8w/tL8u537
UyOoouB9mv3ADmqiy+/xvUHNN7NQRNZR/SIU9U2sGZ7SulvFMLSIurkBNVTvhqJrOPpGT3lQoKKV
ncsC8xRCyIF9RCYR2v5NzMV8YLiO+Xu9esyk9q6FVgtm3DX64whFd9XOgymwIKVrgFEJjjcxXAh1
WvauGx8iHVR5mJt8xnw5K7gwXQ6b7AydvPv/4zoGT9fqpzMKr2ffKN+EAhkVkeGMyvhvlN0VixBQ
+jK1vWa+zgaffQZuRn53hlOZ685vqSMxfEq1B/89ImoQogDpaHKYDiQRuNjwJpoPnum4lIzy/NWr
7NE3Ne1CEERHXtUMMcNWdRmOG2t1dQRavuKWwelNXTwtnnWK1BBIhGTZfPEq7h9lrC9SJsnSsYYT
3dNrv8uzjo290hjjGr5HFapU+vEtvCMWcjbOlTS/GrsuIu5Tk9x1eUieA2BnLeTvQpY5bi1IKHGz
lqNHBxoK9uJCWhcEn1qaLj4qrCbiFlYy57H0eolURPRYTTi457wAeLIefhhoWZ+qMxnnlQal+EVS
c2UuN0NazIuAc9EbTiJ+7cGjF0s4M4aHPtMa6xXHWaeNFFDJxtjViLMjZMg5n9ZoKW8734GmcI54
bXYRZBezHuDQuNxjclxKU7jA/ZbfnGedyvXcWgDahFxR2XuHtTQ8th7kxVKByrxPDHmmaH4LI9pa
o70ziX/8o07uSwfS7P+tARZMrOpljnJcJ0zKlqVq8Sn0re29fCcQ2mv/Y+yzNYf1qP/JlFmmL8us
yrdNZBWGg67642zbdFwsfpwXbYYsp6BnvkFH+OGIXjfO1MDeeC+XyMrldzoywRGm3fYa6JrMwqSV
k5rN+bSjuVYjL+sgWzMfflMKPaJzlVwKmcSKwAlJDWMBKSO7rNTqzc9or+zpZQUFlr/8ziVbwBLM
38PFeUwy6PSKNQ/5UjT4edIgP+hekrYNY7WAfj0G15ouwguqmmTVcof/i2i9UnuQqHMGkj9AEa2X
whTH8WxT4OKKsF0nCxkFq2xS5e6Yaf/JoTagDzAPe+g7D+o6OvMOSnRMe2hE7J5kHrgHPT6fZHQS
KN04eFZcvZmZPzLAyjwfs7xSJzHhYEygHRkP3h9liqfuaNwQYqzK3m7RekpZX6p1iTYQBrSb4OVN
IcwoGTEXtuMH8hQpj/+jZ82aZVUhyUqWnSCSvZntGxcjjcWu74rsy6s5UqLoGXtcKpwVwe7p1NsY
GXzssvv7QA64Ufujbj999srnn8UZYbI3AoRkCqxQDcPKr88JzINL1bRY5026+a/Diz7fFkXZonE2
wpc5M3ctRVzIS/ak1QFgQILp8QV7f7bvUVfc1jaXdZnTgprif7g6ywee3N0G8lTNi/ZFDM/rZxhL
jud36Saf7AGNwL3MZbBzjT3FsACH735s3ca/E76pVV7VxgzMx/YPwaU/M7+xnCfYosecdTxFze/t
Z8SXF5LxYbEICO1UE26hfWeNIVuPEzgdgDS/2ZreEVJxgOwN4vhNrU59rfD9AL1P2x/xAhGFtMZn
Lnsi4PGN8UYSKvxgwRWbAFRWWAIyHtG4ZNpBAwTO1ISDe2ObXHkoebSkpqqsFZx4YBv0QxSaSByk
hTu0rzxITPdI7jiDusYNm8XfPhzZhmE1PdzBZuxEvszBtRNDvt3RW4cesj/qn0Q65k2xBCup9G7I
rI4X5PHToDiYIfUHiXADFfri9WFrxbUuNPfk7Sne7QsbU5a+SQDOVJS3+II/fWvjnW/Ev45pVQ+v
kcpIVyHVsnlgLGe6ooT0gpDDUDYlaK16Tuc4X8MN7JAJZv5GsUcBO3IfkJSMU71VLigw+bRJPNIf
O23DFyw++gc+4DSvkLEovhTPlt2wpl4+9Hksj/RvnRS+5H4AEUlKVc1hhjBq3mmA0EZdDx0uIOw5
BDaW1cEgBPZ9itdDpSjlu0yr9NdLk8Ru4W1rqSuRngYeTkdxGflqfLiMwVcl/OgA39dphQZE31OT
kbvrtKyH+35ScSvTZh6RM7zV7zHrX8qDtgFAjJHFD6DNkP5JYm/QtxoqUHEYfLrg+C1T+6cE0CvB
WUyg4WH7X8rEHna6GEKJeftM2D3boyevIfHFBqmjRfnSn8742x3JkOKH2jR42djnhOOvJiFwB4VR
h2CTIKHxd1+qTbcBHlr5GplvOBN9YHGcXVp0jVzlYqPg3A3vFqpaIgXkRREaMPtk6fagy0bKJpQ3
HT2zvbB2CjYlpErJLbGs2ouJ31QY5rEgW0Zkcii4nW4YTvusYTZkxJPS6kOJ1DUYknqoknd5Sr+O
en2XXSJdNW7LDgQRSV7Q1UyHCt2omfA4+wRrX7NqNGX3YoKfIh7D9BvlZF3GCvF9Q9KRA6sz1A0C
jhX123rbF7gG0vgEfEA/hrQIV3uh4oBsbPpbe6iic52fM0xrEXcz7DdqJg9yh/xHIgy/bArjmDpF
PqIuOo5629IcE8fH1oP+0ToN4rzLij+jUpTViHs+pTVJJlMZ28OQU4fP8oSqK6Ebuj2IVonrV+Xq
NvirV7HPKZFNjf2L/kjgQ/g3c/wQwg6qDoJnCtflOQ+6YRYuO38HXwVPHhvUUH5HKxKRXYf8DMJ8
OkisnV+yr7oZw5viodCX+D1nXv9pltkF5YaOhaoaKuOqvoAx/km7fhfMxlt4rNQiH4jZ7aimx66c
kch5OW3OhQwHkzaXGSVbx381yEPQr9zi8NzjBlKAH1362Us/v7HuvQZcx/amGgXcYe1XO3LMq2CN
/18PNkH6WYypzHrIPv1ZvLtgrxXl+Lw110EblXt086KQQr5Y5ihxrcIUKNThxSa5sySDmhcjuG8U
GOSeGXRbnikyp5gNz6qOFdaCOpy6uCTX9euwsVkX46ktXAI4x8SQYz4fqmWFbKSIziLsODK2GTn4
Fms+sXFB38QPZMjyc0Rs8ofLbi6VXzbbCmcf+IzM5VeqzAYEEZiyKVkbKGjb1lPvOYO4MOnyIxky
A7Vr8O3O/NpnJJo4Sl7akr9/UsDhPuPBqtYvgtywo9NyqWjStC8QU4ElX3WFkb0g9+28exUKMq59
3v/rURavE2MTmfiyURzL3+1m7nTqAN4tbTWvx7CKcwpH39uC8oyZ8CatoCQroLGKb9O3PayGuiIK
jIqTPAzrrLN5gz1f2c4Gqa4jf9P7CCv39n1L2nPHwvN5BZagu6iY0fJqLAuKaHEaADMbW9HBNd04
XgD92lU6vbOsZyeZg2SngnN4Ast7Ki4vN+lCtnJqr2CQrBhpv1fQCzl/GowE3x03TNzeE+B6tZiJ
OEtTnUlrOmxY7xn3Tp/gjFMFyltj6sNHHQaOIYO5fCENUlDJXIE965/v5/V8gbKEXZAzRgMaRYeq
B1AYn/RKJ0U8cjhm8m2hTTTtQP1qBqbVBUtLy9IKL1sVSKXFbwMLncWdBwciDpRwL6lmdFSW4Wum
5Z66eBwCvPI99qbgXqvVRHf+suGNfXQ/LS0fTEZYcz/KycA803Gm5aIRzbpQw48IuCVB08pnlGTH
sCMpJxtwmbXKfffyfJI3ynvD6DuwBRG5urg/uoRtxP7GvITbDhtiHcY9xi43kNNd5NP30jO0cRs3
2iIf306tQUj262Hw/wF4BoH6Ye0R32hN6AP6PNrMf2P5gZa0r6v0MKzZiWKxTk573ISWtVPlgQwg
VuRRv2BK81I6glNIuYxqivti9ycbI4JKlO7ermVKSv+z5SF7K9+oeXG1wmK6jkcAFOPsatH1W63K
1IWz2tVjq2gxNPyocQuZj/Z8skqX6XkKBaVPFFTlnIK6uTarUhO05B4ywOK9Ykv51Ylx4Ke2Buui
xA4AdTpO4JkpcaqbetjE9G6Q4ebyMc6+9Ke5EWOfotOc8FRPwq3SW/fl560qbT6gFefhV9Wior50
+ee/XGuCaYU5aQ89oJMnwwispsD44DlTi9uML+MZkFsijx7JSG5maoKYjte100HoD4h2JoZtLWGe
0HGGKfUMEeIee15+LG/UvMQZzvVtYMLfG3JHYJSpqVfM7Pa5oDpslxqutjjYEFnxdOrmlewtfcEr
n1gHm525m3612v9nm6DeLlBv4b1Jqz9vCA2yrtyJlKQCBdje+oMwFkl3arMGqnwxtp1d91diXO1Q
GF0WemZbrqDdLWw15FwKdTrVc5SCMoIjEc1w/FdlYCl0ZXrMOCFoOqQg9T+ARCQbmwucvmrQMx4V
VQ416J36x4fZ+rGwYk6/5q7Dn898BTEUo/JFimGVJv3YCIeY/9qUi5xKAn0TTfQ3lD+Twv8HNERk
zypbk2SnCjerW5tv1YN1T17SDsuW2RZvQh/jVMPqlf2m2SURKucc9YC9VL5FONbXouTabpZW1QUg
n4hfEsHh2nRFhla2gDqt0lowmrAQQvcsCUY9Ip8Ls11i1QEzNxHlOtdK4w7F4WWDtpZED8yvkwQh
ZXrQnpyEQ+wmcXEGRa+1785NHhrvs+x++IQhC9P/BCTR/XfEeUIiErFHYCXMK4BX8FLxdefmGQ6v
IPIJ5w/pLmkcDz8UioEop86QiAgc1b6iI2uKB+n+6q0fC13CeQ/cnha4RaV3qA7touU8WTWvRSGX
pTltatOFruPATOqDPjmziojgJ8YD2LFk7/N8X7h8cCUzMRFb5lXKNQV37t/n7PhU8yVdtu0+lcbp
svjQQFh3LUxsv00t0YsXrwV8d50cdUrbfiByJTsIZTzmqmddEsUMGqKrmDxXqxxSG/Zt8lvezKxs
7LzJwBVwqvTthbLS53YZa6zfzvacAUOSvfvEIFMF8gRZoSXacQi1YDcrJX5ytZhmcPkVleASM1Cq
EBPEV5mmOmt3b/aFpq5yoO9dE9FiAwomeUYpBYZ86I6OrPBRm5oK9FLKSkiq4hoqrOo6bMJqg+n8
DVV8RlKXlNcn4Tu4vTUlYNDos53DmmkRF5pl3HOFJ94P+2s45ScV+ACG5uzHtUShnM4PwUhpraI1
oVzBTaqgEijN/ihGJgvUPRiDgeBlah12XSC2TYKkG1KXyd9DIiAvsLugi0cA5uadpMMw3MoT52nT
uR+f++H1xb8N63BM1IYS/P4PrevAQYlSsLrjBmzJgKD3v6h9kHQlU8KPe7G7nZocpc0wCW6YP0pj
ZSM/cBhy6sczFVTLfdfKCwdphHrvlNS1cCP+OJzshxeJ+AzFCViYUFeUcrsUrT8ChT2U3rJUHmiL
SGrQs6yITU/scfZ0O+2q61jr5zrHBY9almzVmoGmz136vmPRuKZNwRhhvppcWbvjedXR+5/yC3DD
UyutjGuG/P5snR/GIxUawB8anRSfkDLmihEV62JiHf78uN1RqxxCG6Nne6e5jvezq3kcU2rUUNi1
Ep9MeYtZGpYQMG0k+zxpZwER17KlWtebagQvvmQ0HGm2dMmLp42fcTLAzbVXJJqxYJke1WLMda8Q
BVpFefjYDtgV4QA+uAdAmShxaRSsujMvDQktH6x9ZIlVzi1DW1rMy3MiEjES/F99U9DRKfDAvUcs
ljN03h3NuX5Xbgpgg13Na24bYScAXxAS1vw9hODcXWRQFB64prhLGgnDUdjQZSFB1ANwS/W6Q/f5
WAwDIRfxO4FNGoDimbjDa4MtY0peUQBPCXrXDkKLm2Dq4kri1PAID9Uw4np7DGEiv97purXO3n2V
5RBAoev3NsGVibIHHlnE5OgT3K/mKTPmNaRjVu+3HSvTOH8DSzvFSr0PXwyvsSnb38gg/o8Jsj2P
LquddXzjbdTiOfT2J8bH795dewQhSPOiLx6XHj84twb7ullEq5u1y1ozoB4nJMe4lUYEcJ0/Wn6N
DLClIIowWGsXRxnpDpqAG1IbeIKBJ4UwX7MTHKBrDTcFFdsIlMlAsY0dD00G82GY0XcgBpAqO67w
wGWvvjRyTjEPgrfN4NGgSk7xZIwin0C4DsHFJn93JuhzTNXpO8cxZWWfQSxQv/2ZtAeQXHqRQct2
sHAFJBEywK0Zd6UuvzaoJGM1e5qJN4cqvtxCru/kSm142cREd3mb8g0tho18MCvRy5KII7CvUU4g
cchX2ofi7ie2vN3CZr181bMyhjmHS14jOGdfWhL5gOP6etLTCqoUkofMA45f2JDUzpV5UCUDd6CL
z5ILCUVGHTDFEcXbUS70v77nAb9pvKMAjbPJbqn4lJhsvhDqKzn1NIGXYD/Q0GxohEGfF5EL60DX
mmL8O+zIxJPNl7do8gEVfWiPgDLg3kSWifSTlu/ESJd+qztJqnR2RXmO7Cm29/3N9u6lMyjDjCOE
DV9xSwlh7mSk0PlnDLR2ewSXsDISPOj+hIQ+pWQ8e4RZ92EzSDRtF+Kd1F8U2AbrnO/93ybgIEX6
pXVuHre4RsBPmTena6WaIeRQQDYSPrhe3myoOBzeJ+TWtpflFkzEA+CHJIEhVFxCpYE0WatH7wD/
OMwgggDiwdpZeD2a+X4b47y7umznCBBv+fHudWnNAx/k9sWhfW/h5j30ZXpgwEJOLT0uegp1nd8e
i75G9TS56sDyjRW0tqPPvPUIm6sbPTn5GHgHhAlq1NniieK5GmUEomBny8os3vTAsSLkQF93PGMt
gBiTt2msfpcCM1zdYjlliwRRTd+VZ6Yak5KqdXeCDyhA8Pre5MonxIWW3Gu1AIBOQduJ77cu1dYc
dpBMITIV21a14MmDrW+hzii1v7vXQnU0H8LWev/T5rBLb9gflqBroUyLlLYaAkHZGi/rUPSIQyD3
3wWKQXnF2ECIP7/+/e/GAXlJBL6D1LA2iBlQbQWyZ7UByFQDfhdmmefAwV10BaaIyBXElefX7g25
B7OuV8fndLG4mFEGSyoxaCRYOeWR7YR+CsVndMacnHejUf21JsnCSV5XCu9TpJISKiyMgd8E3HNG
Yr1dyKUn979E42wTDXeraj7IEIO97eTDbMN75w6X5LbQJaQkg71VrycuoAevuYegBpVu/xoBdAqF
W4a1MNAmnOg9gJ4psRIamFho8HDbiNTqhvfCp6gjO/qZkA6VHn4ZGbtH2KxjtoyDgYZ3APpud5bZ
7kKb9f5pzedJ0qFJYaa6pCVvPTZkKTsz3fVpmepl3yj3i9xXg/x8GhkvvGqa05HxeKqZaniDjjBO
pgQIIGl7zPq2pUmDRUSG24mV2SfQJYCr12PSXoQGOYLbYWQIcU24ZNFzTfLXI8DZbkTGq3HSlHO8
xGLjcppLoD66XpAynIVCgPJrUk8hkGRcCq3s4/IJzTwRUUcwFuvN3yqwExw1RiQpG9n26uUErWtN
MWZLvXIMjc6ZRKC6ifwMfXISRYmYL5CCiC3BIhaEhqY+EA3axhfxFZQJykPUv3OxErhvlHSqtYcU
3OMrPWf1oFNVupSz0C3t0iRSAEuSvEfM2SWy3n/A1xLufDzOQ+Uukfk+AUURauVxlHSQZFFbHULz
dn56PFdcv6Fxx87QQClKPXsjCqzIoeofWfpctORvuZuIuDBdkBcxjWoRZs8qLqv5CIwWuvrayoYs
fj6wlIMRMtybhbHJWs4g+fAn5jOxp+D6CprNzv6TDAMhhKiV4XBW1e7wULsvy6ONR/s9vlAEup71
F8U3VVKQjVS/cOBvZCo58sbE63njGdBxFdjDAGWWL7fKN5l11wXBCVebPomp+Y6/GHkdyR7qBce/
2dbGN0ScTnEl3EodHhhhm7Ax+AqaSxnKwsarWFJWiSStOZOB75eCCSlj2Jg0VHBUZ3EaWjG1CfZu
wxlq3YANN62dBKi4BKqWku9kDOyYEMT+CiDFiOoOt7r2zTWHod/47DdsWJ+4UZmYLskUXslQyCyq
ShaRAdLcGmIl8JuP0jy6vy0ZGlKWqAnrLWwS/uzaM7+j1h00dlqw05AsNgSdjtambsX7A5inkaFw
8d92D3s5A+1CqsIrZ3bJUfC/OXi/zU9/qAXzvYnIv4kmXumTyQoHlID75Fo8VhQgi4TYdTLliX53
Y0s/pkNfVG6Dj7mD68Cq1GnCtNUoRaGv+1/Fu8nXUI2VTitQ5j6+6c068MyLuuDEJ0VRQ1ukrxXz
koF4IGDjm995sOhOBrayT7kSh//65eTkJmBr6FJXwnYO7xI7YSnUMvIG14Sh82W7C+ScJP4kDbjw
cE3Ena7pOXJJdyn3N9becJJkM0ucWXPC5F2Lvg0dmYvl/iDLRsc7GpY+LcOLuZjY6QUYV+TThBsW
xgWeGOZ7J211NP0MAfydZBjEfeVU5okpTxFcxMBs8+E4nP3dnG9qxTO6rUCUqF2pES3pEPAbo7Yq
wsnBq9lae0RCisIL7Scpys9vWg9+DQAWOcVRx6QlWNbmrVHzExpp7JihDg1iD1BNCmmOmIXN2OM5
5i7h4jt8jVlRGFEdJVUe0K8fCkoK1iUzDJJY/Qrxq9tXJm1/PNXbKRBFEIf1dlJFZH+bFHh4soDd
a2Z1sLjH7V81npyv7R4ajeekVza+dYK0ivQyLksfDgyZnMN9yRchSmBJr7NW2T+jAk8U/3aJVF2Y
DNEdIxLNV4MfVjkxKAybfsc1e5A7F60Z/s7rHKlrKd2vF3JYs11QWHuXvjjBcxucaS8wNkQaSiho
IVAE096gRBpYEOPLqyxb/4g83zkLZboZrvcBzaVeq0iwSELtgMlbYs1l96dTP0LSt2gTojXI6l4T
kQoe9jfsMwla4LbgRHwKBZJim5c4EJee8nRCnKT5wfiOTYNWYJxMYaWUwE/oUl9F3OwscfGCywof
gEpaLw+v824fy+L8OcCFAxwkEVRbaILSRpnWf9VtNPtMqDsXuwUlVy7/pHiOihzIBtXgD9huKK5v
nl7voUgfidLaErMqTLJcpJLlmGSXbuUdoaOb2jUz7K7b6DMGDjBtAhr1+N/qGeukJhkaR/i/nb9P
hRBM4y936gDNTMisVEzlPx4h5LuXEvDPv4Y29kOSDzPGJxVa3/qUJe1dCyKOUcNTyvjanz+kO2by
f46YloOCjlEdNFXkLWJrRq8TUYbkthxggoCqer8Ki6Q+Dm7AiIF7vsXUB0NEaS0pYTV1fEG5gdFM
NnLmyMi/mpQobqDOHAMipZkyxlXskQ/Ruf43FSVNjR6CcWen2sjTct8ZUZviOEXuh5wCbFUd8KtZ
80oYWodzaqAPp8Dx4II1N8mtnCJFsXJnKu2FGeVI/Z+8uyTQ0HKY7hxWBDtVrsOMS3FShgGegT/y
tEnkkRNztZtCPLX7JMnuSxkVlAr6m7HQAL6cBI/qk94dt7cfnWGztAtYejyHSA8DBAhvJvuEsJor
w5jeK2fLMJDiJreizdYyTKxIpi0pdF6GrcdDCWlRhlSvR1LKO7SWcBc63IWe8o8xNl6AbKHNZrYu
fu6x1OFrcnQ/jwFvzg7p00pRV0hKUijj54yE8bLn7EBZtdoCHDffvER/+kmV7h53dEjfo0HBSclb
TQSO5tAO0bIxt2C7XL3BrQqecBNatelL7lTlxXFTzOWozRXTJltCZTpBpZAG4U1nWAUEK8GrsyOt
xgYaUQjz2AovDk51jNoLimt+O4mzd0Qe1kGWvQbufMO5rsCs4JGm1K45lCkzEHGeg9ehoqIn0SuO
lPQMI5psWqNQqTuHZBYVaCte/KIgspfr74vQzdirM1tgHWuE2q5+6tPowD3ycVZTJmHuECUk4nvj
X2NOxu5laYQmt7d7FFQyrVP+7nZZvRE/j9RRk/WfFzB/TiWUUP/KP7CJDa83+S8H6Edm5L3bY20w
4WBnP62ss5zbLMIi+J8/NSX5GA1CxNOl/4uJNkgroPcjuaoBagakQjM4ZW1f2lPcs3q1OI/5EMsi
fnbEbFzkGRpgCMNMK+1pczNAlziRyNB/KVVxi7+YR9v3Xnt4Dliddu3ft+z9eScECAHC6pPSr6mD
MYLt3tZNi3sxHxg6wB/Eagq9L1KduCwdsKh5yDwu9HFfgY/GSvxxXWHaUnjguI6t+HmV7FMS4dBn
Fn68r2fyUYUSwFOwp3b/erD358EZgPTnBtEptap3dQ4tLtcvZXUb9q3g5BYS8jfrRd5BNBujTyMO
JHK8fszJDYqbLvj3TZIOlCw39ei/WIKZpQkE+WOpSbcaWcOOC3a4QjYuH8/UFSqLNfg0lEg9HTyp
9WlGzBXZR106HIttB4nlVR6G/BKL6okJfx6Hgjl4TEXdInrw5WD0xs+fpuOMMp1aHmDTmXSdmMF3
gWfL6ArYDoilrXQIPw08wUBkpuy8QXHb26ncMwwH3OsuPtanott8/FYQMWgi7LBcmRJHCNobrqG9
lGcDiwzz8wS3+Lo40SGC2Pva15Cfn566x79VqTw4PQnE+Nsl9WyPzQEjv9IUzhW7NOArjPHsMMTa
MXOm0z90k5XDJgweBzZUXbY9jvC63e8VJnw5nt5jGeg6QAU0KF7z59d6pXjIsrVdAH3PX2OIvqIc
a7yy0zgYqepcQL8DJA2wTKJaPd0tFHM6BDqqmN4qUw7nhO/j793Ey8GsIih5iwZT0hMEELsFd8Ul
ygy6HzdkyP3nXsdA6aulvz2WDh5LSraBqX7Cs/BIg6jJPzLmLzLPdUYuXsCItDfHTn/YwIU5EBMl
4OeC8dXiHQ+jTsaskbAN/PW5YvnpV2WyxQZ1Y82GE89swopNRkKvy67Mdyj5RNVE0AynqeNqygzR
0a3yAkfckWQgY/jWuFsaUbuEljM2kCwP4sMcc9gCRyDOjSMkvyBR3ozfChupNaAKVkVCJt7V+dPL
VN0sRnGGypftORyUbu9Oy/t6x8jup1yseZsc4WNqtzluoTMmo7cZtHYwmaGqSLJeWDYdl2aXryOt
0d8Q3oJHLphyG40/9ZsfC+SGIqsBYgC+Wz6hWFNgRCCLbXCqyqFIWHAdrNpHkpqSm16N3eozrVSa
PmExFhQlXlWLBCy54/Qfqhkg/cWMoGN81C9TjXkCPLsM6Eg7ENzEXh9aMfdJVFzWQEw6lRmnYuJU
ld9POX2FKExKcW9Wy1hEAcpe7HwYzIOzEr17xXUY1dtG8yA/8YMa1QZBDrivExTIlaUGFyHSsMAb
hHJTyJ8m8LB7PosDcfoVpSavRz24vllDq4e/+cTFZey8DErhR/prUHy4DjOxlwYlLtnvM0lH0RwP
V1qcM07QCd6A+kxpNGMKgkLcMh+UHAbYhsht1O1J27TnPyuhn2NfubBeV7JZnkZLOZydwPfD1nTD
JqUvOJnzjnp3N7AYXa2NFk9xHf3PqEhRgGv6/iCs2578SSRUPeCzEEk31Cv52fYQGiS3MD5H9Oth
J2zmIC3XIcXfTFe7Bsynvytd17XwfS2errgVIooUOPotkPteAl+B4DScC78IJBSjmKlofzrxe1Z3
XSUwcwT3uDe9EMlZyZPe5xnXSMZzU6D1uHj1QXbGl+RMiGw4UokTefZwkiYtEerotuE7xxPwIS3i
Gop8Bri/J452oNEHwsWPvXkUNxx6G8SsGzLKqVB9mhYLwmEC2sDzv36rEsIXZ+cPSPg94Q4E7kWY
CnDSA1uoqxsjpWq4MoGBi+vXYa7MW5EPWW7MisKVR3wq+dx5JFhMHRUdGrwzSAQRbKPu5NtMZJYo
OoFf6gX3qSrIgltpkukvob7VuMQFfwXypdBKHvfu0nVpKCupIC1STM4gLgjcN6IyV/gO83sNPTfU
4+RVl+S29SKJ9zUngrS+DBt4e1c21OB8obloSbcICnArPt5ny7+EVlsq+ulhO2m81bxjhdQceV5c
4MzfNEIXSL3kLjaJu69qFM6kZJ2YM6Tx1z1v3bmbVpsU4XpqRFV0pe5yNH8ik3c0NoLz5Ku8nfBT
BLK56zD44fmGP2rFYTdqqFFgBCWk0A2DoifDNPzwOyej172BuT1h0pbuALQCAvH0EPMwjwFbI1AR
Lt0IoSmAjdJV2fbCh92lyZlFCpWe7uaAAdWEYvk/CSBHh6cuDes3zqliWJBPuya7Z13I9u4aof5a
Ay5rCgiDG0l+P//pjGFL/oSyDK+4QacTTf3SdOLgE/Ogq/uwJ4oP5ApExQQtawILFUeYHTVYVKoy
C4iSs2TZwbgc9fgZ/jzx6wlZTkwRjsAWuJHsAYXrPoRFOEoi63zZsLhzHz0ug8XDyDOTDcmJ0w86
1nB68XcyhzV10CLogKGlz0K47xnqGCRDfYv2dH7D3p5qaeCYxHmVhz/pMEhXyB1YlCCVU6pTQlIv
2cXImdICuw4EJUUjK6q83ivI1U3Ypnx6QJe48WwnlcIwslerMlUNNceG8b0KFV6EvH+FrScnLkdb
PFe5YGxnX3G2QkMwFHkt3cTmEXvPmgY3x8OGKRg7XEggx8rfBkOkA6Xv7bKxSdxQt+cg131mEqcY
V5HV66godM295YNDXgy6FcIAcRl+7sh2nJk23w0fraAvxjZ+wduGC7AlfvsAuGFXBrVc1hCkS8ff
uC0A+Cjp2uJwN+n8tSUWhK8l+/Q/lKn1w3+3xzcPQVAbLjmzkizJcfEKXNrMHz4VvrCOATCZX7p1
v6bvezoivrNfxuZ/dDIrIwZ/yPtBnv+gkE2QT+6YwQuRQjb8oBAqzE2C7P4jaUEVMbFVzhwxA9ID
aOkVTZLo5oUtWPhysc7PlLJKWrG4brRBb8YM/v1g2Smge0Eq4L/kL6ZIRDb5+PvfKAKV4sxidMGr
5KUk26dsgAeF5/Y5p926AMFRF8kDXVZl41bBMxD8xzLexYt0hl+opt3/DjEjzZpmXU7GwP2qYXOS
yKl59HPg2U7Afesk6kl3AXnOX2UxTpV43FRA8/tLFTB59XcBU3Fn3QVa78JwyWH3LtQ0zObJ6M7d
6I9lxy7S/ASxf3hrii3MZ8fW/MMv0jFAEgVy3T9QUmbPG/Yl7weGwJq/Mr9UcLYB5dLPZBtql9EI
P/zMDn7VDtfosNrb20rFeuh48EKL4gdo2wDnFl20/6Wm/vsUR+SDwEdclmWAOjij/j0rPRialbOg
hvKIWLjJRBe+yePZxmmASKAVruIv8W9qP+izRJflOzYpt0U1TiFrJ/TFQQlo7rm6lc5KtgfBUdLN
O7j1k1w0xDLTs4CntlNPko8rAzleBvZihA7BqH4G9kgbWc4Gxz/OIIFKG19hCHChucCO+4QNgLtf
UP3TUJ3T8PrUZCrZ5TBwAsx+N+kPtcpjbtQVef2DpCt6AXUTRg2789HjXn1Dc+PTwed2zZ0p1INs
ocXWKcC+qP+C8l0zKz1JJING4DSLX79r88j1KBbxwZN+Vsz+gFF1y+7FL0iSNoLsByfN8d6AGzWo
9LhqgOMTmtsW6yNEbxaa9oPOraHZoORNtq+oEutcYb2bWCgmxICht6f7OCeLSXxqLC6O9pfXkRCp
0xjIMeN9kRornc/sxz5MmD486XH+yARyEXFP8da1+/DfqCY4YQM1s9jigc51dKzLPFSZhkJHAOdD
I3ithvFn6hsB8D+pWCK0ouK+mDvxkEFMTCmuMBn6oKUTnyJIevRaV/C+/qp+QzIavyO8ppgCfFJL
a48VAjZgIgg8c9nI5e5lMJwc2qZeunwefVb+V7h96BnIi0P60D7tGsSzIwV5lm1a+dFP0p8Ex1JH
uLlSMK+EzNz2mkXU+cjb+VGCb7Z/h6rlsiXrYfaNvTtMer6jqnnC/QfQ5yyw8i84JyHVk2cTMCLt
j13GwZNKLuJ0PF57efkL+TKrLpA58cG758kROfQYCh4N8uNxKqwSt/Nf70SMGEd52VlvCNvYUO8l
oJKU5xSYADtxa9/KmfvEqe6Mz/FGhXSl1+4YXI75yriUMDoRTOAtD6xKJoEVW11danbAukTNrMYh
cPFHtWjGJ7VF71I6k7GvqIe5EQLbByFciCQATJA/KjcbxhwuP8+yw+LTz+k57tuWKr6tJi4quzgE
ejMUR9Uz0J0jYvCog2NZzn4pdoQysQ1me281n71t6xoWXfKr9Uyk9fymb1UeJfiuC6Kr7xcaAjQw
IDCKPu+wYRxBwVz9Ki/OkHHttofCZMFrch58r5kZVJjIi2bcTv/8EaO92Eds6oF/D4Hlmuex18Mi
RkLVq112pYASbW+v1Nv/QByXxoCzRXBBHy9oTpk5Fm2p/q9XbKDJnOYP33Y960/OSz1fQI0fd61C
r3kUubx6l/K4+XA+c1km+mRC/JFoxMCf4mWARMZUOOx5aIbDmbjTFA3PTiRVztAN8D87Eai/13jl
PHGmhxa6C7FjWB/8ZoEJZ/N1/eOXLLlQiePFKm+XKKbrRkX6+iolYwhdz7EufwLsOZYLcEaocKdi
OADPkNfypd2rNIlW+ZaUjlsNTZ6iDCwqQktBXQHndb2GkSIYMaeWyKv1mEJ5kHozDSad5dK3/3dy
OAg+haszr6Z+UOVF+EJNB45Km7qJ3gYSSYf+2EpJ+cxTncBehsaA51l8CLpjUJ6Fm3d4MTVPN5iY
FIEDWsHiUe5vbbTgoW6R3ulY26mzRAFwBaEGBGhxZ7hTWjcc7wzR+veL2fmGX7MRD24IM0pRvYzH
GRdUi17bBUB4QfR9yr6CTyAWC/vmFtiZdlMbiZIUQpUNzalCD1H5uLIUs9f/G/5KUPTX9ICB+jx1
J1E7riVioGn2XQWI6l9wyKEHQSzHwNgnSmpgNGLnQ4zek/JPBKxAINpvb7NhsK4Yp5XB2d6OKi6e
UqTiE3NaON+jX73pTzbgUVRhe0nTEgJz32TLdvfGumciEKGiTxBAnEucBnKvGoUM/hBPz35X6hbu
rCXtkIjPAA09EIS1MGFBeWReiw5TmpbvpI/IbvN6GTvj4WppaLdHVEUTa3S5/ir+4FMGnxveLSYg
3+WA6/KEJnZCNMTrcr+doQ1Aw/BeFp0qv1HYIl8/SpDGsOUeh07XccrJjGL5f1bWPNhiAx4KeBy7
8cZOt5an8bsELmN+MuvBJqIeOCCIqOXX2zTMUyzKQ7Kb2igBul/NkjWQnJCSUvwVFFmZarc3X84u
h/ux21s0RGc+/W4dFcqlfgeu5cMe+1nYEedJOV4hhElUXAjgtyL8YAgZN6uS/yDhHHCOL/MUyqcu
SMpfddXQMIXd4hnjMuWVKzH3RPuLH69frGBiSAc5BWRuggtnB3y4bp4M5OW04VFl1usAb/Y5vTSf
br+sGytyB5AsL247Fc+DEjvdncWYh0GM4Hzc8k8GcF5uAEad4oz6HQrweQd0F6cJ9/+TQwTUOz8s
PFVGiEg7TUfPrMjzxeddrwIw7CAFGnqisSvvHTF/3ogGtg8AoFbjCiRk11x1VWRue73WYsWSTqjW
OiII1vdX7Q7TPvcyyU8EEGhLgWkX6sl+zdjBzp/veDKF1Afp+WweZrZeHd2BFEet+9ZwZIVpqI91
ClEqMVAtFS6zmKW00L4gt9mbnMUH+1z4oUkXPmCayBOPXoK9I7KVZ2uavrHsQ5KWn55dfGphbzmm
2tEjKNpKfsCIbzEklh8JD2xYICvdFX22+SzTFAosdtEbCD3aifSCT5tV3jJhlYBl76ceRbDVn0jU
74UTJdVe6piNINomEnlUB6wjh4p6TDk24FeklSSWm4V3zNqjZsu5yxaGgUCRhM+auBNcudjPy5El
3zxbPk8j+nsmAb8rRcHu+A4VSyjKnRFIBmWcjEcwNHkk0emkofPDSN1hmrdJ1ZN86vx9exI7jYYu
Y5Kjfx9wAZ93cXVHqT3j+6xToKf7y9D3yRTN0XvWIRWOTKXvxnVejy1/lb93cLVLZM2B8U2HCLvI
4hl+o2uu26GJEevVtPJBxeIZ+QCVBbtGNaRWmWb0nbgEYhqYG88ZRCBmFoSOJDGVRpPGb1WH12b0
V1trKygDAZHiap5582vrphvnZszYIZ8Ro2iuNm+opzLKECa9kcnl+ZaMNcIrHeLhaiELdyL+cImA
JFJrORfF3apYCyJn7sWy4jt8HZiCqC9/x6bi8uuYjkEvVbr8zfsoNg/fb6i4MIQHRmRNBImTT2cB
sX2ShAZMNs+oahaX0/hvea/e6NH77+o7A4wRrR6lTkC7iorYCM9TOC2t4tR40rkews/DYaSWZXeZ
Sv6naHQ17lDLvrop0nWCcWneQb0JqmoYaLBtfdMZzhLk/LMtviaXeKESA8LmoBv5BMbUxkD40JBR
spp8gxue8EJHYnEIw0I1CSGDpOcsikWDQqa5XLygH0/DcjmGUCJtUyIc6BMid/V5t7STUJ4o+gyS
mcU2xMb5UkdLE9kfccOGChtoU11w3aQ6QX+rMEuO1fQLRwu7oha6PX04dfck/ffa54qd3LRYSUVY
WFDG+D6rqzwMS1j37vm1sFe5QQ8nngCsmG22aUZ3CbralImvcouONnPxWyZ9vuTNZh0SHv0rhjcJ
XxAcJUq//DKOjZ6xUKsotbBRMZR7qgdX7g9roS7ZO1/e2wnX/25O/fkD8a2+p3wL8jcyGX+9GUy1
JIpi6GHEqu7V+J7q5k6FR7iOBp4jMNsNf338MGkeDpHxH8Ld0brdWgGNI2Cuq91DNdPNO9LZgUzN
8fu9Y7uHBBsJyaZ7oBxhU7slDepZmz8GT++C0wlGZZod8RnR2ljjkoaXXFmu99IDhrg1KN13iJSb
MnnIn34fJntIP6Ol1vgKAnnu6gYjnKB3CHWtK3wg2kU8/DWxQQHcfPRDQglAzBrTl/rFoagz0/im
lh9a59IF2OPV7nRRcasp5eLveRtKlgGMEjQr9SN0lKHyAaF1xQl9MDUWYlJ5ACtcG6EaLT4UN4tz
UuygfJorWGeEenXMCilpFJCsCuTVIzNsLmFkd7d1ImhAdzirDsayZoQnpmNjywc1mXMaOLkVU/n7
gi+5gqpB80N4G/VyY/MA8BTMxkIu08daK49g7Dxfbt2DUvJXatmAsxFrjoqFKjPUY8cEcQ/Io4jD
mzRcgSAv53HQVyJFiswoqG5/9Erkr7KSeRnvWLU1d677QNlRSkaUMnthJauuK71Kfavr8xCqeUk5
Ozpc1y0o0Ke/vR5voCssCYQkYZlme9icU49rmQA1UWCfhiyZDawISnkbsDdeJVz6jjxKe7jxvSkn
iIyJkzzjH2cW9KnslqrAd5HxYThYoysmBbSnJS7iVHDXOXo4/9eNvztei9WMmhMosB7j2e6jIe7i
u6VZl2xUP4y/XUxRhB0bAAD/vEIjI0Wms5mL3dgN9RC5tsxDAUtToj8vfiAi0/dbIdmaXrsvrw5H
HxfoLD/HoP/I1ptvYx7WEQxTqRO4CypijGNYXaGiCgaUnu/kwNjDLYmhsoGf8G0ONRWWyc2hhQ7N
KJ2wERe+oY+7MPCcHQuf7w3ncmKyh6zMNfR+cOMYV+dWx50AT1gjxfPBTXlYjr7qBiEBvrA8Hrn6
5/VUFO9gifDHIJd/4ivj7JW/mGmDjx/kLA2cWUtgtdbqPS2HJDPq5xs0OphJMJ0CYvUsVJHjHscZ
6VZGeUyThjRIsNSQYmQk6ZbGqr+KFMEQgGmScXjXQoEcYrx0826/wp+8theIL+ZlvqgsZK2na62S
/12QJzFRU+gTzeATxlIEKxnMBuYN+mQptkXA2zxzQCVV/zOZxnLvZcneL8B/Muj8Tc57NbOA2pd1
Mg9JcCq7pez0hS7/QU7ro/AsBGDlOQk0wDiPPLC3fNT+UPnLg/6DPUotQRhUU2+LRgLel9zol4Tp
11DOEfSc35qP8r9zXkPyi4t1kP7WkaSue5iuXNWLKkFxJJPic2+0DLuYkvkMalTmp5apnBWFFNEE
4XqDHlS7tJmHGTvB23Ryw6oWLEGD6U/986mfYESVjy3HReSQvwmFLpuoZ5m6bRXjwo7WHDjyCdvY
SV0KTuz5YGVuCZ/iBOKaaaMMg99z/CFrlnCWv5g3jejPn1/wT2kh1JK+RKGUSicas0Wmft2p0LmY
3YVJD413NMzAj2ErMKXKkjREgxKZjTaewXYDlLxR9Dd5T4FX0o/lW7JQpHaCfvMMOc/4fLz5Ia7p
EbSd04D8GCioN7pKuXKVzh5qe5znB5rZc/b427EGrwwjgODKIv3lkoeOoxXrJ4pRPDIMsPGnYuFB
/HRYC+bNuq4qs3SzJiKgQkkuKhhtKdo+27YRLI2X6U2Db6Np95Em9AJDOtB6hFWqG8icEHXSgYOV
TVjZvpWVmYQiebM5ye5s3Xm8wdlfBEGkvVvrHzMEgux2AJSR0vhqeIHO7paRsrUww6In8I2EyLEy
5w5iJ+Yl8IY7FfskXjc6NTnQTVerIzs+arwZfDJKVeFpmMurwcSrzPuy6AAWXDT1qm6dRm2aprLQ
NXNN29DlZB2gxD7Qg0jP/oNX6GAMiG6kFX4rNbITVxjlBRh5HjrPHez69rH/z6rGjyL0CTNfiXUr
jLzGLwki2522o5halteMbec192ft0ah2Wg9Fh053g7e2x1fVK7icqq8hF46KrsjzCDlXImLzgTzQ
VE9tRr3q4hnnwMU59v8I1kNcoeC7+1mvJySXEsejicbS5KcLOMPgsiJ8o2U66xcecovSkr0MT80I
o+Kr/3AUfq7hKQapWbPpMBu+tHXh3MA35fd8iNPurwWJtHP6xYBPjbxfsZDLPPgEx+SohSpYchNE
C3xO7JoZKSwau4cWC2jCNNnk3syAJ7KZ1KU8fx5rA8cBnVm/WxpiIDz7KAltYYPfgaU/2VnBdpiI
zn17Se/ERBztwoPAjn2lRMiFpeIT8HqhfUJp1XcbqyWzWCSkn901mp07hZOHF37odqXqA9autkTK
HbayJrsDe2Ih+o7PC88wxX39CDZdlhqzz6vZLJdRPlZg1JVpPfnJ1WoqzUq5e6Q5+t2wJLP6tsDy
qjEiYFqCpDjxTYJhLM4fKw2X1bs8dMXqW5FUPb5ngJIt3xY67+Pvcd2kh2JLY2kcFXDFZIVHqbwc
j/zA9TrPlamUXWIGiHC5x4HiOrtZ/RVFpUZRM/H791HTxgEFgd3bvPyj6Oa6qh7+nh907JCSZP2A
VCkLSyN2kMND81pqfS4aLWTQ8EvdDATPUwlRUxhGTWTCxpi0BZ4gy8ZK+xFZKbTzduF/3sTNytay
Y/sVh5q53NiPwoYrSgvTM9wR3hHLCYjTOyB9vD03wO9+/+hU6tAAcfZy9qFqYMaOsxeFjhM3JZxf
UxdF6yXetZOdoVEGriZEVFI/wM4mKqU1tLrpDFebjuEG8eEXToDtU3OLFL/dqqAUzBX8dfKBD14e
AROIzin146dRjDCPdDIWpXSepjI/xy9jgx9Hgr4hZYlAcm1Ol5HXH/uSEuicg+X5Gr2PE87mYUkB
RSfmT8zU6OnHvFlqiwa9bVS0EDaoib6B14Ze/ONJFtRyIsAs+iyn3/ouyKsJKccFkf1YXHwCkLe4
f9j2UxlkLW/kys+eWJiSP4RB1i+bl/qJ1+IsAIwTQ3+pPw28v7NOqPxbp12esU7MwX8MSD8Fra+k
/8zBQZ2GUdau39P7jgMNLFPHBQjGt2FQLzisFcIApPDcH9JoridoYEjHJb7V9J5MmuDc5VGp3F6I
If0U5ObuOGcQSrkTKTxo6bXk7ca6Tsy1PWA06NiBujVhDO9tjNO1ff+fqBP/7Uu4hzwOfdJrLVQr
j7LZx2q+lbcgz+4r28sHz3OTahBdY+vh+duWD2cItbBuIqmTHrImoCsO2jaC6SpNVtjK4R5lR3Gr
r67I16nDzghG5qbkDgGHobFBfsX201lzxxVGQOOvbzetcUM+5slgUSckZGlk5wsCsI18DPELP+F9
zsMFEblhBehs+P9Lg6LTl/VjSP8Ryb43Wq5wDtTY5HJVMYD3ju69RY09CHb3HG71qQtF76/7/0y8
A4T6cA32/DDLX556y7B/BCOXapke+4vFhiGu2Ma5g+wIfxlBgHQkxQ5PTSCdJSEDkIaMMehw7WUt
JEeItupoG9UBqjstnMXRJd5PM4yPP3qQx63kZDNuHoZHV/kNsnoVvhv2td00Jxnx9qMu1F1eJDl4
c4MNr8pmlJISu4l7c9lZfdkSpA88o1lCxtuLUDPpU34i90ByiUqzAtJ8IWHHdut5n4smE4yR92Tc
KRS/6SMfN4LVUBk4Q8G8uJFN9vTC24UCrg4NmpZwxiRjFVYN+lIzLqG5rqE5WJzEXUJLsQfeRAlg
L63E7FW1jYVXQCz9QMbzyKhTy5YWKCqA41EEofbzPnD2/Z24DI0vAJvawrhc9LL38yV8/rDIZwMu
kDhNToou0S5g2nKWi1WA6fnxjw4qkJynmk7UmpgzlR7pCsgpaBDQMhjR6nQQ12E5nwkgE3bpoKE5
30HP7VWAi5sZhj2diSM0hfvkk+URynHkzUv34H4Un7CHn6Yy4Jzf1rPg4BvP+W8+W4DIj1aRShjL
46fRDVP2UB1mNs2cyTVhnyc04QP3MKmeXxzcudwEJyOt8qUR9Bes1M1lM70CpKyBPY4ayZlTRYaj
HsSSbqZ1ooPXRl2iXBZ7K9UOxaZC9WfJaxf6DYJ5e68HZ5/3AsSwmWbrEffr66UBGbrLHeM8I8/P
NGYvYp7CbG0SN3gmS0cu39bm+PVl8ClESKSxhIrBDpVxkRKGhwwSSQ2bepA3b88OK290q13UZNn8
bRrhpi11vLEhXX5NxghzpMrmJ6qW39fH8AxESNiV11S573BEVC10kebc5nuJ0WKGmpECjZWs+lFA
kVBz9OFIMP219SpzuA+7i5/wkCzxERtfSXEAIW64wg9WgxAFWXkuyLj83KoZoiuEx4G0DUSxusa2
s4Fb0QrXIlKm6/wwkXmBkWhh0iXqRb0n2J035LQhnN9Sk9OGY6lFaFYszMdRTXp5dMQ0gRp+5Qdd
emLe3a5mlqtCUxBXkNemi5T6OY3q3+wOAqiyG40y6kZu/1BH/YPjW3IaVIfEt7M2LJM+8T1ZLY7D
rYy74niEfvJZrqR819PONAPZEoknhXDCVsz2YxJ7d0oAA1h9o3sPqrPOYawi8kF039OLfHzu4td8
sM4yA1VnBnLKhKSLHNXVTjh0ZUkoQT8fIGmX6BxWLXizSa/i8Q2clJ/bBnhIZeRL/gIfrOHSiln2
8Na4TjVQtOxhd2fs58LJWM+u53b4BclXEObPQxin0ew9L1STQXqZXOhFaBQ2U3z46mTnZ/jyAo5W
4DtOapLoknI2uPunXJhdHcBpcgL+dd2n62yPHuL0fjRuw/fjzNPuhdRvc3Hjm9j/kQ+2For5MMyu
/zAAwA4WkAqHKIDMUEyyXys1TyKtU/QDNukTaOUkbl1l9F0Wre9zjWIeBIMeOoXvw7K6+HLI2gDf
Y3IGQf7Ra9j2yTvL71BsVP6wBFQvXWP9+g+0kFap2t4qR41S9mVlFM1Fe7pEYcpqkCwnnlbh736W
j92iymdW5WMBmeIZvQPZWXhl4MGdl9Rk4/NxlrfuSepXYZDJl1VYpdA4Erga13u/jiNSw1NHNTew
WSJJem4uccpqqeHFXK3TYdyvzpqOJtu5WPnigdWfm9MWy9IorRNRI6frLiaKgJptxD4WRdOxu4e/
UOwts+qJ50+wiMlWH0sVH6oeFR66HnGVbuYLSnfemjeMshJ2anJvRPQmB5IKsYCe7nwu9oR3fG/p
SYENRZOZsSQw09L710YHjY+dsF+w3nxmNn16ns8se5ehl50/+q36zUO3rQomE61dlbAcsprf1o/7
1xeWvoaGHAz54WxsL4biKn1GfENVE9vVjFjyyYOV7cH+QIfKQSAcP7kMfmx2b1Cg+Z9EfNAE4EZ3
NdbtxGpztEcgQgAOTHc7RZfgBkHJRi2FjIaBSN2KQnDMLWHhTIDOe0/A5wWm/zzB49BO1k+0qriy
e75UFm54Ig7IHyH9DkvgHO/tpdIROQ+kEgO3wuY6aVzCtWqDHcw7jiJvrKV0OpNhJlCsjFqsSPz3
Wu2i+b1wHtCuTkjhPxK5CdYF/TigvsfLyOGrkLWDCoww+h/JbrC/H8uFZBFNMJErHRXJzGm2TjFx
hvaBD/DEHY+6geMjP4jTPTHRFf2fGUJpxLmqq8DdAhK4fhbu2Ed/OuvQFqBbkg+ZZXoPpA7gG9vy
YhL9ceScYXIEQVL1H8syqDdD79RbBELDHJTJm6BTU4laM0BPYptf1nYTRbmDaxkSHQUFa+flR2cj
vqmpLGbeugWTCuUTs8BTr2xMTKSEDkpot35Cm13lL2IK5PPe8JGlSVV7A2LFgtjgnNKyZ+Wu/mwe
IRWzFFAXDXt9Bb7ZHP8OIE2hlq0dyFLsucAJwOTUobsaiLpqk4U+Qbky9SFg3vW0Vzy635ERpJcs
I+wbdhVr82OMi7vgp9fBOmm/JPMV+YtebWbQAn/8l5/lTIWNeKnmsxNhiT981HC/EsV9OLkyixo2
O16K/ThaP9xMLdNcu4BVTA5dlwj9TLrAaV37f0oNWYJMzI/Gl70zJd24kHoSHNJfZ8jVukPW8OJC
5soXIM9TLu3cH6fHfBsEF5C/3+WjlOoxpB5Ig1zHHMt6v1iIXgiuOMHnqlGENFp7ACTprPeP6akX
9SM0MVFarLSQi73E1UxUSWxjK47yGgkSdPFUK/jpfM0MoZsRLe5xDyV4oPwzL+IGCGL8pJ8TTyfr
tQbhM8GmbZFupUx35TltwLciFmwxg/NP5nriOe8atdok5tpAUtFTdsQlSG+ueXb7EVeP40cRo6FZ
FnuDuE7WcKCMe21owEVCuwz2ocjTmj11KypvEHvL9i1qqNFrvQcQ767fZj6AyxHQmLP2nroniaFK
hSFgFB0cmorPkJhob/oEZ3+X2BJ4R0nJU9Qmae879aBV7Q2g+6u8bMv/4FHHn66EmUJMVwwOWYsZ
vvP8AgrT6GZdLA8d3zo9+2AOt0vinew+q7XYbuyzPm3OJoJkxRHw5/kQdZeKJJ6hjmwjTwqWBp4f
CF/g98gqhywyLikG/ZqDF7bW16a0hE6fN+3V6Qqz6HzjEXlW0ePztmBcXwRCSx+XSgRIPV20LTec
Papkski8X6TKazGL9u/qEo2DG3xcl1ohJWv4YBhZEjEz/C6rejdAxjuHgXSv8B75S8CmiePO7Rdq
z2Rcd248SjXjMDvSzL9CiEyaeW/vyFuPkUYznQu/Apx+Ie7Y0JsypaQ1bqxD5BceI+ezN7qZXRaR
6oY1O0/2+tC+GOgPdkePmyIbhqfw9QmnutiXUIaIXiqW1dBpupjYZWxuOYt/QdhhOuru8ABNvJpd
3YtOBha7Wfcza6roNUOZXrsKr8JuKoBTTPUutWB7azBA4Pc5bXpcTg+VyYLsSWRT3sI8M845ym8B
ScYSS4lyTv1d0RzEwF1evUQdDFYNTXldxkA+A085zI/GcFfm/Hd2TtppOvyXkhszYJDusdsyUQ/K
b5Qn3zCoIniEChLnX/+k0i+AMbK1hih3Gx8lATnqw2R7hcS/sOdHfPxuF/4hxkx5I/CtpDrEY/+h
pWEbxWV+hUecriUPohOCJUPxH+cdsFRIHYsBI0yCV6BZzaAnVdsrstSoAV7VU0W0CNEdiFX8O5dJ
hq0SSian222lGOo4Hc4o9ko+QNWd4BALXB7GY8X7rwYxc2NpHI65vVV8eH9rKhfvJs1nry2vaAjR
aZ6bCgX9GM72MoiVHdkKbHNeGUBiPEI5cGj/kva3hbJRQpHLx2C9MawhPivQczmNlmpSZYBXpGHh
Zfatzw+ZVpNMritB9oqwl1HPbDW96Kxu+nNwLqhavRoFgiI2zPWltwKgRP4lzobcHEmvTe/tPnVK
y+l2er0RDuelyZ3c43IFG/8VdL+tNrtfYT6s0PKEAKEYGa/QOpyqy6Y1J6VL/6ND2K8601H54MlE
N07qPku6kjTt52GIPhCfbkjPcrx5AT3T2//lMy54X3JR95xIGoLxYt265otQZposXIeIcwl2G+5P
D1/0CP5dhs+Wz8L8USAlQQTMCJSTn36T4ajeL4FuDXVuZ91B3UdS0xYlU/tyoviM/koopM2yRyYJ
E1WJKofUhH70Exx4qi4aUQOmfkajZhAzQRiHMfbN7GVMU4ohoXMSP0YwT1juxhhUa6k8NtH29Fft
MD2LlQmPUz9lczNF/I9/SDdos/H023911bk1WihqGzFy9vN4SpbhTf+NZO59gfJQd0Fz0WxXwvVq
Vn6vL9HS/hHdXM4cFvTb5erLsaQmvx7VqeQxdtJbOU6Cm2ICdMwF2NYjVZfvoZk7pQiquWQb2gN7
Q5qKnWC9vTF2Mop+ixpNfdudo7oj2/iQ0ehKaBFNH+IWi5o2q9xmuwjicRVEotgbVKkBZAekFm7g
BvCSEqjhOmts7bSG9PNuPMqnB2+j8kt5WV0cjQ+1fBy/aHcists3l1gfeKRmaQP1ZQRrEjaoT0fd
upBpXFVmAXvRx2wEUg1e3yBlnTdnXwlN0sM3I4epF0cXlSKS227EscyYhVCTRXX6PAfsqw/6fk20
mfpS58VcnziF/Xky7fG472Ac69dE0kUPpjCUj+PSMJ3u9emTpdKdVdsmDxEMvyGqHjWLsHET5Rqd
9RlsQHIsPedrsp5F0XxKjXbYrnW7uknXVqO/jjFbvR0Dq0v1e+BkSC6Wv4t4hK+D9ninCwjsNWKM
gzZnzF0vGwRAVtx0ml77gP3O2VG+VAb3s4WYzDM+7qtz15P6h27mh26tm9Wujk9y411ml2V+v81h
08vf0qNMdlQt3H6JCzyMlRcjzRoxiP9LYG0mwvAHV1wNU+CzOtbX+ZSUIsXpS1VZrJL9yjAang2n
yZoQkIvGkWAZROw4hmnY8R17Q8I7o3CsmxC/A2UQEkczFlMfB/FgEwQFNjij3O0PqqylI7+cG+hg
crELqaEORKsTB++RMtRX4h/nANyZikCGngc0fbEJbKt1n0tFDrZLSxyRlU9SmyLzfpgmYKm32Qhk
6v7Pg1qNCWDKwYfIm7ZWlrWTV6Mo/5Sh6soMLfPBCfQYkw9+uljPGEXF43gBSxuPh98qTxfrfM9N
+tB10aXtF531YvNNLuyJL0k+hd/qwcrJn2P32G20aKLriWUiqGALeNdzGwsMeh9QS39O+0hua3zI
otbsDXfj2ru4BflzWPDHEcQRwn+vr2iWn/IjGXLgUP09Tu8wjZAmLVrWq7dIXFv10U1e//uoicMb
wCJedUfpm9EO7RxcgwZ6jJWRYzA41jaOFUvqkKP4EU8xOVRnOvKKRuRxZ7n2k+uDmlRGlktyMt+v
quKRkPia3VBhw2veOBiNlpBeSBipZK5VGsWQ/C6Mk3KpA91T6nBYBvh6OYP7WgGqfpX9LYqeABeT
RZs99TRTYusTd+/bQ5g8H26hNtXBvf2yMw0cGErgM/oKvGIcRSH5x805tekeqInPKK0JkRz3EdXM
qsJXxR9zrSIzywC1NN/c+BZ62E1LzZzdMwxU+iDH4ClL0nWulUrA4+r4uOMEfC6lPamF4w4+r0ku
0Wq84UojkcyJWRmTn5H3wUf0zUTwWTR+Mp1yFnJuJ5twjiJw/VgSvHMmrZOwajAbRF/QlKElk6kB
fEDXSw/GsKDsn+CDl0pnp1yrLgDNcbOFr2cmWl71AcgN2FwZOZ7rTOTwR3bLldRm2Vz5KM8U5vVj
RP+ucIDY16iX4ypct873V3udzLscyqvokgBoWLsSfGrcMh6OlrVeOTfRbcN0Ygd8soCZdXHotVla
SOyo8LkfS/pRZyWaaLQp9V4/w4MNZMvU2rzTXcbAbnTa5G5sRifBQumgZrsTDabtbabSHU/+a25g
fQwSnwg8ozn6ygC9CWS9fGV375Hu6lTZeN0ZzUSLQFp0p4tZbVWM+A4lyGc7U6DNsK9wI11w8lBm
Xb/Nn5glSIkw/fl5hXhuL/BhknR3oPf/0KjbcL0edxC5t1P3timxOjjI7M58BeVrWVIuQeQQw6D5
e1AjkcO1FA2hW2Rdw7siHPemiE8Tkc21AvTfA7abkCPEBTxhl/4i85TF4JON2P5GzY1N7Ngj+GtE
FiRdX3Ta+8hQsd/iMJVvECNw0R6EFAGijH03dGRRCeHlxRt16wmdID5//rlonGywZJuiQxAY3zJT
dQJt87OqNa6vcdSoroqytkVYpIZDktoebIh67go+h84XnS4UguYdpfCtHnQcVqGjq9THw+JVX4Ln
4Plpv72xUXv3T91HZ3vOi7p8mNcBYpnKj12bpiTPgi3ahZ7T/31q5w6zLR2/ORrxd98OrLAaQDAU
573zFfdFbki9NQZX+6vTn0LCCG/bCmkd2dvQKGA688MINlhu3uQkBj84dDhCy7qCdwAwGgwKi5q4
SZuXNdux+UGVIrqMO7VwoeWSbPOQVezxEr3uMEchLAP/48ZQbEGVbsYgkH6caa4GFZtwyB18Z7Jy
meSfIVUPj8VfAcdAnYe438TwAOxDGWlCSp15VONnMg5lK4/0mLlktb3007GPuJy8te4nEBfBC/Ms
q2Yc/LiBJ8/mnObI+qd8a2ape3rlde59dZxgQjoHCysUjkGhD6ywNgQCo/maJ1+X9RqyKKZqe0BW
C61Y3cWAw8vtQDtuK9TP7mzyhRnmidwC4UuyBQjUw/Y5el8blAfNXtWo7YdWMYhRtf+HRieKJX5R
wjNjCLDKy6YaKt40Eqp5MAFwEOQU+KRUMvMfx1/4cJb/71iGgoSWHRd5KB0s0DiO2JXB34XATI2f
IVmCS3ftFyM9bsj3hIrMimwXlfVWbPZ2fT0IEfWNMJafq8VLGBAW2cfd0eTk2G0DFpVrj0ZoR9/1
t2BnLb2VWdOeGQxGpNiNMYZ3v4Uda5nS6D1oM5zRQTZy2Cgbpc1Wlx7lVKtZlYp1VKHDlHoRmCXV
aW6sogvgp4uKPZ352HUz0Cw/XYd9QD0O4Adp2A8jZjeyzxlcNsNeLWxPuil11eUl5tB1/bYdpuFa
gagLwkoNQL630Og+4VI6UTtGvvQa3G6I86M2MtdoheFCHH/nNpckuFYFFevn20NV8y+vHlc+RC3g
5UeZZ1ysuigYhR6AEEqThLXWJO7Tl5IX3xp/99AFMzKYLwUqfaDsOGV7P78eM62t2bWCCpSCCicX
l7L9s5WuUoXhjvRW2f2gNP8BqX6RWQutcs4Ne6SETO7K0NVtIe6vfHeYXpFd5mCVF6f4qdrektT+
9oH9zvkZ5hbpnyaggmAB2Gh+V6ww4vn75U4VIsZoFIeFMSj7/lgwRD4qKam4casjDh2blra9v/Wb
vKIdviKH2ZYFR66qq/k9ORUyi6nKxfBv/dw8JnaZAouLciJLbkY/fQtJ+GpFLtofoRU8gHL7C8nd
OMYUklPbJpuz7XyY+3RtRcqZYqtuOGw8/19ItfDuueUyrgTnZR5pbGQLlRew8LM8h/NFEtdqBqka
xJHMpng5s2ai96PkJ1z3nsgFRvF3Xaj1+2NupUZsegHxfGiaiRkSMVJlk0MnTa5D1rbyXywmZ/NV
Ca99hCia4UupeSKj+VQ/MM9WRl+7Lf449BWagYBVN46bk5bTGsk4+rZBbFxPF9zwY/VA6S2Ap+Q9
R/+6H+IbhxtUV4sVv9xpcWjQYLBR6x3f3UUHl4L/uhOGYu6/aDKqHusjIkVG+A2k+RjHr76wAkdF
IwdkiUcc0m0pDTc0DVfKjC+WB5is12y5oCTeDV86uA1wloHZ6euvyrjCNVmILOAQ6Wbp2WbUggh3
0B90vE9tkjlaJlGZc0F9texpjVc/WEtidwTRHAkkJD9d6VBWt3zfnUtqYfoozbHDKRuwUAwpy0uU
Lt6LfAh2T+1ZBQZzztk7e2AqHU20EQXhr3eCXQSpAxX0i0NjYiTky1vY2Iqn+GZHoMVfg5wyeXek
2S/2VMiKQHw3B1TdxFCffPfXK5tHTkMwjIyrvfd2zzGXi3xxgj3MCw/KWxMIA6qDAWIcoAGyRXjo
eDlIRVn6/GQOjxF9CvxHi0RXKKZhF3+b0pxbGC6A6azj+gJdNv57IdsVmSLlaoBpiFxg2W8AQcQL
a/2ySkvXiA8AP/wMJyKTgH65StyW1ahdMcUHhBobcfyGrleNXqkT7hAluiOR9JnvKvQuHg6gpgL7
eReRmZRJoWm9avAOMyHGqqJCH6i45xfdx7/GNdL75VYx6HW1DtAN3zocKVUOQRDpo7WPgIWbIApa
vNF35gb7E/kXpD7T5Vuuo15R37ZimBL9Sauhce//Z2r/fcagD+WsRQAZhm0kLszZFugxw3GQBLKo
if1nybeR5JwQMbhzAUKMjSIIo5gGEhrKSliSgqCJ0SJC0R7p3dWtpHOVkaHyMWZZ2NcRSuswzpem
U99p1/kbMJOvacvcJt3bw2NgwSvpCNBXGXKJN0/xaLAt9c4aHRLyZVZ+8yZHhEeYKXBWXp3Mfo23
8liyfZtxkR5GO1P6w1XN7V5/dhjV7f68fQMXAoOKI/0FkMoTn9O33xe5s9BtL4azVbSlwe/ufvm+
2OywM0IBS4eQE3asATjNIZhm72/xcMPgQvvtgV2SV5d7Zys3ZzENYZJ2FxmD/hN+NQweFwkZdfzX
r2IhsxogPqaXk19EdlEOzt9XyiFwEwHN2hldTeB/5VJFcOieaRJvGkU/uaLTqvSZIxh/lWcpGoZL
N8KaXN3gY++ouDeGeYux/F6jj2hcrhpkokVxB/Vi1BP5H+xfKrH1UC1R20g7uXbQdkz4QepTlibx
9gAvszBLTXyRsMTrCgrhcmlORFkeH5pGgRJQQmw4Do0KFPhRswNc22k2WpcDe9WH/8Te5ZLdtkID
opKLM0nNZAE567+eSJd6argbnYfxCPw1WoYF+s2pDFRdDbe3eotuVWlhGkdTXAM7jZOa866IKvO7
VXgCpmmU3kxbUpGYY+GC+2gMm9+HmXr9ObEsKXTwphchYAASfARQMwJ+fEaDEOos8r+C3+VlGpG/
6jEVp2vW0V0DbYgkDC+J3Ie/gO968xggpuFd+HR+emtfqCkGWHKRnyH4vG7sUeKas0S+hh3qw9s1
BG5c1DGqyo2+cDkqGsoFDwARWZisBK09/1NW8CeODlFLWYTsstQtSZAQjrvo9pihSw0TOqymEKRO
EZgSqUbxp/iklYb2sJNOLg4YAHKqdosgX3q9Sm7QhH8J/BCMSdrnFAPd+VCFC3pZTQwHUk00eWWh
HvQyAYdhAdamL20aGJwHwABZzKhT6ip1SYyJzNKrqk6BbGVt799UgsY5ucJEAe+ugmTNpNMCvqfz
naD3RV89TuV4ldIsOQhb/8jz0s/iXoytSHJjbSTlCCk7eQ/oUUPa6DW2S95bMdd2eWqpvrVcWihN
ruZaPloVUPZynwUAo3ryY5ER/ORkckLVZnpGpp9MtJP3jOPFsnNrcDczPa8QRFjeHsDOcQ5QQTWS
qDbO/wHErF+uihblM/eAP57Zq5waAZ6JHIdCQi/pimND+013t4XOw99Cmgoko0Xiw44j7gZCAvET
dfZGlk2PRUXK8pRZNlqjR+rM0iTjLaaEM8YP6cjJVGYBQw8iiUQB/UUn+Vs/1b0IJdw3pX6d09+h
PGgqY6wvGdmk3gJ9KHkJnbwVcQ+oV00ZXcYyzjPipOa5NlrIpZnrK5NkX6nt/ZGuZyVaGxO/vsJ/
jjOGpairi9LTkGFiW/qpEw93SlmAHv/6oDmN7NwWQlIsFg+0V+j7ED88rJOzNzUWuaejpX9ctbCE
ArkvNM0wrsbtIXCGL6vIJrOzDqL4t0qfA8s8elWcdReQZyLMXiMA6lDVVkeC6nhrejImaRitiyCc
hoonFVdAveLqYSVxo/NWlSrF0X9e9/A6H9ZP9j9nlSf/d6Hh/9z0EywlMKKm/vBRlAEXzKITTUXS
tuQzhnw0jlIFtYIL+C36UPl9bWCXvClYpD5pnUN9/ar3i7UQr1oyHdLkCeEWRjd3DmciiMfTMbcN
/89TQEHH80Rt243MNS7b6ZSvYGNcB95Dt9IpNzqX0WxCVuTj+J5ecuR7NYSUGOuTsudyNA+I7Sqi
IhpvNPNJx9mSnEqOnlMFGdH/CMZ7xu4jGr4WPWD1LJ7Vd8rLS+K3MF2Yj7lpnuutA3fo8biM4slH
rAHCH7I0J11FgrWyXKKySD/5ptSpw/UHT2o7L4YtSRSpwQ6XzXq7OqlEIl9FK5AijtD3g/KBHHQi
cAnK73vcQo5/wdizFJereDohUevkgfA/YdZZ/1OyrZjr6+uURC+Q5sYX1lMgXTQ5u6/wqPbQ+SXW
sEVR/sobLYUEMOQsBLLtRKqdpH17oROSsAPiqpmrB10D40D70WeUxMY++a7PptvxosTxK4hzDrVl
wfimMav8HvN6hbArW1jN7FYLodav/yKIYtt0TJMCn3A6xe56KBw+ZyHnd8pxxXu96PeUzcNMLIYX
lmQxwN6O1PMjfpz94JDnS7VBP7iECWExbj1VcPHBEHvKxT6TrnfGQQrUP8suGs5IWlJm6rgBppAx
2Jh8MIr7DQDkBpSVlIZUnOuoHQXNtsR9r2cNYdPRuJHSmSDssvxtgj3ZNip8lk2CkoRbnSrLpQE6
46GGOVApIqUK7IdPK6j0lbphOJSsG/i1kxLNl9YrIzXxRyof675qwoPDXTRuBgEdIkCzXD2MGYcY
Holi5NWw0fYe3RlhZ7DmtTItCWUotqeoS/aSRTxYU1OqqmPZn9zwAFwQOmYLHL2MxtbyeYDL2MYU
yb+66kZBDBvkc0vJ5w1OML59PA8CODMCQRf2C30vUVrnITyGlnLw1XVVDTb/qAfYI0pr6I670AUl
pb7MQdUASVmGxTHW2K0zZTYGb0K4QNqAaU95UHHVCBlUHFz5yuNMKQsVXGEOXa0Gb95EndGH7GXu
JeO54nwwqg8iT/5fTEL1ITRA4RkCDLFqwHicoCXspuCOjXttpu3+73cEarl75gF25Rg/A/iQWYnJ
alMBBKWFFYTnNZPTD+Rup9cr9LaOqgLyTejy+FCCxOIO62L5GX+kG3Nbp22M3gNXm2oiQ4fp/Q01
7T1fDhiZWjUS6JZYkHA4veErcYTHJD3jwdlM3qh0S4ud6XWSwvFPTHPzcxjnPYWS+kPHrJ4fUcKp
VMnNmUNJizybZzMufUuxoxdk0QDtLHGuNajChTVNn6Ajltfolv+zhzG/E2FYluREGDQiIFGT1D+R
iKlB9Vs5q4dggLpX+gUWa33c2aww08fcjaWYVkWIjbHTzO7ZN2L21uReqd4cF/HvGMY4HlJcsGej
8oTx+5xBqjaFEas3VLSMJYIsLRR/77l7HhvzKC4Jc/1JBNw7sc9hUX8mZJUFTXDtcMrX6OwMVSFj
PAJRMU8wKt202WplgGckZHUCBThS7NpUtk7gKofujKb15kAFoJsqhoWAO8UubLvUlExQ8SYNg8HQ
QZAZi5bdyi0kyzGS8qhsyMkVYZwsRAQi5tMjwsMN/BOxKo8geucCIUmvQqWk49F/wpo6oW9dCBuK
TlxpRN7kYjQbMkohnVCIqpt7vbP5jcJ6dFTNATN4K7AXQiMz/PewM7eh3vmuLY/RnFVNCg5HkPFT
pGnvQc6yd1p/vtdNn1Btx9dEWNZzODLj4heyL/L0lnnOoDcw2cwlLJZ3AgR/SFjfsAc714M0j0m8
YCp4Lg4mU8Wu3oUhgW4eUOEKoKxUEQu/CGjqfcpeg6FqhBusFH4kucNByypdxBZcCS/dXeqQnWQ9
HVkyQ4T7RlVONl38jDsR9plQKiLamcV1FnHbGEulsjX8esp/tQ03bQKKcduu0waxbeec+erDpVAI
yUaWZ4BSXpsu6rqS5pqRvy2wjLkb1xRx02jNp2hr1ebtU72uYOuaGgoq+BaHLz3XlKKf2PV9buZu
CuUlEEa7WlCCHpfct1KNh11W3Tvz0vzLHpABMaB0EWrHeTZ3VlDufSb7PPfdIX648P+5BUmHtuNH
XJ77w+ttKqnUTFFgHmJwqlxH7gVBHzHc1SX7WaW0+ienNTd9bBQqJbjrQMi9TWWLIpREHv/IM/e/
v83Eq6wX/Swa9h9PabB5cjKr6jl1tAsP5Udq9R3MvheP7nCqu437iZMMMd6AdMp6Q/Ks7VOnQfOH
jRD3eMKiw+g0xpiacx2OIQV9Jaj9eHxjcHDBEXOjsVOax9bQKz0L+vC/mK12BnQwk7RvkC7hA/a8
xi4xSMkfWS6fj69zNPFphJbqpSWaHiwmc6OgEbmIQK+PzHHtG8dp/FR+Nc/TTAetDkdZaKaiubyG
oH+O3424R/zlk/MQ78DUybdrZuWVfI0ClLngGs5CayQcUPcEW1FYZlkHaGKSo6P9vRuvAT97/pl3
lAvAABGu7qfkRFgux+bkpwOJ4A6i8orquv8NnW01vjV9ylpvx+h9FDwWOOKDUayLo6JYWjd5ifWc
0dE5Efb3p5wuOe830iquzTNTtZ+D7wlSIOnqIu7Mo+YIijIDx/DuYv12aRimFqMP/amzxuM+QXV1
Fdf1SeCTIhwoTJsQZVJiCHWvRbcphlkB8xmq3HBXzdtrLT0y3vL7G5mLIon8S67/yhy54PxQZV/Y
0ryQeY2bn64NFVs7iJ5ReFvyjh6b/6A9ckVYU5dWcBVtYh6MKiIbQXzKuOh8JAXaGKRMYpYB+DVC
mKujB25/V+TnkhjBiSEgBrrF1zOS4iZU7LtGIqMQSZZLzVSl3xOpUya//R0hQ+FMn1o3d6VNdQ4L
y7LZ6cMmODk1FrK8s+tYqafI7rOSAsye/YKnqzZAjdO2o1NA+kR55c3Bh+ur5uNwXoP71PWjtUTr
pLQ2hAiPwS1bv5GgagV7idaqOd+ngGDj/Z9NlLqsP7tP6EtN2+yWhsPwzwiAh7XCUoGgGhElOmJu
aqyj1q1Wxo/Vh2mwQABChdMOJP7auQ5qnTSGsrGUd87IiXvKMokVSQN2PyhTduoyWTIzKcTq8PAV
CpoFxxk8hwWrErbKBkEWEmUWpgNYkUYzQnw729+ocLZieS9lOnn7FEeEG1KMZqKoZdY3oG6DcqAZ
CpwJ/gm3z9B4GfTwE0ErbeF7C1Ecn7KaQyvS0pc/fB2G9vbuZECQ7V88tzg46gJc/Y0Ift/1nY9D
juw74hvuia3kAOXgywcPwg0E7qgmYGS6SyyfgxaDKxISwa62kQI+lGluogapgeLKmf1tGPQJYz5V
Qtev3pKvPl6IJRCNXgE8eNfP7ACfPpEtxU7RrsoYtUgrvPSzv1OQleNAJQIaNVSr7zq2SNpBn+2z
6W00w+X4KVayJ5Uvl0HlWakXvNhq0gXVTmXQQsBRXqZwlcvOIfC3SfCNBzcBPhnP7KZAT5C6WOqw
iVUUT64bd50XvYQ+OkJjfV7arBqdUNGXipKaiNw2McILtUp6tL2ypCaPRQmT8+RLK08Elx9u49vF
hGrwgcEfO7TNRwF4ZRL0PEoW9QnGpY9qfgmP0x6NPBIn33+/PoYSabzBJOzF2T1TByayw98Fy6Qx
0G7M5wjXJGKJag+NjMTDC05O22dBoL/UShL+O47EjDPfx0OUDG6M3VYHl24O8BnibHNMEev7PqHd
as3vTHveOM5UjuppF59JLoDTnhGgLRpzvQULFqH2i+UPzVV6cpYp1fYotNl3mNAOsAxs6AyAUR7U
zDlkIcAxLCIY+AeBRSe0XKIISkPSntx+0mMUyQASRL1B+eVLy1ObsN9AunYa141FCgIjoDYnnJpw
Cu0VUz/FafEXMxVWvKdjf3kkxOmIYipZzfYnV9AQCTncWn88RJX6LREs5i9i3CDoJYeHGLRlzMWw
pmK6igR5YDezBSPl6VbTWQFFLrZbaDyhg3u0lu9GVQ9800um/7BM/WZydGaNTDeQrTSPwELP6L1A
T8ex1a79wnHYBf8HvghnsNrddY6k0tgJhLrFk9zvhtnz5W7EO+P7C01Ecl8JhMANjdmQ2TkVL9/C
rzKoaahbvX4OCrxlWXjxg30NtIWWHGiU9CLDLgCH6ekkl0ROo7I5RDEWSfjlJJQh3YuVccsKhaM+
c//z3dBa2Y+nWy14dYtNGA1bWmqlKt2Vj3Lp7R36JRHBrUclWWX99M+u/Ca1jkPPlX36+EMuEOaQ
qlTx8hYh58cg54vDOt9heLKmEvMQpzf1j3T+mGR9rBVz7lrUTgkUEWIJHIIxR8rsArho5eGF2vj5
z3zzOGjiCL7F3vy8JWXraSIF41VULdS/YEgIEB+mRiOiLVVQ6hDGr4b6SwNwwLQWLyoTEB3Twiu0
Pii1NMSYkd5vQOdUGnbr+Ij4ENDEtc7ObL2vhZvbAEWt1dupLIxEJHH6ouauXvQCMwTIBeJwleMm
6kW399ufsdbbTpJn6w2SmFaqlgt5i7gSFstCn1/8n2apkUrAO5XAUkcbcvceLqp67xDGr2Uc+bBL
cGH1u/T0bY+e5gNA/reMqBvJbRaxblF8Wrw2SkYuB2VSW0F5n5vphQzydTsomTERdWkDHPQLDIwj
+W+YjvzTwTlVf60nee4vS2GYQgsef5w4MnCoaWXulu3aYspBDqnj/KtoyCgrzWhMpQJsiznSucWG
UvJtNghv3QWwxN65HfS6Ay0seWtqf5brmoCkihOh8ypi7BoPX2n1K+kyfI4d/AYVVHcPFhH0mz2H
rFU0bNxy8nmenLntbnP/LTW44+AZityoCf/q7kB5Z5KJzQFa9L4PjPAuh94ORaCTaRxE5AJ5Ahd7
GOjrc6NZgUWtRzRBHa287gCLmT1tzoqZiwuuL/PIr/ve9aSGMKRBD2BXJOpeADdOB/WzwFX78z66
5revRK15ZdDR+DRckD++5BKp0wx/t/nPTYO1v0Smw3CcsL6FkY3E1I8iC0BJoiQzFuKrz6O3jbBO
V8owHAXHfQBmPwAPXKYu7dDG3QGbpTzGG6RIr/9svRg+0qKoTRGQsumrwS0RcbaTrzZUT7FAe8qy
gjYG9fAsVmNdZ/0YTNyV5LI5xg76UY0AINAAotXb5Hxa9LeSAtSmlFC8bjUO1Td1kRooBYYTeLrv
X6dt177wLw+wNu1fGXm2Qb1qt+j85pCWN9gl8QE0f/Vnfo9+9RckS0XsZ7WST2e3J0DlHWa5EBKX
V0CXrLwlxALuI132pU3FzsLRIzgjAlr2pE4JR5XmctmnVFkTSzT4vF8NoFHI9oYPD8QBde8LPPo4
vUwtS4CkAtLIc5n2IUzk+Xx1Mp6Dj6cIlUzcX9ezkpeZUuEepqGbIiaE/0tEOAw5/ENNSqbl03kg
6qP1BhBa8gkMlf3Y+oxdRSQmT8WNKG+NvixMTh5uJYxSOrcvWowy7O+pBz3XvHNueyd6KkNdIpyd
evDpClrKHKuB1akRA94V84TgMqhK4dBzictBAZO2M6z45PaPiw8vWwNIQ0GvTwMPsQ35yNlsfUP1
ObpgzAuKW4M6pw4LavZsdex8pcac1Y+T2wPiz6xENknG3/cKY+U8LLhDjsxYkR2+IXbXu7kLzLlj
V4kfyjvzffYCGahesvaWW7UWA3xoS4kkzz7aHJknexH7SdbKwXOAfAVf2TyjCyxFuUR5hfYo81ng
DLvVpFvIS7Oo+xN9QUkr/nfiReXlG2nqEbcFYHvZNgF/1mkyWKk1WwGp1sPMAYL4pjoeLxnwk2Cx
PheXj460mr0wlnK85bd0ADdvFoZkDOrX8UVA+7KEAZak6Byyt3j0+3TLSyroSggdxr1vJlcePrmc
rVzlFU+OcJhEiHXpBwLgJ8TqnOSsRMOF8it8Oa566VHmJvAnc1C4YfsofP356mnQPIB8+72Kzf40
scgRkTTJrxLSZedxXkvdFnszoJvRO6Xc0JX8LOpbfp57DCD1J3HlH9dpwfDAj+xrSvoRLlvV3k1M
rNxJP1NkcDBH7DqI7/Vd2npIiF3/N/h12KPTlcFIEXm+lv6AMc8KFfnfmzk4v5LEmcwG+034dANx
Bj10tj4qvYSjRXjBhrrBtJqELAxE67FZhH7qNQB/8GUb6KmjZwH58DPwoWnutQOd2Wg0tViKo+AJ
uYPHf6NKH7bhRM2PwYkSF0XBNEGuOHmFF6q1PJ9IvOUIeU/PA9gOdpWcULyio4K8/OYEOvEb0oh9
aX3oRGn0zSK6vrgFFyT6WGzY34xYAwqNGiGfAbmzRFoylfX8x0lRASiS4H6P/xg66FT46VHzrMgW
agvgPnd9LMJX0Rxzj0puQY7DKdpCGSuK520sRl+pfpDEqFxRY70aS1YwSQDCtpI29r1pD32C7/UL
vyAXyAJW4W2OrSNnVGrE8QtbLBWOgzhP4t7MjaLXgXf870d2mQOnh3SFZz6FD0Rc+94yRwHAOI/1
K/bUZdlrAgjENLgnHAwNCLdvlAdovbyGrWKnP6pzK7YcTUunNhByk3N+3hmtx8oYS5lR6FwfW8XR
EMIhQrkrh8htzHj8ilK4GpyaUE9129r+iwi4sBE3XGE/9sZSh70dYel8Yf7JZqxgWNWz6DyiKYyL
VLbRxxUFJgfRWyuVCLjDKwhmL8l1/tr6DArvb5lYoC61mJGAr54fMawb7S4donYXX1ALfCJ1cHBZ
9zjv4z6SQ3O7wObfqq/LA3Cs8+9R4s7OdYAZT/tBSo09IZ+AeANCg8H2SPst6bJPnodqipn1aPH0
61kESCcVlKCOxD8PFx2YbsyRPbbi9eNigwO9quMtP0r6jMiTjYlY3i9UIfHg4OxcV+0EWnekYzmL
eVAV0GnR+jI90oXA7RQU82rwW/DMegEFT8mDZHWJSUobm+Aq9vVF2VIht3198kn9Ln1iKfGq60br
wy3av6u9X4gjCyhoz15k9oB9cO5BxIXbkWzzvAqLQuwU+P6LW8eMJMOO/9amMmQhvsEEbWIUMxLI
Wba586AcIUOmEVr9rJBr0+AglfEkm5e62lmfNjIxqGtBQlnykkDY3Kq9VlddKePg5Fim7z7AWGGo
LcCOp3YOQkBUI9k6rWFJ1eaQfHGGMAxxesYI9JpmfuZ2xKCIg+V4YQOx1ZwthwdJ8f6HabIUm6Pz
zHeD2qKYsW0SJ7b46GycnhdFmbqIT0VWahcaYNfEhX6OxkKPM2khrBomAqSEpnbxIU2JDpGzLAYR
6Xb1MpG8QgLejolpsMyl3nqJTee02A3CwODzXaE9YbY1uNb/VpyIT/KPLHuECvkOnVvzDk4g+A8Z
DEmE4Z8Aw5pVizQtFoAHN2xN8P6oHPj5+gY91PWUn/bBUmVZEwMjilVBcBf5AT8KQaXYboGlFVAm
NYhb9eke007dBKjlnxvZMTmBod2Vdllx/vfqjogV0KlBxxn0bvOYPnCACg7NRJ4Dr+S0sSihwyRe
VGCK2GKXJ2O3CuVVPjF/1Tb6RWhIIfnsd7kZ74aZ2iCq4Aw7T6nBENNm4VvkeGt6ackqgmLI7lPW
vRjnOSodmpjGn/1yx6+/bN1SD15JVq4qx0Qkh7lKNgpT7SZeyHIUBCoHwg+r1uLRMYlbtKHuaHfr
WiKR1XZpDM34+1EE+3bY20aNB33wZi1PxyhXTtpfQ80a4NH0kCOs/vahJfeus0aB7cRAySElClGO
Lz4k49nVTd1eqIjFlolXlj6voNA6A/1l3rTaaxBD7itQ4dI6ToDcH2ocohAQl2VpEvbiz0evUXR3
B/BE+8wsB41ImdEYkfJk36/rt4eZNawu7A/+alMljR3lz4JLQasUoKdPsU4uIzRQKXo87MSoPatQ
2V/aNmihWcVKnjRbYOHZVwlnzR89gZSCrvtb3BoUIUjZVJTave1uNqfBVM+0ClxdmgBwJ90aAIek
INDuWHTwu8q90gJSIb/TfOPTaWgwqshJ9SN/8AgtTWQyRvKLEOQR1VwTJbfKMchpj87GCyNmhbxI
fL2eY+ounvD/wrD9031wrthOwidQPKLluXiY+tXoFLB+4etTQQ1B4ro30x195Pedccz27GspFbCw
cyB2OvF3DLchytRYPQYDxqhZKnhmQen+unlTst8MUeUum4Jppt3obVoDQqg5Kjvfm1qmt438C9vi
TqvPQkcLmAn3+nowwpZg+vJ+rCAtiTEUhQuxQagfEUIl3z8tzd80nhFS3xIlhx0lQbS0SoBYRUHs
we/4UOgWp+xL0is70QI/K58/mF4eX5DlA9Fd86Ly6Opew73db/gulFzRqixNwz1m460/vpKBP+t8
uUZM58RyMdH5qkW6KynBZmIyBd+F/LZOzaBXf0M8FEr4y3bsF3F7iOcPTfBy6Pr3tPNs0QliazWr
QmYZ8EH0KoagZ1AHw3CiwNZ1o+kR+/uFzSFMaUJXN96wtO3Q3XbEUNrzZE9PagPrRGwljfzxEEpg
+Q0mBf+tVw3eesrPMLACiqHjSZijoDXkmvEW0u/MGI9OcfGR5Kx0w3yIldGH+qZ+kkGGs1sylMzr
dFnfVVZVSyFgMJfRWusDJi37RMMfW71JZHuIWCPjfy7ChcO4amxiqms/+i3EAGSc2DbNMsT+PTxd
2TXcs3aoHGNiile0Z+q06PaUe69Qcf5mslJTl0O3cNHMxIGuW/fPHZNKQdner6WCO0ztmT3iiQMv
nTsgDuDxjaSp3hetIaNMDtffmJrmQ9QL/RCleqCGBJpElma5p24DxIPDA7SZyH4p+PkTMNmtt5Jd
p9S1F3mTtR/D5sXydjwSl9R5Tfw/IyAgRojLkRHeE6ajDgOfshoOGPWzEsmilzLuQzQgczYd4bH8
lwzbNJM6sw4viU0tOzlnIJfEm82Bypi289sH1OQhDhrL8VUktb0ItVfca79UPZHLbPioNrV9DW8Y
R0TCh3NL4ZlM3wDh9oMAssDdlXGLlyzSZQo/WtanvxVaJCuThga2GwkOh9tylM5qs6EqrgymQe+W
UWKPW6CfWCUG3nz+YwKTiPd+aRglEaS4nR3amk/eO74+/pCeiVdaoQMht2b5nfrcLbTc+v7g7gDJ
ft/UrBHFsRSQxYMKqRvc1o0SPFiOjdafdBJYkzM+8qXjWu4aQobJOg+yzb5D/eUfpExmd+gVN7Oc
EZ5oR6pGVIdCm6iMUZn/MkY5eHdv97jmQjQrk6tpt3sYglnHstDgvBbaUNXzLeeHCWgE2x8YVShb
He7v1Ys2gZsphHPqu8iPlVsuDBEPc+pj0wJj4Qgv7Nc+U1vulokTf8mN48X2hKn4HKS503oz0jzR
i0wvIFbg1gKsjhee7k46C9/Phkf1Qi4lkQcwcMQaqBItArZ5Ig3I98jWDTDijUnO8OnNF1mse4CK
BLagLfTDwudhmCmkDiIqJzF8Q8QEjnxLB3FG7ket49ycErTXpwxRkJIvJT/TKagOeSRfzyzoHpOZ
8uD76z63nIdcb/o3oYoy1tv3ml0ARDaAWuBnF/G8JWoJriuTYAzeKrt0c8RbjHd36hOmtFaGX779
Is0TvDK4HPI3nm4HKGTFqve1D9mFiVZDSbTi/9qbqKn2uFuIzYfQDpsVHNoc+OWSMu+7VU0Epur9
6mhSef5DcNMoOYXX1CgruXQ1R0WEwps+X2wME/Nj+lK1Ch8KQES3Yjz11rLCQAy7PYDcb8Qb9VuN
XJTofRVTkrIy07QItOH7HKGZzSQwpA0HxBMaBHBHuM8lRhVWF9bv9qhK+MzE8upTJ+CvL87Tr+kD
FFwfY2FQ6u9bF4dGGamu09YyudJ34e9QS39vUBT5+tnwrEBqsfwzfz4mBhIsaIthdvDDHxNJ+VNT
+vw9nuGfS3Ncy/7MflRX15800cC2vsTpe/+zZOLbsFCMgZMVuwCBJ12YaRSBQ6aZ6gDEM7a1y9zM
dPhpLr2YI2PAbhtIiwOElE54CuKPypnuB6dkHTAS1ogm6t/rLGd8bdI9bD9HIAJSG/wCP5M/Ke5/
LWEUdzCIIJxY95LrVzsPW09uUrRyuoaiGidHGjCkF/XY1k/HLMHJ7tAZSTIKN15YiBRdrLmGnK0S
H2ZSAzYwK09hV4qhssl4xvIFXHMv5Fn3il0nGQIMbi4cC7CIseg5rZoQ4dmxFtTInsrayjnZ83Uq
BlyECUWXP2wMIWfxVHFH3+difh7agKxSMCGfjKaJoKNCc8qZqOp4zd2OPUTsjgBbAM0K7k/qUmz0
VdlFPEPzpzzl/wwTfMrlNk30i8C6HGDzmdQPRD8qhncBpzxjyxr6jy4HHPR/jr1faU23F00XlTVg
P3SWqnmzEDzGGowKveBEe7o0HK+pjMBBsJonUEs2iyAseRfc2hKlQom62O1tsxM+qgG5jRfeoSH9
X6Ddwsa+BkRLHfvJoDDW2quAxdNBBThEaDh+rSj5vGLfw1z5dLcGZSFAz7zcIP6gIphU9TDCt50h
wvZRdXDrPTFEmcZzsuUpX4fvoy7b01UZP6Qx00PkzoM00COn9l1YdTYN9zAmHPlyfCB/FWOkzdGp
vQitWsZif5Fqq4OMH9tRcgKnJH1/vvMVU+evNr3P/IPKRMuhenQwyzF/dZYrRthv8NyuTwDf9tyO
UFRxQysr1VIXrlif7QZt54gnVQj8WkbXdb8dQchALZu5aYyPvRoFSGLGGgLq6yI+4C8iWO8yMuoM
3Mu5xM01p2YRG6UXdiayl4bJRy4e0YpgYppMKLxGs45RNymIzCdPbr0YvVl4hCC1euZMdZtywms0
r1F5HS0Wxg+BzlSzqTC+Dxk1qxSCTYzqwkRLDja+s/BbjzwCm4ot2r49RVPu6jAkiYk/e6IeGXdf
bQ6q7r91yXyNRbR7MjI1uc0fB76d52IrgJIqlnVwz9GOzhAxGKxnI5nJR7uvinfAMKvN4Gw5jOQU
dB416o6ZsMNIp4GyU6M4ZYAIZUGxolzUKqikAKXbNzVQe8DGugWBR/xvkEiO2DQUlugJRa0Hc3fM
Db1kli7TwGEhrxSflGPoiV6nMRzFrKaPoIVFVXfjhdSVFHAUy8nWxuwhI6/II3GvPEVjKELiwksG
G7LlyTjv/VB/Wopg8H3ull/pv6gYf4PdOonjqiJq1NveT7GkMAKXe6OfoN8GZXoDo1DXd27SAp63
Y5hePiJ8H3Gx+krBG5EGA3t2EzsHrkvWEOjSP+PdJiMOr0kJH1JB4xF8sSNKz4TD6QL0CkrWUxE7
bmB9uPwriggndVLaQ4ohZL+/eZ3FOLu1UIr2PNzwNUy+wafyuTOZS+1zTkHrAS87sIn1tB44N68g
dxJgz4Gd3mBpSqGeD3PMG7XCpTubulcWxmN9KISV0dsJFLWBKGQ1GvX7ng4nRDtlkMBwf0hF5bZK
LUxM2Kd2aKyqnadjRfvovwPR7CJi8qq3yZMVrMj2VkkAIUWFyt4XFdleS7E6bYBpafQLBuTF0zSO
ArsPhD1PgG8oh2k60Av2kBrmWjRJWlbq1YonU33bAPLuo/+9oO28xTo9cQmVd5Ergh4YkbU4IM5d
4ls+uvfTfsCM//vbUBqfjJ/N5Nq1cjoJJSbqPJFkHzcJovbKXPhbwFqAOtfnnCWfxFJsVCqFFLL2
KInoe+7K4n7gTx7RbuyWPT3QFBzEkb7jX1MiPcKgugTdceaWl/gcNk3sxtKzRUI0umHilx0VGqCV
Gl+/u+nl7siTyzYq3tBaxjLOlpqx4RlF6y1Bi1SAcIJlAKh+u12IeCasg1dfEMX7jPy6gxnj7d//
MVMAFWsJAZsL79KHJdzn3FVIP8+aUb0IwtseDSjFnD70AHWjNl4MyjtPN5uXu3Uf5xG+ujo4wswe
EzPEN4WurmK8lb26qPdhPHWTJPu7DUNaf3icxpy7ARdaS5Ag/PL3Vw0lePE6AuvMYjkvZGhNYpC1
bPczqyA3tXbT5X6wKUNziu/0qVo6csH8hSjOsEewMiUmUi61Zi2yG4y53ndqYKkAk0LKgknS/Unr
NK0JdWexjX7la2AxDso/o90szpXuwHG9wS7DRdzz4tfOFbvg92whc4Zwhs+uPMUS9hkRmuEzLyoI
VZdgz7BuvNjuW4EL7d2c1vpugLUkC53JOomwZR5swbYArgFZcAvkOM8wOXZD5X7cqHuQ3/oa4ai/
KslE/EdEkN+wkFtD7ZtyFCUUBJnV0FfXe+uoTgY7IaChZGXHud/F5Zq5z4JXPAgYjbqm2FDMMQJQ
4dkLj97AluLiBJR9ONyw+trUWX7AoAp/o3tpf5CdId7AwlPTTh+Yea7hlQNEPQNOKwyPN2jSgbkQ
tvmNFAtb6yqgId+rOX11yA9Nnk5eJxjew0XCCaqrSRBOPrn26O/yJtOq1u4m7FcSYL6vrYXtnQVU
Yu7IwsMophd9MHLo13vWpt6qRGTSBWZV/Cq9q0vAAxHSUObZ2i+6PocdNfGDrsC6SrSY4Fydxi5S
+XxwFV2H3Jx2CXGWDSuqHvYvAtB7Is2ngLHbO3WdsAgK01T+4ZcnouspqI1vm7L6Rby3zQ+VgOct
S7oGJeqFeQTrtttPdHc88lQkOUnNoPNU/W3RPeEwfUfcyx88cEjTn/u11QbhDJ7GXlCj0smIvwAJ
FWU8gZxdksJ3x246YucdcXI9pWXMRhu7FXNJPCcqYik+M9c0IbfUM2SqfcMQ7hy62qsrHeW8BI81
T+5GKfgHbu8NFGFv/i+EDxCHuLeEddNg/lQOtY7r23fcRP0Tp4Lm74HDJPZthSt2OFBuqpJWYYnE
nFWwypVo9wFUZYDM1WQsBUq7c8SxBPqv2UYZOTU+LQxLVEqbN4CqZ6Mw7u5YW27GxCZps3wzH96a
9flUzLWVUaz9GXmI9LMdDC+aVIQclvJx+sdFx3TfM8mj0H1tIrrB9DZLfyztNFYis7emMKPgbaDJ
QDSPVCJmnCIvoXJl1mnSFFUZKPzCi+/dZT3sRAa7nVtNTAiCNBmnKPpQUKGJggjs4zcUJ48Yph1V
wjsLJ0ADtY0tNqsv8ljZjDv0HThPpBnwAo74MxnkBUI7g/9pShkh+4dLVBqvtxZ4OWqR8e9uXrp/
jjVGUzV/LqR2YqPwrxubkNhy2c4T3HQ2EVsKJXgn+aDYgGFDIDk9pJt9GFJeZpPuXqY73Dm+Jv7n
cRYP3AbwmShQ49lV5EmGpI0H9988dR9crK5DVSwLEGA0Cf46B2WNnuyIePAluikU0kITkRavTNzz
XEHmlfTS+A7kFO57po8pd7mMVE4/tooZgmEskKFOO7gNtD5Eab2EmwCr3d88y3avK4scTWgRuOBr
nQnEYWNxme/aPF6Fi0uTVDx2FKZYocwNFtVVajIFJj8m1iWo+9NSrzBCjo50hl5UY9zez7POtZ1j
tWUcTnWOjPJYXy6V8kChfAVjWugohbTHfTtTdZSos38ozFzJb8IZP6XG1dV585bRr037CM67sdXH
gfivqRWD9JJaCElJM+Bx/ZCQHmocVUwDRxvhbP2ezOT3Igyas9mcZzeFidGpI/K4IfFq779n16Qi
oE+X6G427zlS/iMNB+/mkWk5sG5c7uKQzV8fp1dbGm87W3expfUt10T6O0GruQgM7lTXxGp8v62x
U6Qo3x8dtRDhXxzraI9rsonpqWAHY4Ow/h0oCcYzCgCDKS1zIa78Vqp1HurinYCCvCUDcvJp2lMD
mGwMxHWHC/+JrJ5vfs1bYeto3TJwi5I9Y0RBDOgC/1vhiPixfgdWCykRFDdoHLE+cuf+ouLZ2M4Y
l5Q2SQu6tDySEO22NDOJ4C8TEURMH7jODglfcrXEg6ad9iym0+PgvtsEql7BKrOtFLwlvM5kEJ4u
XRFYXz9/7vLrz7FwjyyCWzPyxgjXozUVHdSGCyfNXUJqi2Mn8CzNtYgCKhnE9/IidYtc5psXewtc
VEwHHYlENMwY+2fvFRtfb7INRysgyXUXu4giiHsAutDRLNHci307TNizX5pezOouaaTwHyvDWv/o
UF4D6mthNbNDBJOwD6t8PhU8kmOHBVf1zYVt+7W0bGwpvEqUlmpVzjHizTfzDxABTyBxCqrYUXwQ
wVwJ1WCG/lg29f0ruyNXX6SkRoezoL0Wdg2go+33rtZZmGdjlWDTK9BesMmscm/D5jdTyd9wq3sf
wFrhmSyg2Mjo+uPBf7UUlqggC9mciwAJDwlbmoLW8xbYZuprmBOz657SIrztWk0m+Bq9PB1dMLqL
JAnDiqymSHxket1VtHMJcvEi44BW+GjZqSE1E8srK6Kk+iVY2jVKQKu2X3mfdHg//PrWrgFEMy7r
DAk88GRPYUEHxy1izhIAEQU1dlWdQiX5iekv/9V0kCG32FZk8fS1eu4Vq7YoloDIZTxgWFCChZmW
fV56XaA3JtTfaMnR9gzSa/cDC3SPFtTGhMU2U0Y6djZF3YJCeeEXP21H6zbtCCMwi2Tl5NetYIFg
U5DIPd44sD8AR8s9qEOOoiNioPhhircIDnFsGEsNg4vsWClKATYcGMTBTpwJefbaS/DccJNmhDA1
iIQ3NYuGwi69bhSfayEIUGQVDuCP5N7+Od5fNPWhAIvJ+vee8i3ADHz/dBA9QIEwTpKDIXkwMcyM
uu95l/MkhLrMWJkCF6jchPvUP3LddOSm2MNHRHyiHkHFl2jgXA3tep9rTgFUvMvacoCei+rVBH6O
yvn720qMCPibDS8vkUvS+pyt9ErArS2FmL+Qq1sJIBp5TPCMZ42nc4YF4nlfuKspecUKGIxG5YHl
HFBW39cBClNhZVXIAmj1F+RMTwoSnf6TkZQGsTUwldBUBuWfw0x6mLO6nO7plZUIW+0qiJF9FKMp
aXX8E+LuiMsOO5XDC/d+ExRpCQu6IrLik24jQf/lnq98Ij3QngESeA75D66z+6rG7is5Nd0ekI1H
szwKzpbz+kLrzhCXpcAPydXKO6wV8o7HPRjiABooAMKY96R9GB4YzGHPPQnHcsCkxIwNGAuLPhXe
Gcm7KaCoARRfHIPsT0Zj/SLg0ewNuG7BqnhrwJX29nfa4TM80kbJyTtX9VhS7a7rlwAtwBP7zSUm
G+XmvK4u5C4QrBYRVdv0M48PaP5qOa/bCSIXtDv0rG4rjNDoUOHPq0Sn9KJOvGIp26N0cpqTw944
r46fMgyvFuYyuuUyylsIzyH7BBzbrqebDNi1gDiBlyfOAZytT+QDUL1QSITyD/claxeCTNZVyOAi
nDerLBW+pkjV8apsjhy9oe9mhy9N+vMNljPgwtT3upcwZCHr6HjENdSjd7Z47A0gujsLa6at4heW
quiee+GwGjY9zYMTE2MZS5zXYCCWiDOKe0nrGL8qpTxZZ+xEYuTO4UuD6vNX4BY2Zfvqq+L11IYU
9lYBOcQ2Y3+BPsgyC0y+7CrZMFHsyti9Qd4jFqdSgTwslar/Q98w5VghrTzCIIwHCwwRjL5y9b4t
V2ZXGBOmwCKFQeHdVF63BUuHqScIYu76YL/zZKuP9z+Qv0HA0pJ1fRzSNqIR1y0cptWwfuU3bNla
WM3hk6FypvxGYYUfM1e+kbdFOds3fkG7qIwqF7DpqgcL5DAb9ZkJQD2sp+kaAVInRmc4/thp8KGo
mA3rsK+xkXu/GsJp36xshVW/vYOxshhg8Z4/dt2Y39ZfLMC3dzHHufIVt2MJAvn+Gu5byxytBEBd
o9aokX3h9Y/gATPGGZdKckn8OdvbfYgbtXmnSz4FJD+GEsYna3vswRM7exp7pIKWFYpOjEQ7aRsL
1W6mP1/xb/FbEJYiNq2em5admCtxHcng9z1Sl3iTUUvj/PQ5srWnm1TToBWO0YkkDC1ddUQb0+zY
DmWi/Msj49nhs97FFnzmYOCW/7soWt3hz8kmSNfMsG6pjH6+02uoWtdzftxO6ObwbFXB5Rah1eUs
DX1CdwTTHWHJRcDILMEdjVUQmulLDKXQeyJ8vLBEccHPC67fdzYJ/DZeuF0aOUBpisv5sOZHCOyk
iJUuCWI0xCyuZui4gW9Omn6pVtu44ct9PummwQa1Zdf117VploWnKpM+aWSgodVi4xtUioT213N8
XWPSAVNl8rtt3mxtoABCFZZ/SV474D5EiUv11aQmfC6Fi+SrEuj7ZRXymCqPi3cejhBRgfpGEK1R
agAAlBrt5K2CC2GKnZUx+ds+4X7UGOszFgHHfjbezcZrZmraEPny45xc1PfkZeo1P9JP3tIhGt9c
TyyGi1kuiIf4ZWkWuFweMhhzHZrcoIDhmtGfDISwaghQsgqJWc6yHAizeDKY/R2ERzGwSyBzMvQv
YPG7XfV90qHX5lQjN4gKHiMZ/Zh2T/9P3Ssjjm61UFsWdB/AlXMs4rxLVe5fqPAHgGy3cl3CkDJ/
iCEwXZujL6X72lkpnr/3/UbdDgy5DZqMGkaK+CZxPuLySdqrl6jYuDTTJ1kFo0/btS92VJfc0/w0
XTQ+FJk+oOnMLpCFQHixwoh/i0WswZ22lQJ5d40UM9x72OPvLK1c/JoEgxT3s9N7OKnQpJ+vuYpw
VcN9gHs2a6DKyIaTcrS3FDkB39VVDPAVQVYc1+lk5zimr4frqJXvBzwZPNl6aAsCiZJyVbd1CnjV
RvnXN7Aa2HhgcMcRZn3qHIL9tNZGa9W7rt5xAqTWCHBe4m4eR728EZh/U4mmhs1FdNnUpWEwisbJ
JvTUWrH7AQAfYAOOT26OghlLAL+fzLXLovxMrfj7HyNrNMWVmZK+M+R/yxUy//Pg2QijuakWqbu2
2cOVz0LhMwKEB6b56rCmUefUX/FHgzFoXF2+pwhXv9SSxTbDga4/g0D5VjADK01OGDV5GJ7otOYd
YfCHEiVGJcNGr/mkcIj7WYurxAAughDAzOc4hfrgOqJQEB3x2niZD6Qa6J3yaPqG4B6y5BFC7fnr
FcLcRXyUQvUIWKUASisBd3Ev4Z9d+lkNoezpP3NV0qcZWkmP6KQZtkTwr0vMygC5WuW+ebosVsMw
t5WsgBJ9HMZmyB46c6fvWG30jT3CZycqyq4M+QQboX2T6CYYfsCopRYFu1lRM96y8dIljdeYQ2hA
IpL7ixfOGCPKKmlhTXyO6WEDC413LKCDHRVp+3rN6iYD2yff1lvd8C4GYbadbZzKju0k4SUO3mSr
zJXt1Hj6FDfysAdqJm/E/UThd3sUpND06mbZgRlOwbQPPB4ObDxPFZj3+/HUGLl10laXuwQRFWRx
0aY+Y7WdV+B0abOjn45pd5zGlVk8Lm7eNHqYsFha/UxkIoSVEEvmYWdec6ATeY/D8GawnmX4Gizh
M2HjLZxUP5xaRDr3lPzinGPo9BLOr/6GWtA+U2T/GjhIL0s+qsOxZr9swxEanevkOlCZRaPfJWYk
4R5cSdNUqpYbOKvkpStHZCevfgrwD+S0IsUTnWS54izCqSe1EV1bh37T9m3sjAapqfGEO1tX6GhH
vn63cH1TG3zzWEK1HnO8b9IsmvBlZum3/q0mVUKIqqYSI6hJW76Uznz1VLClUm7FGuCCWwbvOvbg
PPCPBW71eIMuI82Rj5I5EfMdkbVJxyAt1u3WUcN7EVEhyeE/Dx5zPss8k/EMFUIfHLpeehsfctqm
apo88B4hlOD2eULPmpPQqSnuZgMLnMbrh7ms/sT8D/koiX5KZ++C+7GSjxQ3d+RlM5VVMwF8Y2Bn
xYnRhAF+Ed1fYceh8fcHZjs6vvc9mWiBYQlUbNsRTu/rq1liDihFHvC7Oji8hezXQGuUUbT4jfAq
zMMU6mXKsSnts2LQkbBf+IF1guj3WsZbJx3vluSJj71tmnUKoox1YJcnB/6XlUThe3Rz4s2oJz3I
F9SFtIQ6PD0L4WiFG31Y/WTw5TeW/WN2SKO0Ta6Hs6KEw3PC8LOPok7CXkyI5axVQKsHJy6XVXsy
FL4P3dbg/FSq7GEbqpak5NhMf+7GUgDUsdD91lnt86KbWPPTi8PxRemqkDuoVohJDl9J/XKQlUpi
sjeEowVbdwkKQJJqt3jXmp++1ttPjkP7h9qKpAtxaQtRB/k+Bm6pXvc5HSEr8XSTvGBeE0HBKigV
sHsnOEQwBr3UedxAJNTBHWx9nlDSl4yQeX/bm1nnlrafg2Q3lcFHqfXgPE0yjAS+vStqDA7w0KvJ
7LC7JQAcof7RJW1EYfuy381HPP7H7YqoyQEw88DEBDHawnMzhhm4fF3+3/1Yn0oJPSZLT/RZZjYT
5bTQ+k3EgaYhW5qKs3v6nYhXis7WAxNCeem1ygqB7ajK00p1At5KrKgaoSgHRP3IBAwyAWwC2zoX
onzfqXMBTzTU1ZzTBQMLNhCr/qyN8zJbwRJ0rQi19h+XfkBKlKZqMrhpWbZIt9F/vuL8mstlmccc
B2SEVoN5R09/wgSx20ksViReBJQLziDeOR/JoJrVjf6l/4X4yE144KtQuZSjfd5JnKlTxV+vRtWv
4dCu7w1bIKG2hzC3IZ+jLkPockoVtdSGMemWsWU5zUTDJPcx/3a0b6Jbkr5uYyXG9y6LnjJQv5IW
i/EIKyoM7jigSOCoEKL8xGWjvoCgITW6XRdG92v+QV9cnNJobgPSBvBi+ZsxgPhrVZu0QqoGJLVf
7WDN7Jy8iSNkdHNWaf7xsJtuUjIfVylRfuEXUkxzW6fzZJJ+HEihU4aWMOZMbeyN8XciyIgGusD0
Z8fxs28Iqj1SryBZSyogfxnRn/mDQw499MNm+3vAceTjT49AyLs5fhVueuJNphjaKntUT3ba8SSE
mtS4DvED2JfB7MWXVBx7bmicyVa+HgeOGgAonuH1DdWOKCs6XNqmbr0XElnE55U14+adR4ysK+BX
CaqSWomEwMbSR3NVwNj3fI6+XJNEPPMOR0+6C25Z6jy7LMeECZqV3P43L9+4aCzyh01FQS+bSAkU
08ovbvwkeuRCW69L/JOpl2GHViUKJYYgPd44TzpXQ4aZlHL0NJmSo9d9fPYbA3xGo5vY/QLeW+uj
7pqewS47jlghKOskXQ+1JvIWwPUxVVkWCsIIyJC/Hfy56rCdbnJlUt8iWowzSno/i/D1LBONPSdm
50Wvi7RmlTMcOlyPFj9Sd/+Ad/BZEInMt9ZbECgHgsxYGagr6pRKNHYCdqiiSiLskxuBe0mezFWe
z8PnxUIfQAauyMKgHDMqQ7Lht5XW9Y5H6Ra46rMBvxoe1ZhwDFvmmOhMdfZMLFnQZ0gbP4a3f7HH
47trJhEYejxhQUcbBhaDaHkLTQV4gMQOABrLJjnuRGDRDLxq2DOtvXRK6Bel9F5ekb0yNd9yhX8N
pD47pBmqTXWrOZ2x3l4sDMAkeHoawURPSvgN41vdGRFJ05fPXMXetHL38jSsNGJJYJ8Kex03XC4S
IM7Dxkko04mv3gO0hU0g7PXlBi68SgmPzRnFoMbv9N7Zn2EMslB3r5R4ZeWfCzfa7FD5fLee2crs
PU8l1wD+L8uQW8YYYT4eT8w8/7XB+zJsdQaK0qioIOh9IKjztpLVBPGRTPI9nHBtzrisB9Lx8chX
dcXq3duisZPliNG9dTbR1FlETcVNFDDBqdgmdyanN/F5t4IAFKKhJwNMCtL9jm8EgISJ2Y5nvxaQ
n2H7oKbTIej3khd/nmRfqNBHBck8pSNM6UjAHcMKJFnzpMPqGi4cP5vJmvgf3CcZxeP5lPQQ9efV
e035HGNpbE5ZRbfBRLpXY5S5MqGbV9aIZH373umYZmcCOWbI3n7we9npm5EvV8Qz+/+95RNTnWIu
fOC1Kjywa15HAQyjSFwdjKS78HNkxDw1qW1dLO3sunKXOyNvJqSPe3KXVAP1dNLJY9oVD4pMwqoX
WYzM7V1Xw7AcvXBqa/pRY89+AWzv0TeZ1RtRxrONlpah6/d0M3R18MFttbA77gsV1+dGGycB3InU
Xux0tyYy/kzl9fflsLZGciWNqHmj6k25EV2TAb59IVSKCCpfTdo7YeEKdjCS0QwsOJ6WD3mHqfhE
+FbT5IqebcITd6d0xxZthOYhliepGZPdWHvl63Os64h72I1Oy2jEc8tp4bQeFmx+Oa7CPDdlex1K
O2E3zNwUzYKb62EtSHjv6i2hM0boChlERBhxJ3PnF5hiXq7mHvlf6N8AR7oGQR2jx1IozhFHbDv3
CZl09ZKOicHebLpQyYCMWTCchD6Bnk8dL2rIx7/68hJ1c5i1C1hFb3pcV+zqLDZ9QUCUwn5SesYO
IOkRvh0aBbehu6RNNwAKqWfsa1DUm56c5IJM2SWeZUo6KvyRCvC+bCXqQffdYH3zdtKq1FXxxgA/
Wo8ZF0uDlvxt8VnORngXxzF2LRb6G+wy8+0pYgTalYYViIxp9EX63oQPXj846QVmeLTjBkll5LcF
0YFDzCm5BtyieQf75WCHrEPBNp8afXT52gPD6mdoCj2+wZMo0TGKjFGYrQdNv4l3AkmHc3/F3AuK
hyVFPWbeWk8BYf72NflSbbQSpFgFgyKnWfVFbfNMGBHQnwmIhyP4fbj1fj3BjF00SiaHSGoBp3HY
sVAViNDbk0ovKmdnm4XQrh35q70baX5497asZUYtQbuOVG9ya5XRSOStrE38tUQ1V6zjtuZ43tcH
l5b7kQSQ2shYfzf+5VEmK+nCC9a8G5MwfUOOnLYK49c9dJvGk6d32btqXsOmXaXvRUC1pF/tYDau
4kvYEMhSRO631akfYjYmeLHlqvbMDnpDDEglPWI4fgiToocSQYNwpYh3LnUvPpROgLCzO1mu98WB
3wdxriJxDNV1tU/3QiF6rR+qEyIVpIqD4CRc6sfCfpZCCSLMcbRi1zphCNy34Z+RUforZcoQK1HL
zBZcEry5Q7zP4drnKJqm8oiebvipmctWaynZo0iWvivbiSWzBTyUhpmetLKR8aZiaHTInKx2aI40
9c5CNgFMczVLgNczvbL/dBY5W+QdiiGV2xxck0XP0E0gEZYJ69rI6tNBo7C/kjEcD5zn6a53uLnl
NOFZk48pva/OMKAw/oRrud/bF7W7EKYkzHTdUJwGLppjsD7ykW+eLzaGXyTgjDI9pG9cS97m//K+
Anil0VQF+FTkowiK/CF7/sxbC0mbVmPKbB50xS3CcGzVzQCHRWc3JVvSTnRF3sKqPatOn0ANiTFm
qLNwZ8NCjoSoECJQ9gH7EvSUSBJPhnOPiEUUMkh6ywNFBjcF29b8hjW2uAIAi+qaeKb/Bptn832l
8VAucSM8l6NDYBRBsWc6DHtMFkP1qhScXHzGuUAIT/rh63DpHcElzihEI2CiRHTXDsumg/eMvETr
goZeAowN7+25zXPhmHKdVU2wZo0YA+BkIPPqnFULoNI0m/3WHM75c8RSm2imqCJ35h64sxM5iIBc
aygFUnhbjHvhqEIS1SN3l6MNeQ6gWBZCl1D8C5cj103MZbmL1THqIvNPgzZpsuic0wuz+qV9mucu
0AOdWYt33pIJJLehLcOGzW63SU2CWnGKeS1EC70ZfExInT4D4eoWATL9HHd/QdSP3oNcCkjv5zNZ
Xp0qbzY7B7ZTdKRnv7p/qKmc5tL8HtjkQrf1GK1pN3Zyfhb5xh7tZ2NNFLWIMZi0hWUiKACrgkBC
hu/OAI1C0jfzEYIdbYZCGlPe2M1aaItcmjBTfamnx0pk/C9n+A7xScjn8/lYedKOS9Ww29Hdo3ie
h1XWzwpkUZ0A0qZFvLa9GS8hv6LN4NskXpbcGPXsbQRUzmV2Nv0ti51DEuKk4tVOaJksbKsQgq3R
o9MaFW9st424Ld3Se8fmg9754GZHfm6i5ZjeBT1cW4erEqPi09EwTA/+R7HhoarwFNYIR6BaSG/d
q99F5z8a7N7kiEXL+NbYU0LywFG4nmhXy1rIXoeSLWTKC6dWHU5EgwO3KVocKkvfe7Oq8A0TPY0E
uQj1ymRULJ3p3XPlCDkaHdead4maXuu8OEjgCOq3Tl6+OAxWZisC6VF8iPI0s5cSIsFkOibD9KhS
MJ9fS81gB00fK96wV18C3W1IEvqa6/IjDwoGsYwl9QA1AqM5jj2/0jmfGQaYoUfaKWF5ybj0Fnud
PMooQNSdXzNxh+x5EFSbsjF+8oFW2dKwmzHOBSXVx6UPx8P03+w8/JPfpihaGY7B7yObK1Gy0ONK
zFu+I6e30WqmEEL60iOS7eMfrXSi+h0T5Eyhp3AhKRAUixmKBcwMKEocEdF2kulAUeI44nXb+oXH
42x5bOzeZKW3PeYjg/rR6MOHwlf7hzAP1aOpZHyXxcX4O/Z/P+s0MMC9lBcotbAIvBLoGj54HAgA
27flh4J4RakxOtNjwoBSRSka9tv9yqq5lMtYn8MvVP93qW0y/Q0fk5mA6U9eafyl+R5PLXD/HUxy
r5SXJLopx7VGKo7A9uRn4PbaOb0myq77jhQWS0H9Sx9i2HgOMBLVrgXqvJJveG8yDC+xPlHdZ1mR
GHSRWXfweLylDQZ40yOjqp5PysVJO974e/VIXcZ4IQxiSrL3sfbiMInPyzkDrlI6x4SHz0XmhlwA
LM1eqiVJM1Z6B+zuKxXt6e/Mb7qitXIFvpZrqeOnTim56MetxAGh8+POx5Ne2Q6ogCwEhQpN5G7d
/HR0PsxuypsNtqLFtNj/PLCeyQQ4t0O9s2E32Na4sxKlj+pur/c5rAMPHubkBJL9aqyU6oD9fXBj
uf5MkhT4pSkrya1i9rMMthLXggsjk9iYmmLm5aIcEfUwfdO8UBQuIGrazCO4vy8QAhf/C5oJvDit
TyOMfxbTieEdrlJa+xgrkuJzxJWxMDBSFRrKi5IsYqEjreCLmSMlTT6FU0ioo+BuJLb/sXxiC42C
FgelS8cxH1FV3lIJkFVvUeqtciEiaFZCzT+Fa2XAnTVX8aR3Owqv0JZB0knpNfbmwuIw0OlknE6k
oZIN+Dyy7H8OxXM4lrOElU8bTtuVO46N2gJoJEDr+wp/s1u3AsWWQsCOfXIBFearlnxAhWNI8SYA
IydtwXZqf+Q9xZ8i9jdE2q1xCfq9hkbPy2IbP56b+nWuxNEbDErKaoW0son9t62YCwLdlmBlCELl
ZhmSZfTQRjlevTkia+vPpf9QvmxaAB36D2JNhwkbVqYlsquFzwNU8C8o40vClCj+d1pbm0Xgh8Ca
qhdxZVM6Cm0daMivptuTKHQHD8qPp7zgKrcjPedhP3fELj5e+F5zvbk4Vts+8oGAqiDI2L7N7Fvd
Z652OjHZcegPcb5QT1MnQjYKU1JaHif6Drw2DfycwWa9fV08hsp5hjlVVTuD72Ulnblw+0nXACTu
NoF99Jep0pvzc2FOeF8Z3hMXcj1hDcvIwtO1g0tZyyheQLuLw7J0NVZNe5EPeFydV8obwCbCK6H1
a/57j6JMsDhCOKZT3bn0hh6awd6Nt3oN/owT05yJ+lHL5U07By3YZnA6jI5FwyeadHHCx9Q8o1Ya
IfG+em88ng8MKdUlcxcNKvDPqEweY8ccYuYseTVy2WQRp5c/tqYygUQGxJErde+rrbW61tCQ2w82
B2TISnZQ6NLSyI0h1Gy2iFWbhtNBCfe1oEWvaIKbgB6w0lfm6Upzls11Sm+MznW0N1iZONVJOYO1
zW01op7xAq9YpbqeO5ERkRMfkcPMP/GYD0vaXruSnNsc1mY+JAcwkN+J2Q4UQgGimq+IKRybidMI
MfQi0nI/lha/tMmQmND1GfuTUuHQMFPW/VoIfNN6GdB9XerHbADxzy8+hL+lfAzH0wSXgfSYteQV
V9HHx8O+5yHz8/Tpd4Y1i0HQvHG/9aqlqNpl1LjhHhjnNa0L1+UELqtJ5Liv2F0pwUOlLn5S6A9M
LbvjHqp6PxKk1MuB5mAjpLha40EGeG4ldYHKwcGKngR5decLZ0thqokjyjBU4er+KNKIRq+/HSwq
u8Mt1QQO9/+gNATSvCLHw8fXERTKGn1AdAqk1Ei0ctolW7m0NMmEjLPvHBii8FaWDys4eAmH0+Ie
RAjLOaZMZlYtbzZ0tjASJMD0eRZ0uE2e+cNvlRdaaZGB2Pmf0mNrvl4M7W0LFqn4TvCoWWVW71Oa
fp6BWmgBT9BM5l7GqSOdmwM0zEnKiasIinjsQZaohnjQx+PIhdS/XSb+o/teOgoNNF90Z3LoqtFa
TrYhHLzYbrLyv9vEqK4E/ZaWO+GhySU/NdR1RIUtPbhZ/IEv1GsA0KLiV9Gl5OTRIfOK9SjsctcA
9K33G+uWYo+9OmJ4wvs6ZbiOgUvSkM9+36+eeRvJBOsQJQKXrrYMDfAZXII+XZZh97hBEtD8TRtG
AxWSv49LfjcQkTVajrD2p9PBXbtrg75P0R65hTSIj9HzuFP1allwsH7JMEiL70zowEg3vipi8Emn
o058vp8MzmosdVofxgTIXLHXHhN/i/lY5lw6K4hlFw06beuXONLz6aBQlmvLSHixpM0mX2Hfr0Y+
qICnMKkDjG14mDGvyaXDQGcWIdGNXUvvZFaojf3F+PWVgNgxwhx5kY9ZisZdWFR6woWFkJLDRhaN
BKTunIwEIaZpJM/VS2Me2G6FWGpSHn+zzEjJsOvnVXVECuqIl8FH4KZkzZRE2KDajFcRzLxshN7i
P1uzBWaDyBJ66o/o4YzPB2mL6XEdZ63XDbMzjAxp1Mrxsw4MuTAt5bJFwwIBC0AZ3u5uXSRnXzD0
i2eItyq6B6fJB8jFlIWHtUQKcwdhgJF0GRRiz8vVnivhIdmPwdK6L7kV/Nqh890RwB6hOejUaP2M
mE49sM+Pp3wCIPxDOTKEXa/99z5rm0zD9UCg9+DuYaABA8tKdRAwufZ0cYNFPpASmhC9LblNVcGp
k7usOcr6VkKAuhn5U9E0eCBZ7WBuxPM5jV/OPoIA4MKoCJEgnZe4Uy/uM3ifSxeuK3Hk9uqDtsGj
3eUsEXYQhbhYUnHmuhiiXGcSfox20B8Uq+s8mW4XxE29f4dzj7e/qWr30ikqNEPaFjLJ78WBdiR0
9hgrISchOTBxWzrx/Rm+He6zrY4BuVuK4YTC+JVzr5RqYXBAk2x9BnXIgmVnPB2/wjN73clS84rd
L7aFs8mY8Q7ppAUiaBZmePnNmRmmmJaPOeMmC6F+vL2++ZsvzwLhXMsDMDa9vOqRxYGq8xWK5n0n
Siut7QBeO1H4/ZZqp2bBKWd51GZXLuf0xNH1CBGZ07rndZIVjIoVH3coO6CUHb5vH5Zb9ZSQ0tt7
sXmKYiYmB3hTN4oHF+kR+gZJrJGXJ4qFn9u5gDYBRVOY5U5kdg7ohxZEDQm3+jBGqvdjbCbHP63D
1IGRvcgQgJBwzEWK5mqL0QxKby4humfHDeWfF7YASw3K3aOL4G67RelOiu8eA9p/BHxMgHXufUow
TGGKnmLFGozYmB72fej5SBmbwSYOC2LC9Lu6VVaFqNo/f8dyw8Eil7w1QasMddjCPJjNRIjd3yx6
7tA8/7KJoIoVKlpaYkZMOC6epJXbwCefpgFkZ1jP70kfQ5rauRDQiYPoZfvAt4OXc+S0hxw9FSYJ
tNkob6v8whiBf0gp5t71DV2g10DKsJjAX4nhhJOVG3aC4kAMXLbArROcO/JJG7bF5wK6vC9NpHRm
+UTYgBTDU/XEJyJA2/GzuedTa3QFitwyZ0brEAvnIhOgQn4Qc3jm5JE2cVnxFMljNq0IlTgYragQ
bRufNcJO1X7zFSWhzFWt63hBAmsyMcG0BgK0RPlAwPKo/YwSti7puBE3TwzUzXsZ1N5Dms24S+ad
PuNqPKpewm4hp+gzlaXTVqM1XRwMbJgjS58n04UIhmMSNdZuPMGOBtUvh5h3Fw8+a9VO8YX+sZgV
/8x+tLA81usPB0YYRFwUCAgjJs3zbxe1/U56kWWhHalsBp9eh4mboVd56YaMiaCkXPOJz+9FEazm
mm+fDmsTdR14mmlvSfthBAunUlR6jqiHmx4vbdesik1ZZDPDG6zSoI3ITnpmeZ7gT/0DnQnonJS5
FyWXbVUpslcBTaW2ofbHwOoYWRtIG8mizkuSvCQVm/GG7s5d8qAsPJhicDJ9vwyZYBioCCVx9Ptr
UwwN865h9JmK4mZFAAlUiu0Dx7ZDo9THTomYFEfwqwImX1Vh/gIiPaO3JZhFp43RzqmLdYe6trUo
F2IQ+TyKQ6VD1CO9PglFh+CKS4BHfE8djkJho7epsiGzN2hd0fucnR+eqV7uJKzTduLTseP8jI3c
LwNHrB8RqUEKRt5v7Wf+gTLJKmieg/Oxvt/ZLGZ8y1GrXU1hBd1I/tyXyTe9Gzc+mmvosgGSEPv0
v/3SaOKxV4Z8f7dZQNy86T6GmDt79CO/HgeBRrcxeto7yhF/zAfHnkTYu8Lm3RwpefQA8rTmhA6w
+/fmzu/hB6nmkQX+fbeSHcL262E36evutzODXLP59SErs+9XwHug2sFcXNTI0T+Por5or3cK5HCX
KX7jXj1FEFcxGyiML1ChoT3W9GN/X5+SP0oHJR/2Cri5uwk4bkcUUkBRZjDBpFzh8yDIrQEZboz8
diCRo0JXNN+Yrj/t0DoSRLnix3MtDkbkx/xbW+vS1OlaCvzfRpGSzOJvhRHA6KNzWNH3QZbyivVH
isPzwnzhER4coUXQJwPAU8Zy9teYxLovdShJ+Dq9fkj6xRB2PnIkyN6ZErKJCHUaDNJLmezK/3vU
eUdOEkkTwvUT3+L8zKsOCsBSVa9FI5yODICtbCk5N/gAmbs6/0iN4a8JRf3TTMOk/dCwf9c68na6
UmzZ44lUxfg4FprPArdSGCkc+AbxYTnlngEgapLHXjjBydHNK23LZWx2NblirIPDizNh+UWUzQqw
JIh0lfQA8ZqvwXQUee5SlIIb1bH1Svs4OJgFFgY4XJYCA+DXrxQtPZS+0G92nQxKbRvGWA6TjmOA
pFCL1DQNeVUseXGbqMPdQs9Slu+B6E9J2doD+wVgoi5ADuo2vUimJaeEnAOriBIJ5mBeYTXt/Iie
pvKTJzPsWr4KmLbBUvPDALxTYlPqaXvgZ2FiJOBkcnkp3Q96mXDrlcelPIRz0nFJIosxVNaOy9da
phcbXYqiQhgp7wxwPD607z9PVLbzrlLiMmbSsKDfWG+F2klwVljQ2IftI4qx2e6N6RhamG7BxL4n
jpmTyE7NmC2btDj53JgsKj9KzhS9MgMcLMeVh7pcJq2EVobowmB/t8xhCyN1FajtdHO+ij/0TpAj
Fx6FUUIdQs/Beg6LrhLd+IdLalBgfZaujlSIajlCEc8ZRhQ5Fq8XXL0UvpnvxObuvuEmKQNTHExw
eQR0ZJl7YYZHoLQMEPBRvepifDfs5QsdBeLOOyIFP9Z4/wlwNWR3LHfts2Tm/xv70SjJ0aZ6xeac
wwSIbMUF8Y0nEgb/RWcC2G+KT+wrQCErEadtMEBXe9qJTRREAcgjIMhUAvXXWJEsogDRKPxunxuI
Rkxs0p3jCuFy9MEzKoHLA/W2NDzxyk+PwmSrKfxyEshMNCQ2EJzfoUtGiO2XxtsKcTKxyWq4hJPI
ZA8cbnLf8+iZgoDi9PzIh4Tk392dCdt5Ecr2sH5NdC0ILkCmlacfc55nXCFknYheBG/Bq2BC2OS4
gbGOfxkXxYAd8YOWVq7yO1oFoH3L+wUZ4mNlulKNgGQUJSEd7UhMjRuCzBXxsFabsgDpPGjyivyS
dwfpRju5ey1ThTQcZ1Evru+phtnZSpmiY+AaF2AXEcZ6iV/R5Lcehnh7/i7i2gXR8nanlGc/i/Cs
ej/Gd/usdj+yncTD1jpBsW4qIHzX0ZyW6YgYO+aC1YU8oWD/Ka90LSGOjX7OK/zUXgl/54OlTy4D
8je6vbt0Kr+lemXBL9clPI4TNY2PWxiO2z5Ex/+S5Rs30S6nu5Y7R/Bu31oxH67pnL7DZfQcR0Mk
5Z3IH7XnH293+oQJIGoewFcn6lpF5jxzSSxfV2X/JRoyhnwBXZzltNo+J1BBYAKadttCHRQAqXv1
5vDuyqyEEeT22m+MrF7F8Y0Vll+ZmAcr0/tO3N0WUEd9H0tHNB1wSjAstu5tSFPnffFDmGn4pC9u
oVujs9o5547wkrRD121ta5Im91yIPUIHIyh3HEI0OOHuQ5im3f/fVHtSmhIuiXzWJyvRECV1QQ4B
/euRTNjRrZcbMFcpUTcubFav8udpVNpZzMeDCkB/+z9PlsVTCVLpCjh8fppStzCdjOgPrswlgdht
XXccO++VTiqB7a7UTAl5wN/PCMiHJUdSuK/Y4C3XqAL23E61zRaAQURgDJoW55xtBVQU26M3fPFj
hTSH6q0ilzhd68CjlbIAndMIyz8q+WCdsbOGbhv2vjNO73TxIuqpGc3tWulppWL9UwG4kXbMCC4W
wIvYyIlkLQvVyho0hOX36QWEa047pKWIGCk9XujsTt4Ifl99rxQOwKNJo4yvXwZv8UUqZOyYN41d
GZC9A1FRWeROktBX+IFQf+th7FJGLQ+JPAvLMELyMeFcCEO2EIQohFBZBlmktKvdN2kiWBxSAwiG
xFCFGEFOF2rTeIc6xeBboT2YjVatRwvvjfY8zDFjwj7puqhLk76+25Xaz1exZQ/W73gnVotQy0/L
yUDWmL2COw4+yV1EMsyuNpcjqy3oZ0JcKrmMR2pbAg83ODGliM8eAWYLS8zFp4uSuoMB/q94vVaO
4DEheZdXDdXhU30EF+2fdhoR41/a8g82vJIQT++d7aEWeuyupNdUPeHoK9Eca2Y1s9FEWxziS15m
OfoBk5d5Ms+qomBY7ltHNdzpCCU2Ev8YIoQTA1Kq90k+x+BjJ9z/9J9rJVFmmRRl40rWpjkueRFY
RkWXts+fJ6VM/ZjGDBY0iDKhUcQ1uEbae/EK2W3QvN1hkQZF3qj+baY8B2LWlhRKdc2sS0JFaIkc
HLAoyHnJpAsRG1nvfJ5dCemhl0yGx0+nrJh5nFDtGkp9aUPNeSFuFltrjJOgYxUCCQ6+EtiQ2Gx2
Je809N4uHLs63DW2kX1RjMV8sjU/sFNr0oxhM/eEWUYq4sKajFz7gCyn5DQSGi3fDj4vOOZx73T7
+bSnxUY6Jq/AhPaZTwS+bFBi4Hg+hWwjVZ0j6UjoUFfejKp1yP27EpWXBWh6VY5bNkqr44csw2yG
5Wp5Mq+mK8eamHHTfMzIWfGcevI7at+qcoNm8GIRlfAW3z5bmOLrHHsrXaISesbHTQ+8tSCoYgVf
r256D0XTEvRuRDzy72qIfJc3KmXFL4TimVCyOoEMu3a4qmhNWKsmCzDehfExMARsFFxx0W/Vlqdd
RG7NnBNDKr8kuhcmN2cDWfUIUNSuI3Tmbb+iqeZ4GluigBWOZTcNeAMcVmHtiLck4wC+l58oMbXn
SWqliiM9senfRQcUBraGnH3DsjGvawvvEEQQVCMrAGSyuivebp6u0bjqlNKLaQBvOd/iv2/4bmDv
4eINBesSmnmKI1Qt6u75EunXh5vsS14ZK02/NR34uf9zA40//Mdbs5hY0rhAAPdnGeshTD4m4Tw3
J4XpR/OS3Ds6mp++iPTmUysf5iG/MPCYahznTz6BcLoVqg1gBsyqKOfLw+YPEAT3JWdhPK8wb1r2
1NmffqBQnwexuBCW7gSZ0hkUxJjsB+JlM1YipTaNrRsAYWTmO7rUiUV3KJFWKgxOF0lies2VnOMa
rXDeg7Z/ebIqICESN90BcqmDnA31/fR0+DAeyYkhP8eXKXHppiBao0HWYQSCJzkbe5XBCuBhJbBJ
wLVQdKd3Mfako7RBgdq53mFQJsVwhk3Wv4rUyd9NaLfuhAu5Oh+KD6gMHU7pwOe9pfDNPEJUe9zH
GkG6sH4IQ7keacMM1n615q6ry1J5aOIWoI+HwoBKYyjufyOfOGhgM6N913mQ+qp3VdcI7Sk01BfR
8OaSRpep9Xq0K5X4dsUBEsdZGdPRCxHBJvMYc4lDxLwW6O96xbybqJta6pLUtT9zKtIGsaKnPjPA
8HV3KPxt8L2VfsG3edXEPQH3/52YGVl4+JorUx3crKhAUqfaLHhllhyGKJQERQA+C/YdaedLsM/x
Gj+6SflG3+DKdTPkSVhntI9MZMwu2yznNT8lHfuIn/RcJrCUA/D9fnuEH9DT0U0mn+dw2bwZlu4Q
G8fenRvlvXZ02U3xlWr8BjPI/KYX892cfHwLRkVgpY2qZ39hdoMlwjedVx3xi6gLl3OtgxAKClz1
zj6aGy9x7dPFWaQqMgxOi9Mw6AYR08aDpwlwJuY6M31lmLQTwRUy8XOJHTuMQmiisThTKqOPtiLo
5cc2bmYo0Zdua8HTBl7d1UEDwZeWeqMof3MFO9HjWUa5oU7+AAXLJqRGcrUvnJXlxF94T0b4S4Y6
EuPuzqbHKFSR/muaiSDTiwABORWOm2oThYP2lnVOGwvijkZOAzJR8HipXXofgufl3V57sEGkPv+S
YblepBYt7B5szi36kpq3oPkYuqRwnLI0le78PtEUhva5VSoKO68FXzWgYFb8JcP4yc+koZpPVqp0
NrBhmCHLj9iMMo7DUpuUfON6mqZLCwX34kZUXQ4EpN5jQ1phjc6WM1VVVj72bvd834F8j8e3Nv5W
VUGcJXGE1UU2fP/0046G/DsefFOHIgwhIb7kGRcbq1V8iasVwTfixXmQhm8heH2kMeOj8+vn91jt
XV9ya879W872SM/SEgw+Sw1xEk33bfdXh/pDSg/bmMDoEK9xFu6p7fCdlWfxUyWe37Xic3zRBdk1
TuSxdlKBSBV7Z5imZqCbMjhfCPWuvF/bPHc2eK/KLPVFJkvPgr36UN8VYIOdcIHz14ODXgW2cSDX
6/FC2Je9oTPCeFID2qUqllLs8cOm/ra587wGkBaRfB+LwhZPE5OGTN42wQuJdUfOilONr6GWeKgg
BWy67+uugmzmui8VnI7UWrRNjWVTesHomTPE3JU7fdRHGp+c3tDCe/W7/FO4yed6SYqqK+HaEaCz
4641bCA2Cbwl/SH2CbmFcMQGhCUr2SgPKGlRwPtT99X7RBc9Uq7R1nPlBQsUES+i06uViDr5m0y5
owY6uL/mmVDCgmVtJ6D7y6Hs0wkfH0sVq8t87od38YfbDG3OfCte7hX/LR26I2egCu/ZxX28zFU5
upfdeyVIXnKoO3X/48Zo79RcVepyfTJCoQdMTvNFkIKmY2TgEXoDSkL0Ly1K+/VUkT0L/oxTKsEp
Wwbazlb274NxRjvdkipKbEGb62HiwHsctj0JIAhIWXDyAE/T56Jc3WzkScFN24b0H1eBaVjSBVbQ
Cbc9rRAnz3HOL5ZhqHXqFWbsrUYbOnXr0W3WAqFPsLfox35nDXc1o0Y+XMPNRpc1B/68nffYNRb/
VI7tPBAkXokokHca1AcrHpmwnCDzjt1MAmX0BGu7QxcGgse1JqopWwXIojwO6DUZB1jENpMV96H9
2d60fn2r3BVmt55Y1dQEIIgtjikT4xHHF+4ta72eQ0eBSxtNHdbl83S3DvFc9QShLKrUBOYvFnVR
Nzew9CdbTM1Rqs/rxkCSw974OhXLogIteDOTeUknKyYN0DYPr7JqjjLLvZ1p54hvSDPZZxThydYB
VXKiIgwKnLP6ztE5gpTz/npEtdWvVlTorAvVyCl/n7Xk3ZjsNcJUD1quiz1GwNzyEWVBc5jgwh3i
2UvAwvXoBq1MHpsw6KxKwcin0+ragBGHn5ITis36RuiN6NRG9LpWjhDeQzs2UiKufBdmBcF+fWEV
xae6KmqlXt7LjNVIO+OLXCct2msbFD58K1Yzm+AjDNSvK35rZ+wsulC7rayFRpP9fLIMRMaTg0Bs
kfIOc4UjcUd3nWzAPicKWG9qCYwIXw7c9UAbiyQP/+7MjJ+uabTKLG4r5TgPRoB+VOe7QI9U/Bcb
qrFQ2hJ+K/OI66wprbnarCiGDH2jMZAT6kwxQ+9/bT5EHP7lyO72phVpSWLJL8K2dxGBPH3kIt36
TdLMjBK34Udl/jAripcvXwC2aa0x0hKd5eP5tpMFp1TKLnb2AIGYMCSKTdbMFVwLEyPRRQeG5XFE
KjmZMn41WliAfuzP5QJ503fs1vW9oWEsvrxYjSNxIPVJqL8iaiNdSkGjnkh6ncWzCsKdhl4LAmKE
2X4rzqOjn/eXMepiYoz87u4sGKVCRF8hw7DMCVk3R9Af7M7Rc/+t0uh4AYzZ9aexmnvP7hAhWKwD
HB7gpM8WjzooIqb568WfBhEo6S8ipaMhDElnmIcOrjtvEp4x/GEOw8aNElee0wNI2HKWsgXV0ofV
firapQkQNIItWWnd7PnsNewiQWvRfUMEG/QUMzw5iksQDrIgpoqUMlxgF7igsas6+kaduqjN18l6
tDCqqx729ubVulvzP+1RDsMZtVRKoHwFzY+GTpZRnL/ooSwCEjIfcA6lVwaMZ+EGQiI2qa+7uLpt
JPV/ntwHju+NqhdIzTTsTBR1XeXEqmQ8HKs+sd0aeu5r9GB6X+pG5WHNS3F6wL6PXAsfsLNb4Ldb
BAcU/ZVkz2yKZxzROrH40ixVa2eNg8IgkO+h8rRIQBbhrfpJ4j5DVHXl95iFNmUZcSKYTKwMpSfJ
JTK3wHf4pHYF90aPbX8YO7PNFy7rST0mKUdEhFwV6RpeqI0uBzOk8ytua709MkEPyEBz6hAiwPN0
+55jyQM4Py0IvD0RqQMGC8dDgfBkVi0AzsvplebXdpuk6ZW16CIJah5jYqYxmgfpgbBYIDv7zmI3
QSVbM8PyUHkpiOCR4ubs9gpmo7ns05Y6lHi/uGs35CSl+J1zYFcowRDMPWxZYEC/PlsDWIP6ZL/E
/XtKd8Gr9hApezB7MFoB8MlVp0LGgMZiHAb4db9HohbZI62D8nwBV5hNj6mcdcRxTuKti8LhxENT
AkXQhkAZV3v7NSMC5fjFj5Ov4/XdWwrgonrSdtY8RjcW/4AsckLTu6f31JMl8CJV2iY3WJj1n/ae
qaPBqeIEtoFPmr1BurjcludvYUJlEMLuag7TpXY+yOaZS9ShKogehhnP0svCUuN/NQqet/dHBy0d
nYI5aH86+5Th7+xI+2Y8UsDfO2s16i9iahSPb+4sJsyumTOXsQks4FkEdeAC6wuVVVCxPSB436RY
cEj4/UZnOQVLSA5BxRX2/BPnMAZmHNDoidWyt9XgsQfpyLTvdRaTqbiUO7RFZ6J30B1YPryB+YJD
wN0hdgKN0ZLC2gXjvmXlChe73bvASkGOEZmMZXUQ+X7/vV+HRmvrOmHGwLHuXGiWjW8idNaDOokE
nhXP9QbfJWb1zDLZoQHTOJ7ELK9gTb5b9d79Taj9wGtTu1dlExAG08L1hk746DWuXTfPMeJQCUpL
3AOsTehzKGXUGMR7kWOc2V2a7PhC1HIMOlPiCP1MHBy4ppCpPZonMSj+bGxP3iihnYy/0CfyzDUj
q0t5Huy8vSt7WixuhyQN4XIotqrhfM3TvOfbuFdZbsrnwzdMWVRhFnloTTogWKB5uuxg7tIjrVpG
Dbzho8rDKJZ3O7icgOvrJXYQTI8JmmRrInc3lSrzqGKZT6hkbRAU6SWAEGMlSfoHL//MXy9TH0Kr
qvP8fpr55unOgeqdowuaS4okA/JHHW3Oz+7zhRxzLLPJFTzZRbSIjhENeEWE8wDzmTvgY7WaYUdI
ZRBL76+Absbe2Kfxz996YGa6mWMAS8lUtTiqcjkRYQpjbxBCLGNjjeyjBw0InlCL0uZGEob6md9E
XdAZTvkHK6iziPD5jJXXPadgaJD9Nngpk0eaHWH9aLfoYTPa2vyw4VUZLGRmozcBhQM65swqDbty
xyiWn0YhJuCagjn64EpouvpIUarkTe+KtMvUzG7ZfHwpVg6uIAFAaRl5Fjj8eei7CmxhfecS3M5w
fPtQpSqPylqD6G0ZWXwAf1tf+zFbJ4dmv/9oXbwIPan156dMwDEQuZxY13UYXrSNiiUFnw3OUJMO
QJqlr1gx7iy5ufy/Sk5d8HYomWY40RYGSNBJMsJSQ1gSPPSZsK59XLguMFGV10TGYn3hgcUnGIaa
+d4MTRcnoDpxban9gm3bzbvWj0IVeOzYDpXXMJJ6f/EKiPpexEOGRxubJBnR40J14r9mQAOPyA4Q
sf3h1upMhRDGjVA1FiuHwhyWrrJ03uFQp/0kNo7uy/CA/4QKbErGG13v0ZMG/dK4jFfyIp6M8dbC
KlKrD+Er3VGG3y1WwPWxZIT4TE0+DRXyWlhHzdZsft2GZA7dN78t5UD7cDdK/RDDCa26zaGRCsi9
wEHPqBpjEO5kWeKWHL9mx7aZb1CGtVv/CnjwT0COj5Xf5hbdk/Zoy/ujibD5FhJtihxLVIG2wPqF
66aJQ7ciu2UQDcvVlQmm8iDyYNFs7XSsJOe3yAS6digVtDIJ8CPsLasROSrSXI5Q1a71J5ri3Fyp
Ih0JwToquo66WP8E1rm4Xrf1oBpOc09Z19tLUJ8DZDPGVRIiqDkEC8yUDMu7taFfP4E0T/zgdrXj
Un3gUwj7Cad/y0tdy8stv7inMUGzBPj497qnlCSLTs/Wl9aXf2W5ZhGt98ET+1kK7YWD6uOxuyue
nx7vM0nbkd83wbk5wY/DBVG8t3ijb8QHIcwsmTzxkwTrMAqK3Kc1fFFEdlZtubrbcuifxZB22crf
c1kwzJqUkOe3aiCH2Vsmc9F5ZHpD4YeJoGSYf7gNWXasa/cBPLywz2TDs41wLw6L65giqdi/pbRi
jgOrmbhtOckqJptVHrmMkTR8cAMu+dkJM5dhRwiBpJD27Q5pvsMfJWQLZZj0NqL6NjDjyJJpF7YK
9fdT+2qgiCvDdUkiAHBdm7j9sbTq7q/5PSj9x+o98Iz3Gs4N87HMPKoWOW8S3oFy2wvsDN1Wu0KR
QQLm+O5IXWfpo53ac0LNYWtYqQFC0vUrvyLL1Uc5BrpADfw/o2oRPgHGYCIcwOPGmljcWc1un4iC
Vf4iEPBjb/fAhyCbKydrYK89H49YlnKEAgST2BbozbKcZ7RGdPTOfENyik3aafvo9QAZcrdUCVFx
ty350L8m456NWPAC09SzBNpN6OETw6fagPwvFo1YhkpuxVyCMXxxEWT3EajZJWtQeWS1oexVFtMU
L1le/9iWiKFjFCWrHdd6DzQxFZ5Qz2bOEOI2qLFrvGjXNq4xgjNWE8S4RsXacyERk8YguRT7ymno
XxJRbY3a07FsyVuqEygPQDJssQ4+Y6AKfxOsGAfzGlhbDscDqLvcSbTVFcysXRXJ+l/oE4UnJBvi
GBR1aFwj+K7cQSwixkA1U+1XC/BTBAl9hMifamZcHU4u17S2XDAVR8vEML2HT22eugmEwPXLi1Js
4zq721s/XBacjYiE0VU5vFKOrSj7KihIBnc2YIQmUE01nbK/NpE9JpyOR285rnStSlUVyDc7vDjV
gUiME48/T7VsyPwiS4PTv3CVJOIwSAtZ17IV73+ow3e+5hujNAVjNlCf/7N/829ErNE/Ks2ivinT
6A5k9GxgiMg1Itt4J8WjJYK/Xb0tIX6NxVNfiob39JcZb13pI3rEOYxR9tcIPkfPgUiW1rgjVJ07
Q+wXYxqN/B5goNg2Esy/V9NezvaQlGyfI/05nbpXL+M+IpsqzmKvHYGUVcFy40k6qSbOvvvY2PCb
ogJOJ2dwobTjE9zc9wCJJV9KM3SrNJ/FwPrm21WPZ2ZoIzOctEy8kOwv5mSMYpKlMpFHBND14HD7
wYvD3GnsiJqu1fM5qno+IoNAQ9uoY3ZpeuiUaIy+qbrt7MCOfcyB0MbjhfH6Cch4uGfmUf4q/7Kw
QTrC4pHJKwlk5IlYdZzKv6ZdItjcDbfHPYLv0fy7mDWg4EKHNHzpoFodaVzrRdGo6qaRAF9n9oA/
dfh2yJxBJftKOZ3Jz1scZmbLwkECserUQgOOVWOHb7K+L9oc8wxDP4ZicSEyGL9A5Kg2eUGBoV08
trfTp54z1Gn5vJp9UMaFJ+7XDnKSTPQKEbipCwAioYPhRTWhrzijpc3QQ6E2MgjwnbP8a0O9YXDM
GzdusEMZPK0QCBFDHdxykCDZZHrvoXwAhdFtQ77DUfw1kg6swMBeeDgD5D9DGF2OYXW7SBh3+9KQ
7/5tg0dp1Wi4h0t2gYYl2OTXR1Oi/Z25II6SUucZYliZmQZmfsDiJyJThv4mK9hIaia9KVgLWTEF
ZSNWXj1WbMGkesF5EC8V5p+16ccbH7dz4+x5DVIfr8jQ+RfJarZt1esWKiP2UxRioPZfV9tUINkt
byL9SeNBloy5ZEJn9+29QeXnNOIUmRKQ2EQ8gtnPtsG9fmvtj86Nyjxi7ZmsLLGY2QEKo9pKDlM3
qwYt3I1hYnS+gneP6Cd4AbIe1CAnELj/p+03G5xrXyWYDqU4aoDRnju33VGVHsgHJDaFVtqjbHb9
s/O6HriHN6UEPaRztjhnBi9cAqHXnt/Ggm4wxgY3pXeL3zX2ceVf7vR/wvl4PKsxjCE+D6mezHhM
5HkMRmBZuh3jgnhwJfZsAZ8FK3O1r7EqAkJf1fG/1KbyfF61Jgizls9RS7j/aUbEWrQJPWXZpZ9B
8jT55gJFGY556O4xtVx0ERyoq/7K5/YMrxcdyOPQWkY20zRbEMy3Os/pQJ5Dyoq/oBupzirdxJBr
ikU3MRE0BRmFsdqgTFDlwUQPoCD4w2R7Apk49rIWB7uKCCqmRqoMLVhsycIy5+U4m3PkQYsYz/h6
i0FPy2iJJ0vs7jw9KXFHS5I6oaZwWIA0m/KdHo1poVUZ5knn7DzlFH6Sf+AXgEAbEAq6hsJa+3bO
50+xhPgUe8jXY6OU7nQnAk3zNq+Q1ldE/wyrIrEVY/yf8LYYxbmnkmwdiCRXVNK8y9iYi+sIrjJe
bdWdwwd3fpH8g/eMJVU9QWSRxOwBdYFiKug6/930uNgtjqetuhgsWPZMuS9Km0lDXEjUYwPth+Qt
Deag0ufodk//VQPjhQUihHXwUJuGior2IhiZGg/q8EGEMzyjVGsFArfKBUd2pOGgEDR7AI5S6mLj
vqCXSpS3hBSAhgdIuaFJpJ8HIbGph9vpkTTqeRkxSMJdlE7335MVMp7Dcd6JGp1+PTm3++7k0ysF
YV7OxlQN2yrU2PMCIVDqmUDa7Vj2bSCBkpoE/vM8sErvBI7YZRyAbzvaADki9MlDYJ2mgHw0Znge
PYksKHSOzqvNZkPCWU3BZ38xlPLNKV55aVZ48lBeeP1fm5Ufb6L9jPxwNMV8UW5AK42epM0A/E40
wz0EqjzZiWNY/ESpmhq+RA9uQhCCWlmbwnJ4ylS4hcPQh2zIyvjBhKlM7TX17VjNtR3PoHa9RY+w
wYWimyaXvCgHxfVDijbqKsikSRo2xvezTSUU3bqcYm+jg58y/9O91p1tGPJLTNG8mWWnel85GzqO
JUByGVTOxnS6lU8q6WTUVY27AFSNtIatN1BA0gJD/7cdV5/qpmQ6evORMK4rSpSSB2v80C2pISV+
ltsr1PnehMRCjTH2NDSSQ4581pVowJZPHcBP4GFh/jfLRspRT0K5b7XGnCydYjTVGTd7gJ+f02O3
wDWiU0QjG9w9CLhKqgdJE1vwfbhZQYqpNDFIRgTPaJClwoS7GKpRwbd1/T0HGd2Na0UmhhnbSNv8
jjOA3Q9Sk3pjId1GgIJ56p6E5AFqfn7eBFO+y7qF97t2BjEWOvBQhZV+U6PnsJ/zoRaSnP/oRa21
NjlLGul7GR/uB5t5dTQOMPRnS81Da6O2W8U9mhkcsTOz+J4ovel8PRzHQi9PWkChyk/NilGTsXDb
I2ikQutk/hvfj5EX0cnuNeBf4STX8/n3on2NffJTeh4gMvb8lQPuvOuW5iVo+eB7fJdYa19nmwg8
JGZTflrtIGcONqidW37G3t8hujoVr7AHFBJaPNi86vsw1d8VjZOjHsrwDP/oxbhqTNIO4o5qnk9r
AOhJFQAs9OLrnYOtIwve6FJJV88oH7emSTLdtrr14xPWmkx8GQwi7J0sDf4BzXYrZFAdyj//Du2v
uC+jbqCeR01oD3v2Y3MzF0VPTGeBVM+iekovKQb8EeQKTJBcH/3XDkp27E9nZEqVz9AgxIJq3H8r
o3uY0cLTo+p+kGW+1Lf9S00ZPxYu2Eflxyl7JT/LCTEV9LQztSYBp6oR8rmFX8GuLxIleIoQNaEk
ZO1u/AoK63JaPhs/jKcFXESdBEuSZJJyrAI0CgxlKqIbOSbXVTdd8Z+vxOiPe2ZHyJhJiPXCeiJB
TItd3T/VDuSdlnuYRdN3aBwXbyHjw4UQ6lbSsNGbrYrom670O8e8LoU/V7TiQek8ShqN/SyihkX+
eSTQ5ZDjVCA27Kqha5eVd/n0M+7YfxiQjqcYvIZ88Q5bZqMw80GMrbaOXgzOzpPFQhi6Vrf6UdqH
jOn6ZAXksafi2wjRvzSCbJ2sgQuoA/++LfPbsIgpGa8kNf86SvdilrtP47BCpdYF65r8hFNJsmN0
prf3fXees/SZFVdYuznfhCirPMpBkZb3L9IKytQsyzkkuJENLZ5ixBgJfMMPWUgdipeVjKCuPn5/
0KGZQF83EVmv5gDg90/MsSLltphMH/i6toQbRp+6hLliZ4lt6DjWHIDSYZ0TBZW584p0g+DrXv+Q
gFnl2zowOb4Cquxx+mqEuClk78/gbqG23NKGBTFA0vi2eZypKsjPgLdT82QYhPVt3N3Vx/Al7qDa
yQfwBXesCzqUtiUVLiXUXTkAQyHIdDNfv+6ti7+ZrlNu64/7fykD2u0QBjpfqnlDMKtWHxj+TRUa
/ikJ57RQNlz8vA46Y9KhEaQYRdMu+usiaiDDpPuM6Ey5FMmzC8axDEMhC3H9ElwheGKoLGvWyutj
+cMTl6STSJPB1txP2mTnou/0TrnE/6TiXFW/jnItXEVQT/AgDdX/u/20Fie+GiW4/o3l1paavLE+
lbPBp5VVu/K5LehQKBN4VdIWTkbomoUROJmTx4O/cZQ9i8R9SzkhC0HGFuvNqMuqV3eGrs3Ina5p
DhpGnW45bVzvDC+pjORDrv2JKffZU87ZizSn2zub07KXEKSFO6+QjV3d13q4zWFxFtvsUkiiQrGC
iXejX30XB/yUij2pkHYpABO/3e++OwPdYquyMVFBPorBa7cAwAsj/bBtfu4vzJsi7WD8KA1vdpZs
0mOvrxEXsLOEY5xA3oVROHH1qb43DzEW7UwZW66xk/PuuMeZLwmma5M9wOE1Fne26vS/RsS1zhtX
IgVKzLfcu0fnXYE5PxGwvCUKCUHs54h22cbqGED/FHPSS1/sraPWKPpqLzJyaPTr1QgH+e3w7PAn
UGl78I81ppZsJgWlAa1VfENCn3AiQmcgxpYNXpB6Jx6yvgxq+tggeOzeqfBQVwBkLi2XxQIECROz
S4kBdMeSfP6O13OgmWJJ4bztqjNNAm1tWLrioe+94Q79/bewf+wJxqP8XW2FpVbk6cxRkfAoQO37
6prRdUQdLvgnRZB5xUG4o8xIOgED99pUrlpW6gHyyuqcdgiHmM+YN6Qqsh4pBEQ5vy9MhEh8T+mU
5Kex5DbEAKVGS+ulE4PrHTHMbUnj8P1xmKaZEmlnQ7lejqDV9CKt8Ba+AFFCm9h9by5EThXz6Xiv
7ok5XJbeB1pFbPuEiqEaWKV1OdUAregWFJB5RgWKTHAMxB6w5nwNWdGu2JQKMtIC5z6VMLo+tq78
w+OIlbaj/A+ii7gF8zeMAkMkHN1mspHe3kLiV+HcJsKC6z3J1OdlIIN9XhJe64adTjdgWHIH56/i
2fAXIFtwQiI7eEteghNh2JXtRrHeCClY+Qs+rNfMx0rr14u2tDapnhzUKRdAA6sRL9LRp2lFoBtO
wvJW49jVFIp7b6XIDDzrz3mYIT+EdI2xiuqqH3/HlWDlsRRoRrlOk0vQRlwOFj+lJHADTUZmd+Cq
6s+EUFajtqkW9jRGTHPw0yPVGuTPZJc+jr9dJ5FA32ujG/uM/tS3w9KtICx8Q7U78QHDMpFq+akg
2rsEL+uVP4pXKstfoMqO/SDgk1FVOZVbxy/XUBvsT56bWIRlTA2g4C5woBi+GxA9jMblAaQbXD4u
c42g60r6etpi0TPdBhzJeoGKKAdoVcPyZC6fZssemHSA7SG11rWi6zqKartpqk0g2LSy7/sR6Dry
tMrxgKj/182R0YVWmFv9PZbivIzR8jRSyfqd7GSZVGN4AHmNlH7KrO7/z96iRnc+mYJj3Sa+2GrV
xFlzQcUPviT+O5bXE/mO/KNPCl+JL5tEF0nuduWvrjlvjxqwJ513F4GN2JH7GyAbHNaIbjc6eD1a
GlvyHbcmSewghWXkqZfxlujyUVq8nmn66zitZ2mDx+zpv3pInlvlRE+Kx/NlQJQ6WHaNXUvDeWw+
h4i4cpzH8UOZGwIFEG8Wy1YSLYRqo4HTekBjg8AXtQbbMUK05y6AL3/I2EAt32p8EarF4Ph4E1vY
/TOvLiK7ICvArro6QyRRA17ag8AbXgih7whcGFxSKfhfQBXOnA1yS3F1qnDT08PboadfNZ79JIos
bX+5v1b6dBLA92cLlChiiEUVb0lhLSEdaUcPrevWjPpaACkA+z84p0cI8OUAhG0bXITFUB27Idog
pUSZrJXyb9GhNwVnect31GorXlsTyKg9azvL0de7ZnJlg3Y43dMgedEC7Tex5YK71aEq2JlxmjDz
wwtc4/Fd7kMW8VQrATSFWDcW+CTn4Od30mCEpMoXVAtClQdKFJgLIT8hLoGxFetKzEJsdrapvX/v
OAGPZ5+lq8TMw7uMP+4IZekFbcFIo989hUofoVGoJFhnnQ4r/7WCZGGXXdmyiDlV+LWaz5ujAYBS
mkFJmRGmZeXpa6MSWPJE7t6bD3chbqGDDnnxfDLULjHAtwZNPM1cAsSi/MOEsbhz8lzsYDFlSacS
qeymINnn+Q0vcGT9UeboK3q2FV8uTwvjwp3uvpAw3L1aZp1VwI7fPgw57U3qYsHj9EmOH7sEcFot
kRMWnyuwhnRbnmATrwbx2jE3YCzoh/hvLXTZ8pvrdsCbczYjuUQlIkEbLzZ7YvApD7cg8VnjVZ2R
DZWfjGHQyFrJ2cipRgCfrvTTN5CXaa07ZYLLer04rTLlt7weEZhXas3VNGivSbStyvnXX4fPO4VH
8EmmMgesrDyCQfFgjjnkfDoFfjwRvlSrMK3wvTMii+GyVURLe86MFBk99w/4NrpHhNmZ19TOt1k9
TsAjoXe0t72SBCkwAc8k8YDwUmB2eVY37SaaSPA0hwaDaOb/Uh/UJG0uEpa+cu/sFbH+Q9Jsnflq
m4w/SqqfEy1JVkwO8t+Rh8MhB98Uknol66YJB1RUdskGR8jdFk4aEONHcmSAZXmCMckaT44eTssa
Icx2RBYuFPuu3VBsSaFwqlsMZHXs4NFheZ7aT6cH5esCd7GazKuo9dFNCzjNhh1DXEw08NK/crjS
zkuRCWeI+G9rXuEAr1zuBOka1yJ8EtuyN8TgL9JoQqCQs51CX+Ll9Kj1fYZYx8NZIyeTqTxWwxrQ
juvBai/xZ+0Ep+vr4MeWCniL2TNYoHkPIh4GjzLlf3/uxHGhMRkBZI+YagcJ1jrsi5XLAEWfbr0f
5n8vaquwA1NIaknoVL6Vzjfm+UgPUNAElUGI1TQDfy2+KYuimY28M4LWVNVd51tsrdZXv2MnGW+A
Gecg1v9xxu4djDjKTeXErlIfoyNdS/60dXpLnHWG8H3akjwK0nD6zYZj3y/+ejKXQVITC2hVtCQo
DaVpuItMAHMktdJfo0/w47/HlUsuoD0BOoG7NVtSYS3cOzpun0yXXe8LXp8m4SOsazHZZUUWuQtO
mzbOP41L3dlaUs0j6En38MgbPYJ7cYRTd08DkESDl0z8jzfqod41xRpoj3ac1cEM3sM6SL75S9gp
ODDp8rLMlqqv0JgRaAbXRncRPc5ziAzHcQM+aPXKOPkkHHYuJe0g7QqoY45usVJpRUXzO2760Tdt
auTw9Oi/jIvSSrO5QUM426L0NmQW6H1B9G/y4sA5wah1i4sHjjg6A9zJt0pH/yC/jr0pyvZQ3sPJ
HGFJZrkdarAsbL/1RqbCHyy/mU+TC04u8uGKxkpX2R3Oxx46t1nteTuBMbBPgLHBa8Dm5MTMZGDO
zFVqTjo/BTNvqSVfhNI8tzZ6uOy34i3FetHrkpzUCpGsWXtphzLw8TsLnZ4gwtjE74eL7qtiXK3Y
r13Rvd6nf+W6k88jbzBVwm/mw0Ruah8YZmPpaohFtPoDMX0+zjXjKqLHg65hGKG1OfC6Ba5wGwo0
M8SssYJj0Z1851qvVQxq/zIeBk5Fpys96Ft4IAog+Y69KyJiQqbDGHZoBBS4tF5Tf+z3K5QS1MiL
nbiJCoYanC/WOvGftwnwRudoITdMNM1bheZlw8vW4p7z0JafO3HTc1L3axBTIAaTpiYYEqD7pcwz
gduJC/H/CPVaBOyqRWeawtlMQRIpn9GLyOUOKc7cW+5mmxDP0K+ttcNrPsRYdssEvRjqWJFm+p3s
XgKczVRMjeXkgh9X+7/GF8I+9sAgm5CObv5wCJWVHYVMk+68vK8dPnrwQRd8w6s+pkITDkiSFV/B
OZOMvI3QSo3oLCQ+SQ86NGPcUWjhqhuZIBsUmfaFDt/rn90pF3owMl05ifbT3TLBkn4XIWafvn3V
4Zzb+RMFqnCFnisfeS4nw46FSoxdGPKs24zENtHWzzREotactAyvEV509EBSAW36PY+JXN7wvnhq
utr1dsxSRflVEyeaL93tsqaYzJQunimCbbJZCJeicxgLX86EvLAlxVgsXtw7A7ScuNMNmXFqMgHs
LfqEtqonua+99aB9y9NvXs/NwxduJ8vXteMqTsjWD4I0qdqp3WwUq/yxlvYZOn2uMDTNDqluv0Ga
rjSHaQZQScsByjqgAm5+FC1wfTWbj8vVHr1dvmleOCTs335nYErPssKOxzh8kI60dlVbmmTGdFSI
zM9Nud36Xhu/2M+iZGxZ83q6ey0FGozfyj8DJxh4ZHIzLwCXIaoyp0SCIaFRuCTZvhIagc+j65rX
I9NRZCqpvtK64UVipij2AEGrQp11MVBNpsSqwr69Q9lv95DvLZKJlcjStiBtW+AsV9CRdk0x/XAU
jed/90KZr5OHqI7xlgNNGvyPoPDXFGFi0heKWqWWCooYaEfmohc0LEY5Tzptxl+N0AdEjEGebzp8
tpbOq2iF6b705zGjn7ZeyOW6TG9XujdhpGxL/qfoIqdvvlOBQkZJKLKnHamGM6gzcjUYH/lgprWV
8loNKmR3yP493n1muwgEcJy3dV0mMT8NHpsl9XSI1z696Mpuh8JsbOh+mv4t5tvg9aWqe1Kq/J7+
m8hXolE71a0BVvumxWIk2v32OWcRcAWoPMACG37UqoPjOu89cTEi8JJdK82hXJXydwtTpcPHAPtt
VmcCaBWmB67ofLoL2UiazVXpgUWehPyauRKPbxu/w0ZqDoZEqMoGkDnYoExbi8xF34jzWx+/ga8T
+GB7s5TWEnpkOPk4PEaTmZFWUNDsTO5e1QZphdnqXPOgcYL2lmw2779pP3axjXfq9u9gtOq7Sy+Y
XDoaVPiL4YpF9dskmBE5JTEHsOeXXHn7mdlje+4z3abGXOwgqOSvwCKatMNFv6Eu4VWkdNv46jJw
k5HOqFtRQvVY9024KENjIkIRyA3lUDEkHDsIL/V7Y4FOkh8MKb6mfT2ajIBqVVoh4tMuXgS2gqim
JUMRb5pVvafpdr0ncfYoCAWuM2C4+mMAQtjjB254cjYPVqD7i9IkTnYsHtGRdaFR0u39XRVLWGyg
V/h1fLQgnZb6TD03DH9ZJpWgQjOOZnVcKAAqhUb/L9YytrCLo6si3INxkaV5odtHQI2+iw0wU8JJ
/2I1VwdbCUGQVgGqUnnewNppM5kKKo63A9QEhuCKHDLfO1xISyF7t5U7ar6v3zSPDeEqk9GiMMBg
ZM+z4BEKK6rxMmiQ95jIRjaZPl8ZD2VSG+gX1aV3u6KMdd6AnohT+LWWuSG/odVchDebPU9gv3uu
OLd7xiloMUHOUObfPDSMd8QnnsXeLb3sLpFOTRbu5cnABBqTsDIjE+gSobnUUiu1DzqlAP3XGbYA
A0iWphpU2eUGDo85qRntooCbe84r4WfEtWDyQGR4vkijdUbi2dz3qWJMAxjPo9k/Ndz7ibj/LxfW
N2eIpq0m9FESRU4n+Hf8F0qaWfXX58YWbixwqY4bJxU4/SE6EggkN9RPLK81f9N4mY8wIkfMaIv1
Ym/wctQJ8o2TstwO794WEDU5RAPHKsB8wcyWDmkrbjlPETTwMEUhZRhzGtY4My6vYYpxedGlwjgM
FZpN3+GpJPXsnracl9HowFL9VTuaRz0VRy6ZZ4T+lkj4J5JAfgRdukTemlkCsXC0ctTaNPm3N0su
w7LL2HqLqnaQtnJ9YUi6cYqRXs4DlT6r/pd9zZg2vT7ZU4+aiA2KiXPdK0EjQf/rkSf/cfVCxdvU
zveXr7r+XKunuFaQr6NnODeAxyGv6RO9Q20imWKomx6oiL68aS3LW8PIoM3j9OWZWEFqOVdnaL3U
msdKIeXn8FiV8MhoeIyy3WCiENWXMnaRNI2KXPY9ICSxcbv0YfcCQxGRUTBmpLZVrnjQhD4fPUZo
81vGJ0h0okxqIUG4b37nf71hylHCr+1XfEzsAt5lom+NlQi3TkXkYDV862PeKZ38FmfcHqSkxz1F
7pqg0lkqjVpqbLivZM98Sgkt6MQBdDltLgTlVZ3RRMa4AVS3SgrD99jZrbu0kHNfuuo2hLof2Wt8
02cE2/LH9Rp4mbTujYxI+7dBcVOqzqmwSDB0fgM3SJuAbwGOoRj1pAYzTCW25+6CK/rY5z8qFlF2
Xm8rOT/cMzc2M4ICSLPluxsrSgsj70yHLiRnmTrOVwJmsJYRpZwS9tjs8fxbuZgWsBWKKjLBN7Rl
AgjIpZ/EJVTz0sULwBuXcCodYonrY2BOGNzHf/ZWNtTDsxn0H7bg30oIBFUvzaskmRmd7PIMimvI
TGEtSgHS31xyoV8fqLS4wQn20B/up6XLmM8PrOoH+bD221xdT4phqUOpc43Oriha6ko7vo2QsZqd
CZ0Qt/4p0fIyyLK0JAKJO99wGAhb7+aOOZ7qxojTQVmYEljHUB8rL4VD9pjv4Fzrow6WfxE0OG2V
j06Mo7XXtEgwSH0JjZctcJcagKsXTywbfmqiJEVAqDH/LOPZmgKyhzpWP5AvW7uJCLPbtoCQ0zXP
kLEK9tawTRu+r9blk1uN8Wbtxj6hwbiCdtRV2/N7aZHjP/iZBb+D7HU5BmPx1hVzCc7VQQBKtu4T
zvj38EOvv4NurP3h+yrBYN9nuD0nlWRpKx38qY39xcZJ/MXXvnNKXodBYOLqC7oiuaBgLC5iMkGS
gVsICCe+G1craloggAMDG/Y5oB9uPz/+r/nEOcTE9VC7HVFRX+/taTrmsLo7CoIr6U+BUdOVXTlp
fdzIBink7wed73JyAp6kcWh19Yg1o30mHuxM/82ONZT05rqEtgQwCp2G2H5JnOuW1AiNLHflHgNl
390zJaak3e8sZNVMuiAApQh+IiWQTm2906dpZM/+ze4SBMhxXE75EAAdhUEzhEWTMfB7utJM2lR7
FOi4nOMyRZrdpaTcR7i+8TxUy3XaufErmb67Y9qVcS96Guz3VGuf4dnucVPaZhjx1R0wWK78jn9f
D2JShdAcWZlbzXGpyFe4qSh69P49ReaR9E93r9HoHCc94jIk3hABQvae2ykIqEM0Zs0YGBFUjgEH
ecNc3TDyN4X6OLcC/k1Q0i71EcBbckxeh6wszOZ7XTXqtXt6wGJoGM5daH41ry+G26YFXp0qYhLh
YeB/jFzhohSWlRnq6piEqGvuDUlxTiaj4qc+uIOSP3RE+RojTT2tZ0PPCbms+fe4mU1EGuefpuTK
aVBUAHrE+pU8exII48AaTz9kDz58CV+D9yBgD/xSMQ+jEb3mXnQmVNSMjfCgN4mFSR9trcmg6tbg
zk/7zPIxMEc5DMC0F2eq/UM6Fiicz0DktLDKO/l6PcTLg5rNNimZIiLHouTRLJ18CxPs1UCnJEma
WDsHVhJXgXfU8KCR+pD+qJsEXHDPaRCPom/OXohysgzH3dmhUzBDggFxzAHgGu2kAvX8ediHbwY7
KLP+GzzQO6B5783f+Hr5Ore010R9M4wz8VnE4li5+rUnOA2YJhmAA+1oTbdK20OJ6Sibf+bl8MfK
2PlrzbSSA5CgUzBwmKqydCC1snLmqmoUpdiFmPf3mGhjo7MfKJJbCH6y2V7QA1Y2TGzMeiQFQTsN
qeeKJsxkjFT0uL7su41/Ta94dsllq1298ExbDrM8k+Na8a7oWi0rM0UC3B3OkqczQwqv4++flrjQ
3XNH2A/4fpBGrLNTTmB4UuhZula2iYGSXCVSB2hkPqZNEbqG4VWSxiUOMMpaxE6No+OjjqPguU8c
QS2PucAEze/8fM52wYzYY1lj9ZuUw5ZiIsx9HBGhph0qVqF3rLitR5w6NGjqV/V5X5keA6rsc7d6
9WGfS9cdAnrzzMJ1lC1esA6YjlDy129kqSqsS/2/Z7rtSO9EirgND4iGo3CBREvQfXXtNL5a8LNO
CR95xu3vP6uMEaEBt+xHwEh/ptQB7jltIlf5Girr3zLzDwQgp1WRTN1EU/3wMfMU30ExxA+xEnxg
InABdZxePvm5fOiy0wvUcyeci8Xeksu1ZJEcSVnSRVMkdEA75qW0HCd/RLcFrYI/o1cH+6GcsPQp
8D9HpcZpLKiN652tZ+Y5loj5/ns/Gl4mz8OW0ZRAYG1NJJQe7pZAZouRDK3yAZfACmh6Es7QaMKg
CeeXA3vWNOGs2c2p+tzPoLEaNHBw1hlS48PYitTk3WYGUiZ4jrrZnnuYMchuwgzcGJfQ2DHp0ltu
x0Jh065UtamNjwVYMExG8U5AyhRjPmCloMh2aJ2aqdLomKjnbY6pibuH5V7NTVAQ2g8ENf5MXI+I
ooNU8EzNmlAV/4vGf+S4VLemaCp8ecnI4DfAa0c3XigeULacSWhVj/1rVXtkrFH72Ym+eSA4cr2J
t0d6XaAf9ZArfGcTSXbPDTwY6xz5nkevaFdfa5sN2pblSxkwRfMhp0FhVFk6tr6m0Rp0qXdh8fNp
BY5qSkt+KRV1pVOIv8H/fo0aFyJvz29/XH0fUzfUl1HTXGszQqh5WVaQYSPOwxx7wd7zIBEjE+PY
tSkHvBX+scZQpL7X8Ahv+9ffDdBooCT8vllDV0iUhipovyrH+SsmB5AzOc02afze8CSZ17XN/fUt
mQd4Msq9Lu9X6xE1zykJzU+oyzh8xVsBPjlZUj1VXax1h7qO6i1k+WiR4X5CoWLxibaxkYmlMBX+
sZF3oxHWCR/TTntXEiXDcbQVl+hLcn0FkxkfJLO18ObvzrnJdYncq3qKVFUJDZ0BxZpUrQPzsr0L
/UYVj3RqjbnxXrax4cbPweBI/fC9q/9G669Wgh2MhpyDFT74wpxYE+6azvonRqJj90kegNe6y21B
JeNIQexNwrLWMTbJSpXhj+S9h7pI5HnHRBvUK7W4wcgHJ++9odW5M/oBJrZ2gYz0+MhPWaojb6V1
BmSWoLzvCUB2k2Zp2+95alAYRYch+TeImaXx6re67PVQYaB46LkiHxHf4bSucZqfffMgP2zc7L5S
VeWYYbyAvG7rofF4apu2e2furiQwFW+HqeoX5B6bUP+a3Lwxd6bGBf9meHouKYFFBiahRfEDdml2
Izh5z3wjM0QpA3G6AmnJJRA2vsVlLcSXgjcoVhUrQF4A58CjyCsQdmf+W9BFLi0PCdZu1VAu5vNy
2aLZayNFIKRCg9FPp1aX6PqdvZRWP2SRLIIKzOLufM0sWjIvP5xBlSa3W8UGAZXhxh+39HAKk6Ks
oH769cser52MjojIunj+Xzj9/y5MQPBPcvBf48HcPsY0NQFaQ7elyu5r59atuqt0o2bHII/eax8S
io6kwzuglQ6TW1BQ+kgj4aCYKSLjZ3sY7nBCi3bDflLM8j68d0M9rLzqvsdImHKKqUWAuRlfoR6p
e8LBoseE5ClL8ciP9I3Lxpgr5p99RS+0jW3IdlaghBkMvwl9Jtg7s1zOPQqUfrf+J/3bO15hjFyU
TA++TJ1JqpOCEHytwRZYDvBzVqgZ/oV1Gd9eJLRot1dfurJtBGjkAitFCe5wNngdJ94dBFTiH/FZ
4pqStf44qnXWNKB+YQ5Zy0HCmxbjakqE8ivhSi55gyUSLdujWpXKRFWO744MTe0jrkj34Xir34n9
lmt5hghpzxWwoWwO8/L/VgYwt2DZQCodhIyVWYBCBWCz+O61m4dwtO18or91YTKw2Dt7UcnLrbuZ
2GHzmTCSRHRjQ9VNnILYqUgdfP3N7jWrHiLiqAOdHOf5a88SoqlYeLIekZUj7LaaqrXbuHtBhsTH
r4LTk6qf+LMMkTHKJSDLFe58Dxb5AAR44GdNsWfYY9QMzTkDxMxpFzhCNhPImxxbOX01ZkSgRwDB
F+NA6tuvHkR85+Z2eKLKnDVVTfXbUE0cEdkuMS1LMQQvly63QInMBk3ex7H7pC3Qw1+0/MK0Pv+x
dK/c985dzh8m/dTu+3mcWQOiECf6Dxw6cRFrMhmsJQQKPObd/VjiGT6NE7qnPJn/L20iGduSpzAV
nw4mWgyC93AOdblPh3v+83K3qIEK4nlzLbgdPINTos35YbkAXvMAbo9CGmpVuW6dZmSyxI1x/8v2
Qc45qwhp8Calk26xLg5UdatCEqP37ajripjF6gXiqbd5rmcQ4Irv6MQqTLdU1qblZsfnJsotaU6F
VvKH/Fhjj8WKTrMnLFOTozHLhPN9OqKz7UYd9zRnAPaT2zUkRL+YETH4exgTC16uNSaeUqM/iJnV
2aa3bZ/VkymwpkMfpEhVtCOgtvfW/rM5rAb5zi0KfSwXaa5luZkvWB8emCVquFeydePNGsPADzgH
smPRn0ydUzkGr3aJG4Pk/vCpN6SWiv96bshBWOUv1f1dRSIjQDrPR9/FvTsaVzA9dJmM83vOGEp7
2CR7qjfRxlq8UQEatOsKGhy4gR8IrvmMGmsLOO2qNb0xI+9BE0/7Wk3W7kdg/XoOybiaOHjxYOlM
CVSN6XRP6lt3iRHDK9bwGePehZDoG27HzraxXUTrpWJpFrmhuTskIAYNZ8JeplCmjWh70i6sApR4
aLE+xDfXAPfaaZXLSbK9HoUjbNCKIFBzBvJ7XrMw8jva82exJGjcX1jBhaUPdmALFoVPFgb8coW5
sTkGrmr4p5jV7hxVRY9BvId4goQmi6TiKHi5KCT/Scqpafk2aOUI9RkkElmwrc0atKJcqWK5g8dx
7wzLH8wbUwhpIM2jisL4vp7EyEXBdbyi9VS0CV66mF9QxdK/ggkeTKglII+QKq+cDQFOMDJS37d8
JKWlHU9D+IGi9UIS5bj3i9FcmBu59CaBmb5v4Yh/AJbEOGeHjdMLjH/+YklGQXng8suB8EbiDMoW
MeAMccQQQGJF+7z3G1S+yEdoumf2JyvolgaKAFzZDwKTeOYwNL35rJnlD1VPnKLiHG7K+4icQGAp
dgbuouiRX0u3qKtb8++8X1eGH5XcbSLG8PLxVO07w2e5BtwXYybCPs3eD6cvmLwD71HMvfx8dVa3
UYwaaTgo9yodtOfcGQG9y9BCPoYaOj4XFBnEqum7eYcldEUFQ7h53m78DPKPhhzte5dyejhcGjTY
6mi8Td372CYTIp5O7I0ZmtXgdvD5zV5xfbx5c49Cj53mmlbMhQydjgivEbQ/vvi11GBwrLjsFhkj
sem7L39hfz46fo07iRbCKQraVQflnGjhQ9XHjX8sp4Jizp9lCJxXb3paxfsNhQMSHKks3yBgiCSA
Som+rgmwL6jeY3ieHb7hXWWUtX9BFHTch/TJ88l7h3xNS+G9H7yzFaOQVF6WXjV5bZDnRbxnjXg3
OdAUBllMeyHp7h0Xr5Hn1fqSD07jnstlCB08XxOnbi5Z/32Fu+vhCe909R/YMgtWDYfm9MPyhblZ
ChP1gUy2RBYy1uegi2z0K7bbV3Wxu1Sh18B5/WbnjSKpL3JajtDCZAZAd5sLiv75iGwGaAa+U7jJ
KeoCw9GCQc8ZfftFucRbyFczrKxyn5vMsVmLv1OfbxP+E1T2ZI+nU8xj0Xp2BUXNZKIzLXpellps
GNpWutc1ZMOojoV+2hgu/B508YXU6luGkwztfJ2+ME93igNy0iq5xtKSFrnrSt9epgf/X9cFxF1M
GNQihuaF9P10GZOTdlptDL+kBib+WE335MGxQFdA2Zi0Vd4ep8Moh7BSiPiFGNT5pfE7+2cJY7rg
eQf3HQsA6bQhAi2fcx4wFTuCgWGqZxLCxuj4pNVqA/3akvCQe93K9oV9kVPdb8kygnqaN15hF5DA
U++qLY5a+gFGozM1iE9U3e6oavRBPLXdb8FjR4diIlQS2oNea6lYt+Swo06GDDKMYQM2rYfseanD
t84vusPUAmBqVkkm1Yci3VtzBvIXxlk8FlUDZDqu9HWPMw01iV45DXnmH6eS/rMKuum/WCCWgFEX
EdeOOVWh3TKNrQ2G8KE1AJJiOh7H7B7UvpxyJuR9p9+0nriF7Z/+Rlu1j6+Ji8aozML8tqJ15U1s
5/XGU3R96g2wGpa3oOQvwsltCJDLZTIwgYd5nZTsmLjoQKDE99VD7tXmtniMYWN5wtbkndX2YRf0
gkqMRVbh8RGjCLu6VySjg1G65v8zyz1vtkIIfIRvYRXvPst/H0dRBeRINoJwvsdtvU5UzuP92XB2
AzjvOhDvuioOtLkjx61e4ExZY8O1Xmn0ZEqaFHSFbF8PUwvC+sioY4AWlWnlHU9MjSKMtLbd7WlA
XTQ6mRSnCf/EbQfUSLQsd2mQRfGRM6lJJNjI5CkbMtfWd9Rcn/gH+glCxZdkLv1Wu4kbVU9YxwJB
UcEedgI94sdqtlOUjvfbKKrzlC+ieo0vqjAuWD/aIIZMqFghooQJwWMslZN3puD2JRg8uDmRSQ8V
SIuygc3Wf5KL4lUy7JBVlQgLkkWZLshFNrcSR2hsXFAweKACcLhlgDHW6B8Nc/NR2kKR48Za6zDg
D9IUUffkWc2gmT9iayt9PI39MZ6xIR4k0SFWJ5Tb3FGQ6898Yl1Ugu4I8mVxKpRuG+LIM1KZ3eXE
XaFL6AYMKGexo/qS62JtrmwOqCf3eNGFhgD/CN/Zt65kofbyWLVUYS6gV687Dgb3v8Txd0dBIobO
M4fvFMI0AHmH32hnJAxcSTnLJDgIjW6hVSm6F+w3zYDEwXnRnbizPoH44liPJp+LNbWch04mQ/d/
azpLgHlizBRePYmYhcHaC3Df5pLfjJ45Ny0oKD417vhZdq2PfjJVO8HNG01Di9D1Mk9GaiTqhuSb
AxDuNkQGHmWclbxFG2TGaNoB8BdAa5mEQgYhAfMIa6AHIYRDuyS8+Y/5ELqYkq8s3e+TaXMUaIq0
DMOL8v16coQXGVCzp81Bt7wi6MymHAYkNPxiESssh0zXMAlZKYZauUniDXE+xxrPZzKDOae+QOLw
fnZwtjSGc+dozCM6qNo3YbUYItB9Zw/B1DkB7zN0H2hRnLQFaBenFzPOhVZQdMyGBWK69XffMHd0
EL2okAvcPzIqaXP1EkbEPlzd5tisOJShL+W3kVByypXW7/8K/DLrATl4NdlVRcZRbAll8fHVOk/k
ZE9ZD9Jz5hfafVuzAWL4RPBrnXYJp2xQt7ntymArM5R0VH03vXbz+UZBGvvWkmDDkm35LLVh2vCA
Wc2F/1wadGt9EIpyCfSv4DYHUJ8rwwkiIuQwQsPs7lbNeu1FenM5k1yKfKaki6+jjfbq1zZMeg8V
dIYNrzSOH10rPZRezGUqdCNuKvs2/SmNFx6i7l9DLB/u47TlmCFfHZhGaBeMkebxQ9jUSEpfm6dV
oTmF16TpSyg2ki3fGiDyxmTwhCPo9g60NsF9XjwaF3DSdvrlwP7YHUC29Q1Ef0vIsclR2EXA1kER
OqxxTrtZVi9h10Jf1u7EDJMvG7rZEVbDO3HOeME6ReSFl2HpJ7XFthU/zDmddGE55n46Lwn/2w+4
uO7WXh1aYGEEnezV2zdZ3k1UvDTeIoYOmRHtjFfa7rI6GpQtZNk+1xE3ilGRj7wo9POdv/zeCBKv
qZ9AtMTbnRNFTnHvY1u4Rjk9tRHXjAQP+pVyPEXie1zI20lIhnuEgQFkHJUrkuTsx59HKehaHrNC
pi1vs2QMj/9V/Nb0ic3yTjuQ03IHyUMoH9Sn45rt8ewZ1/3v0+MotPP5Ok/2HK1qZhXpNLX0csEJ
4s638QZH9AalnNPj4UOXwLtotyRoIWZdOVz+HFYRqoW6RlyjOwMAYES6xGokmN7QNGPhiLfQ3/z+
NWHoRxkrH2EEuZvm3Jzj7OxGt6sPoRXImayP5SxebumfBT5gu/A8o6z+7NHumMCcer0U85VffHYA
YIeIgD9VDnssKs3cKU1PNrXE3LOpsMWrQ7zRh/GIJunkwUdM7Mc2j15QQeUWwNMPusjxiiaof23m
F4LJm4WFJjQWfhNxcFZcGup3ck1BtlhVJsqJ346M/q3tFwXMsv+1woeyXUX68IKNXeKSvBkeDWE+
AocGebG390p5K3qUmMavq7Yfv9LVYiDjLLfjcocuk72U94Z/sZR/O0hcuL+VkhdkHKd1s5OKt3CL
uRruHYnei0g+MZQHxVm9/zaTHE17z4zyXaEzbTRu1c2xYnrssT+74bJv6gqvKwyt9qtlW55LzKDX
ji7/B0NtGvKlZ3Ii2sn9zh572Or1sIWxGiqegunaZdLU5Y9hp+Z8uxS9wmp2sgIXxDIfsInKnPWa
mTwK3RxODg0qKHbWKWfTcu5FZ8S242ROnTCiDE3ag8swycTi0MI1y19IQTo+mROj1Lq9jsq8z0jU
7mPkayuTaJVPiy47zBjRbtZjzkdWa+idisjnOCm3+gDaXXjwkuGq0eh8TZhvt5bFH2CORUzzppzJ
w9B/Si0Fu5O8pKGAvfl8CuMJl+2h/H+6MAkEjcDcHaSvgf+mOxeUXxbWSuU+26Ic3UOkqMicPl/n
jJM97sNq2sujmunBwet/I0FZv/35Y2S4PecaNWJqA3n00/0RDRYJZ83TMwkDl/gDFSzlmIha6F/A
dEK2YxnvA7AVRyI7ylRbMHywPjJgtAI6ie99CkgPZTxUmKFqFxIjxWUUcYBil5yfZwDAmDZGrgUg
17U5rXTFHEXn/hFf0hUgwdPEOfM0bnFrZFTlk6poDXXIxslOcN5ZpcfvS1HAAROC00q6rL6aTZTZ
CyRjM3esen2Re1JMjQ2qkN4ww0NszNR/qpj2Vf9lPrSPqxIn1afjyKP91dH+oQSz0IRGjPQiN6W7
n6EbJIgIsIXCLyKUP9pcQeSuEIbxtMdAYxGPHmFluWXP0ffaeUw8juq5YTmKudxtLbNsUe6w9bzd
zscvEdL/FtltcfcvM0XmZu6ZSSsTnSvdCvxFeNasI64X0Tf1LBfA6dlSbqQeGMpLMFXkQIkjichW
ngksCpu7Qpu2J++w9cOYwu1Y1CPbpjZ3HXArrVWvBU72NcK/4f+MC2xZv0O5bNgLdWDbM146Jagk
+iUx7/7jbjKtIyi+EouyzPF6tbHZ90sLQbCTRBUW25M95ek37kZwMiU1YVPBmtS1OjL1DVizB0HR
wXoskht+4oC8/vsCb5u+gkxTwPRYh6MrzA9FBmNiOfDm2VhRS3Z7iwXRI9IkL7ORWzB5XQJw6npI
g0Xe+4zAqscZNqJpQGKbZBzp/JilsmL6aQvDGi59mU1InE+grgPyzf6ZQf+LiR35u0j6E8LW1BGv
PxSaqRiUntb2e5c1C7EhIgO1HGr1BvfrrP2ev73liKa7IsxnmHggVsxzLv9ppEdsZKoDLHm6p6op
8e7ltrFAJKnu9YMMw/J9at6xT9Ra7TN1OgqMlFDDsAr7Sr+Ph+kQ3NGgdkUWjgdh+jpDcfjDymc9
/QCGoBVZDfkoTtSwQsPfO4P17Lej5CPTUHiFQv58dm+x1DTSlSJsPjP2KEON7m37MdFTO27r5o+K
iWahvAWXoBPEHyU7NnQVttErDJ/bpucL8bxBxRsD6DOef4UBUBquihXRSDiMwHWbI+Osd9z0KHdS
ZU6dX5pXtME4lZpXlqD3WU5//OsYGYCz5LD73+N3oLouDc6N+aKRN9A55VhpLswyNhyl4fD7wZO3
oRkRxJFCZbFVM0Pr0D2mRZRuLHgzaPB8RfQ/rJZegOgYGhXjjIHTdtWBlbf+C9jEtiH/AG7Djzkx
waUXY87z0GPe7LxBJdRD0BpHzmY83E7puaaS5vOqqWMUQFPqHfcmb2IA+2j/zKF8EEPlix4NEk64
FWGvX6Hl+twzBwirvtOoYXpYnLm2Hbcc6jkZJ98wOkWljGBVly3PICXrREzAU67+wWl7gVFy2gKp
sydfEzoPuiGhjzNs1gJkkJtk9zba5q/P5zaFxTuW7DhZ0DVr3K+GTBh5ZbUjQOo9oHIXiLHgJWeA
4ivUJdU/LvAFI+0Eyd9h8pIhNGuoNPJrVwCepFszxDsHKEUp5UE2sywA9LZ+K5SNSMjP+F9lXzq8
XrazZZSs96vazXaYWscdNuTW/En4TOyFchxzLtWd4zKKVclfLhjQGfzq/K2KwZXvK3AG280KJ4b4
m5dRSevSXzLl6KicVA6idFW2uXKbAATty0YDp496IGfZyk+Wg7MyOCpu6+f3A7O5Eu2/ofxkREDU
aqx0ZbR2VAtXhCeenxYp+qUALd+J5nVR1IuyTOmu35+vesZc+P0NZML3RHjDGHAQLD9rQkGDj8ll
rcfmYUO8K2QWJ5myB2FUB5ZiwMn7J5kmFmYfiys1Gi5W69KOpCxCKgBmNEkkieNRZaCCHll04dOJ
Eii5Ef2tW/xNn8V0rjb+on0UZ4PW1sm/+k3t/hiHbVRkzeZcAa0I8eZ1Og0ZsKa23a2zbxkG9m7M
qrCdYnWbq1i0wKiaIoJ70/aT4yh35xq/JfatWpL7n6tqcGyKTW3tfVl+Zeg5L4DrB1Q5lquYj8bR
NhAZY4DnmuH9uYT6R2+psOS6ePXlZFa5mIoYOulaXMI9Cei74B6Z0FlVGlluqzLknBTRVQKdiAYt
rKfhR1LxAWPqMt+43c8xA7bSFoA2pmYXLG/kvS9D3Ru2oGr0DZPHYFhd9Y5LsALMlF4nnK3SY4BL
nRsyvRVUTYwWrJ7B/6k3VdYMVjZ4hPcvluk2QESQVNR7+IqhLx+K9WLSDBY89Sui/yx34ARxkS3a
EJIPnD7rSYb+EhqDWtR8+6RkokqGTRnLYZSLvkMjcwY50glZVm0i1WzYo6xB61ITH6lKsO0iNxRJ
oUEqr/q/l1d39x0U9Obil5u6+8riy7l3sL0XQRVkAo7H7UqQ3MYvslt8cLmi9Dp/u5yzfquIL8iI
a5iH3+ho0QtYPqJLY+70NoLJeU6kxuQoHQUQ4q8GfjfMR89COLe9cM5llxWQ7oiFAM4yh/1q2uOQ
ebZr2xl6ZcPVptUCI9rICtk21j3/6fR+M17+nM6cWGZO1gAQchXV92CL8okyqv/aoobsofL+qQaL
7V12erZgfcZKy6X8xsr4tXysQYS8S06Efl742lPYG1Pj6CtqsVwyaK2e8krX/tcGyNc4LLVzEhht
l6TW3bX9GMkNIWUsPzRwJ7BmOr/ZUU7AbxMiNftQKXqCKXJdyyZKAiKbki25MVl+uP+owruaJH01
WiUl8uJkPEgDiE4pmHLm4ro6WKN0LTdn6xDVtXqLjqcvPPIf/J3YdBTrXZyqpE5jVbNXbpiT2iCd
LaHSsiuVVLtuC3RB3wpSPSGhMIkw25jk8VA82oU/JZvpsyXoH3VvfygzgowtdSrgbuRAcijiuIoX
/uz/J64DAbqu5hBBjM2S2o32kCbm2/MlncutYVxX6xFEHMLaS29oegFNHwom7/UFi5r0NAp+CnPQ
o4puJ3dzpd/MncQ1+3XqtqZF8sjT3fNeuBFrCENPnpuPXIX+1PWV3kbSenXLfUWBUXyeLbNehYAT
r2AXrU4zHZYMIUBd4Lqt9c6Zw7b54p3g9wRxN3bitVydtIrET3Jp+FUQAXBKlGX9obKojQhE9hE+
MpIusxiAfkHJh0emJR81pq+PA3Tysf+BYnSS1W65KyBVOrSP5oZkLk9mQmFpCd1IzRs0WwPzbdg4
emNmV5wHe2xlwkM6XVruY50D9MwYHzc/v0vHdRlMBqrb2HlaaOmjDTf+XIjZaAMjjHkci0OJuJag
E0/TQCNa/j9kjogcmxyZj+Ue/Kfk1WlXGvvQ/R6s4Se5QMDuJsCv/5VW9d+cvbpLZfs8zlF7iiDw
dUEZufANeAb120iu2n+tOG6RXx+0f4JJPk5hRYT8eLNR6NdBZUF1vyxhuijeWnsuutmP4muAu3Fd
enOvm9/7cRE51ynRVgPaNzAG0Wchq2j5fHYRUw8dNLjvOtZkojjB+td8Y1Zuw3wx3/KRPenHouiN
RFmcT4/WgxZjOmZhONX63o1U9sT/2BUjImL6ly9f4yk71YrkPLi4lu6wwvGMgMkFfQwS4rEZ1iV5
qBCVqjHTK6/1eoWceH3vTIqCWa03Jz07CCpjvFbP8hL+t9RE/2NlIoou3pHxaHF130ve4CxneIk6
mDmOHoTt2yTIKQHRrqJ549SJkFHedPUX3mW3Hbg5VkXm0hGcyMs72JQuG0EUd108/DA9hGiu0PKw
Syec3752e6grRZaP90Kyckisg4rfknwkkLKgnjorAe/BTKABXdxcQgUp3+PSRQTWOcsVswcvrAoy
dgDuaDRPmue+Qq/oCdPzjD3W/rzswXDB2W+//dSFrBqTth5jodlyI0Lh5Kbsm6mv+AWocgP6fvML
PawNkiwnPnpV8BcP8YP8HE/QcuENN6APYXzmyrhAA4oT4p4ObNaF1B91QDAanQ5W7J414R1OYTXs
pQZiAIv64MpttGrjsr7q2Ly1SPGrvO3fbrAGzheoO/fp3jR4D/l1g5NYm1RdwHwzl2vEUVsxm4sU
jUohn2/wUopPm2eAlHx4aB365P8t6glY9re8Fjg5jpgkroU5MTZmhE9eobZR+SjnZSDWoImZ3UDM
n8zmq+U7joqeEGG6E5iqI2BQlGSinDZU+UMDcOLYC+pP880/KNxw5ht/wrx3lxnYQWjdy3nIZcSA
uOxheEVyjYdkJFbNrLRa1AZUlXT0zQsBSiLRT4Zt1hFUYJ1qaa7Kb5VMf3fF2NOldCLqwVgTEyO9
aFDDjtUv8B9IKSfQdQ6o+M/IohYHZf4994C2+MfpXa3GlvSy5ywnFvUa9nb+3nSpCyKs2347//6Q
Mee4WcpYLc14SLBpJLVginHapHbZ3gfWTEvdKfUCEDaifHZNjp9EyMx0+ddoFAD3EFz8ZF7cK/wd
bY2h+J6XBevxOimXTSi3muVoOIU+gAE8SQa4EDygo0RPVNIBQJNJc5JDjtOnQee05tBKCqtfMsDZ
MRk69ryNb0NhVThMja1EzzSdIWdowExyyd6SwRZUajOR+FrZW71dbgknPyIZRifaRoY4hWMH1PLe
1twCJM3KtpnmhdAx7bL3laBY00iQ2+O51DeczcpQZg+Q2heQsrILPzBxy/+pziWMd1Pk5Bc5bCx3
SrhvXyZCfrKEMGJrHFD4wOWP++Vr9dWwjdhg3ImeioVdnove6OUikAYgvJTal8sAQyq4orczdwsK
n8q784MdN7N9eYl4i1TKEntsbHg8GquN9o1Zj9157p8NAFpgG3CAFlItD23S6OjR/m0PG6v1oKkG
5JnFWJyAbtEczxnx1bbYodezVUrnY3uFv+XlVf8fZxz0nWIuaYuFyVl79bahBuUKDHuK9gt3Hrv3
ANKYm1Gn8vBsNaX+7LpVU4/GYeASMOpQOm7u5KKVRpJxuDbURayVwKf5iOovNrRscAzVpCrmmM9W
L3LBJnvuA3GgXz/NxnWh+niP9P1/Mt0K/Gs4R2AY8KnGJ3fioEEyadBzc9KC4yTX1a1Ws9AP/ghh
66QpfCVmJ7AOY4himo7xSn+YaMsCt9YPPZrxwNNJSAPBquGF+rGM6lX7Idwt1KIvmrmBpCOkapzJ
duOkRiRfRs1zolg1BGICbdKRC8FuDaCrB7DTMrBvQRjRtpJEFmKbpnvDElD8p2AoTIUCc6W8UoP0
5TOvaVLx7f/kKvUSLTfa1rmbcYZTf9oaYFBrMn6oJosnM3s/D2cb1Ob1rewkaRkNPTgBuRT21XjB
xHhsRteIiem6H2GX1y3eXMJdD5BKEhV8vrvLPC7M5sLrMkoOq1nqygP5qpwMHs/cPfa9qFpYgC7z
7ZLwm3UIz9x1NjmiAcGc8PBGhmcA1ThNpuB0wUBP3w90XOVxKS8UsiaZEMCz0iDSeSN4wZlGBSfn
i/Wdfq/WHGfcv63YbH5vcxqq9XZyziYREC6u0UZHEERbGGSpTYeM1vWKBfP9Pk8jHJlYc4lNLLv1
Lf8Z+Xukln/p8DsCc8LBpbXWJVM48vISWnZrULrJM+Rd10S7S+aJ1rPnweC9AkwYmlA3W+UuNy+n
sXc7GJMzP5QfOs47AzZeMTvGGZPrsjhctqiiBsEIxOf7g2d2YULE3imjxZ5YTBFb+jOTz00ItuRs
xeoj/IQSeNPQvMC2QDYCBG0yoUXv/qGvEtwdDv8ITs8mYeZwJaHwPBx2SnNQXNkb99qgNUMvErPV
BNdRYeOP+2ow0Zfqdt4r+gzKEHaiTaUUpn4ic++TN35nRByLszIwe833JcUibnYA6CSq1xuQK6fm
5De73xju9VmmlgUbrcftZuzZT3fBm8p3KNJ5V9ThBIS69xPlObII2b1NK2btu2xFUJA1orj70Cty
wkchEbzn57pCt6ToFa6cjpKcBqT3pm5OwsM9evHMoC6e0C/FWHFqtao0XKrJrNfNW10qnYter4uE
rgUwspXct2W+qtj24u3RVddDNY1SFh+cq7dkExnTFR2mSokWPVr2qfOgYhHLvgaY8zK7DpfNn/M0
ry2IGuD7tUUfRp2UKrVENmzqWMpsqN86XumVPJCMwJfh+mNl86QYY6/RXdss0dWDvVKOiGYxSsLJ
h8mCzgsf+yHTwF3eiPwZ/qcuxeNkunORQOlxbRxKPrkVbHyROMFCKR1y/JiqY+rUeovc9+u+diGJ
FmXxu8+HoZ3M/yglkRUbXTOuef9bJdMX5oZK4G5bZaWCUl26Wb31pFt9+1I1yGcn8rWa84ilIf26
iBSmba0g0ZBqmNF0XnwXgvAAAhV7sUZAswBq4BLNJ+diItashoAhjsbEa71IVleUA5Ad1eVX6yXA
1Svcyw++WI6BQqvyF5uOzQrkJ0OygpBoA13IvcsiXhsJlsaODleWW8094tJu/AeiyHd5rp5ZkjgP
+OTW2DilScCD/V5MGaSHmh2OMHisC0dKZEDD1ORt/xjnscKHIj60Be/HlZmZ9bQo5i7yEq7SWznf
UcFQL+YgKHCnYXWvNGbHK+Yy6HVSdOKZHcqZlBc3dhp0W40/eSXxMX8FWKHaWnhwqwQDkzz9wYvt
M6iughtPipov3KTM0CynGpO4kpu0AizFmQRo4RSSe2SLiqaS5BHzCWdwQV9+DP5l7w4kWvYErlO5
XCroBnTS7e+c5TkPNKv0f1HX6Pl7AnrrNzkFwBKJx2W+R9fGCDHFmGivASbwyC2RhkBgBhdr5Ima
GWtADZwH07I0weOcpJj+/Qx22tNi5AncW5aHoSTUvohx5ribNO0oOPO7kUPdL55FfkYSGy6Z82Rn
GME4sbWa9ZjoxA5erxOEbasaPwU5SdEJuRdT/hlJ8Vfc8h+tFnuM00rOODcdZo7S22zyzF3wjmQ/
dc6QX3XrKE2qBk/OjvjK3566ZajpXg3Cr1ylf+WmU7vW+cWJsXHydRf8XX3WCcCtpWDzFKqFPLLx
+Y777OGnw5qnzqQOdgOfyOQpc7rdYPkIOfKfN9Bidkgul7HvRh9sQWN2D8qqSgY504+Vhw/vwKUg
lqTgoC7/F5QRUHL/vzMXUnHziY96gHeekIVSBDOrDqSVSEY0vM0DwjtKd9YrRy/k0vr3uDew58Fo
hnX1T1w0qZBO80yaa94krwBpObfUVsJFai9dZPT8Ct7DmncPf2nDzA5z1XYIcW72qqRYArSSnMB2
WBwQwRG2QUy372SLQ6UlQF165qy3goG4nyEO2zL5wqLsZzXsVMqxp8fqo8RzHZmPxM+rS9an634G
20SXWwaPjNbQ/CBCeiWThZax5p2RMhqlDz0lcKB55uxDdyIly919zA6ltclIZYH5ztrM8Zsm8mGM
bBNkpiZOULzVAAtqdY1FBjOSywUIuKXla8Bx5JcBv8IcJ1klsgQFtuAzV9IVrnYIJCzwEGaGJmPE
ozbgUfJQItbfuCkIqO+g8ZDYDa/tboIR0nWIcXasncktQEs4kLFApdamCw21cLMOytCfj2NaP2Ec
j4Znpp9Xz1n0MHK1Gw8LGxE2Bvv3rG1KDnBoLR5Byyu1bb6KJ8+9aBvvA9XGuxrMulxpvVVZhD7H
0RP27pj3RzyRawvl8QLcKmeYwsGHrUwT5hdYrIxBh1e8cwJJw3zTLBqdWaT1fBwcEsLGJx9Nsj08
rBd23/o8pvlrK5O1cQdsRS5Pw6yAG1F2UE8vf9d0yQyXoNWRsC3TjXEMtzkda2igWw2YIWM/E/6W
fmNWwSwdeKc8cwDrzb8Ek4enXr/J1YW5ql37Hfhh5fPMt/5KLY5rYJoIUsyzNGr+yraUdiTHQDkJ
tKgD9grrhuC779xR7EhetwG6ijUs35JoBMp6kXFfIqkJlE5pz9vMYgqcqC4oht+XdnD067LL2cvU
dHzXcw7DuGGczMHhKnTQMsQJqOuEN2Xuto17dRnvAbpw6b3K5XYEYhj2QH741tyjGfNyLIqnS0Ak
1Li4SDF5BbiM/NrsVpABhiVrsRTQ8IlF/dIsMCG+ADuXnG+d4gtzHqYaiJNeLWoNiLyN9W2hyQEA
ZbxstKlz/bXeM5Jgyef6xQIQ12vsl7/xrUeCTFGMllGawA9mqnXs+HwI6xJORaFewZza7ZX2Nk5O
FDwTCzYJqT+Q1mAKNK7CSV44d2YgFxurtDzFdgdqD/DccTnj6H3oJVjccDcmNihAdLMfgLF9dobv
PjmO05ebVGo2GoVszFA8o3de0zysGMNewar36orgrH5Hzv6hfhlUInbpJYGhH/TEEd8th2HAl0j2
2qYmXCzbu+8YqcXcJn/S9w+UFIXECNz6XVzy/NwHYS0y6XB/6FiPrOte61AMkq+0XyCVLlBToTLS
Ks0jJMV6bEGw12WKVRE+0VlP23935c0zFU64eS1pt4oS4JvAyruwJQbdbbuZXTzCpGT0MVlFonA+
aU+WEAXiTFkxE4jj20n+PeymvB+RQiB3hxpFM11sDgkkN0frLSVQqkrSB9EF6djYQFK5Wdu/qy14
wPc2v6dSK+t4uAI/INOvNEwaShhcKr6EWBB1pe/UvfkcHMNPem5vPzVghsl+/ZWahBpral1RmuUO
4FpNBCEGytmsoyRx81AIuvECN6qAJOtRWfFrXdYd54VUiI/WsmXBBGGgAgHarla3XIUrLbMDb2lY
ZgTqfhxyqpFfUKrFmGpE0AqZhY+0oSho5xTOLc3d75f7T4JxRWrA/W39YXu4Vxg5YeZ8kUfg3wsn
loH1dk1EmjcPnCQtZr1akELz6LVpv9HbKAw82/egZUMLyB7ZHlDb6JZ791v1Pf0xTHrcrYqKrEcx
uLhAtkew14pycA7zBoADUegerT8Wp/nPrTjXKlghV6AkeEp4hIqRrcNEKiRoreUpDPykEIGeh5h2
FpUC7ghMiDQfRQIhzx1bvOqgXdgB8s+IMmwh3WqUeKbFsuuY8dwS6I+f0W+PRYrgzATZWerwKaDE
wCeNPXFdCNNJn9datkKYXRtAkQr7QxF4Gbs+uzfPOZwg8SIGc5aaGiWqsEHpfvQEogGeDzuSkHTJ
EgIFrCIIYz2PGMjA/3hvDoMpv0FMuFIGzvI18SB87GfpKRxK1ZH58UD6EC9imylovWrnn0kr8Wyz
UcvlLbyanams9VTXnEDfcHAXhKsFHPng+a3p3WGDkSm2yIyL6GmkMhiIDf8wdtSa1mBFKP2E7EFl
kRsKRzBg2ZJ3q0toFpXbE/RNzZKyKWnU9UY/i2B4E72XyU0hNc4fZXpmyBzXgY+ttUNFeNzekAYx
kSxAqsniuvF3X+A6+S0zDv1cw3ZP6fGVyAKXXJaf3XWd+RcisjH6oMbf4YXqXcvxtcwtTdkBO5DK
VV4BTN44TfNvd4aO7tPEDKTE0R9Pfvgl3a3HuK6JMQj+aI6lXqcMY+Ud35Bm7CXe4OtMYbp143uA
g22Y1zh6bLvS55wqYoQF3kpKLTaUbfDQYkdq94ArHgWKwbvxGg/FGXOHQH88UyDSRUkGRVj4a0O6
wndi5SDbjAKQZR0EHKf6X5Mx1glBTD9QzS/mgcu4yluzoSN5ztxjeS2gdzRefeesD4eB3869rW4G
215p+tDEnV8rpeKc1cDhREfrTjoukVt9R/uMkWdnkY9bTcH0dBEy/YZoV3ETFZpqOv7JVApu2tH5
z7+S9oDgrOjciVMV6v38ToYCuHqjTz1LfK3HP3zt0vZWzSU7Qy+Q2axDVMaaiCNUFxLbvSPKdGUK
MyH1KvkQ0T6ZnCa2i4fkDrUgK9SYLvUv7djbp9l880Zi4MemJGmD9W9u0GYm2yv7IWlVEP6YZ/nP
uAtYGBRfi384VxJLb/X/1vKyUkEIVddd20uwxE3313mKIkpEBQ4ReePXLd3S3qlvlUnpNXeZokhf
aW1OCegYX1YD3rkHfs+9heDWXgWlF8oaAvSz4SMQfReq6UW++QnDY5tivMG7be04OhC0XiBt07Ne
y3TBQW1uO+gxZJiMTD8IsB31lcwzaDYgUk4ILQDs2MQJFVfzCF1X4hmLEKfLJSN+0tlPntzyszj9
j3buLviP+RPFo4NIfn1qPwOrB6b/aUSt+Av7oEU8Af/VVkqWKI/9p6MF9Ak80iNu/8nnonnCCa4c
aCKPDomOogN/K81Fk55q90Ra2LtfWtkYV/L0alBnkQnRfebGbtE4+QiR32mTCi83Uj+uiF3b5qHt
nQqd6cHhUA7Wk1OBCQ7UFyTTxLcYwfCPmIngKfW/PuQ3yVI9OQbLpOLhJUvaNpEit2mmA6umVVY7
1tjoXNnX1C8+ciVK+u6PqPXMFNGpCjlNeXYTL15bv9tQesMInrnD8JakBpjRHi8kQxf2AuUeaoqN
c+dA/KmAZ6LPPSZJUJAzFwBiXRQMO4kCSg+uJGg+2xMzf3pub7+yJ4bsSi9LayTRF46QRzOZr/1O
UIM8cbNbB0A8vgPzgPXYCq12Nqzst2DMG6z5hwjWW5iqOnF0z43mrSp8X7+5PFo0pLu9zvvFkguW
IcUDEL38IGNfQWSaaBgk9kuMgC7lSZS2EZ7x92J6ppoqr10vkxZs4mBSyAoanixbeAqw0BlacC5S
evklfhNXD3YwugxvrIl7urMJkprny8HG0pED6bWqHpQQFOTaF0xCwtfsuVwH4Isa8tMaHpoudPrb
sbMxRFRslTAT9gE2ZnXlfF3QOjr2DOMvYRXuT/YPkoPqD1xDble2xgIqiM+T7tah2QtHez/R50+4
4t49cPq0l8Nkzfyb99s0Ls/Mm/dtDcLCddJEJqwW6SxQnj8sR2rCOO/S1b2iXY4RC21aAfDkalrA
I0kdiyNyzI6g9cmcd0Z7bxJ8Ede8+SpPivcQHSwK2ysnGB8hO2UyhUYu1u9v/IKj/igankfEDCvL
c/Nyb4ar72NwZ++5eLQk1tNq4zpYo8wRFs6H3JfUdkSbM7A2ZSXi8ZBDgNNxIAK40XpLkPMx1SP+
cwNVj7iEQbT2Aw/x/VaLDV39rEvPe3T2+u4VI90NesSg8qWNL8vH1KZOtGx1jn0NIyUx/Fi6mM/H
qWK9IIdq9tygZN5Xwu8cKZVrVNDH8MvhXsbPuA0nIiLfaxLoRM4KX+melUhcqBqAS7cV+x8BZBke
fwZX6cdCmInUYbyc+6FgOdjjCWXX00YIKOoyDnqV3IirXVU0lsQ3R6LSVnx0QN5+77IMzAEYLb6u
BpfkHyCNSvqHD1YeubPU7p24ppcK030pyK0w3bN1n99imzezLaTXnz4SW9Ud7xwIEMYwiDaSWy3P
DpV5eWROACWG5tXyu2khify6kCbL/yqmEGZQdngy57ZPSFLw+BEmQIUpiLndTaJC54G12SWP1Fif
t0M88B3jmapsk4Vs+LdG9cowTfKyboGl1y5MmuRCMsVQoySOXw+aIuuP08pf0ze+g6CSUr2xw8S6
di4rdehCfhLu/K3d+3ijBqIWKFtniVUiqcD6LOAzFB7odk1S1/F4rgPM8kYWb33Mn2WXg6CAmcxk
n+VLua7vy1/GqVxeV/mMiHIonj9R2GJtCAn0Fr6SLei5j58wstINcayMrhf/OWlzRmoB6Mlr748D
49SqsBv/RE2tQt5V7ObGpoOjNUaj7TlrPm9U7xn68tr6AHG21osQvIrCL82rn2AnbIH0Vd+r1T74
wBCe1jubwfH5Chlayt/QC2kPO35TUDlmQp19+uxoM3YG3FsDI0zblc7FVvU/t5eGyTgEYL+h98xb
3/jqJ3Q8SiJ4sBf+gOb+3iXxQcGXql4LOTgJrDhzRMm218HjDiCOvFfkyhndK0Nm9u5kN7Vc35jw
IXar3rriJbt36w82ZgatXfhLiteTPpXXQbMO0cpv5zxcVqIqQgYtC7rdR0lUPDMTpZcJtbvuk/i/
eWG3443yieSYvbwaBcMWI/P3ePCCl1sR/N56Xfo5tRynvVbsBj5BqdP9cOglikPiM9kCTiua7rgv
60gdWJdXXUKFc5oIh7olooZMfOlPLCLuHYyeYftKdQIH9BEqyHqu+xE2JV/b+PkV0d+Y2VRhR1F3
68zM1xOoF1nXO0sOIPG3T3dljpUO9p24SCsXJbFN+PiCZ8V0QOWYWhC3zeB4FkQOb/wYMPRSX5g0
hALXCY0xQptqFcKpCz+Uo89abvr0hBCGBXk77WztZ871NAuitaqKDoyOQUpXnb0o87dc+iFJ+o2n
9yv3D3agQkDREZuhUhUWBn3AoXTZkPAveBwcq26OUvOJB9k5qoRFdh+y9c0xRORlJrKpXfuPdai8
8EoVVgAQy7zLpp41JkmxT4shRcpC/pGg0fBitOHLDgKrRsf9HzD7vJHHTYK1TpTi8Y5xt4aeXRN/
A71sRvN6tdnZWhiB6fJXSy1xxEY6h0UenLFqzhl6QL9LhrnhdLfyFGlPbuwrvjJNKR3iIU5bewuD
QXcTdVJyUPQRrUvBJwFvPpUVUfa9+/f0h4ALHFe4gG8EAsbii6s7MdNlb+CpLedHG6FAPVGXJ01f
0nopacgI9WpZKMromWy5/SxcgsSl8Wtqqkwgz+3vOlxBT9t9RUjfej7e/B4fjmBc78h/eitiDjyv
0TEPMhNCv2dskhunWhkX2MzXiLSRZUUYZASbuzLeMsVS4wlo8+MEDT2RivnEd9j53Ci4Va/+aexl
L5WLBQGjfIoWxnzIXnNP/iJ0xr+kKf98x924TDKfVvtayiAlCEuVjS7aseww1jU1Czkie21As6I5
nn9SdkomY6EqXReVPhyGXymyuDVibdjKp7ggOz0rqpz7cCMeA/4bJ6ylVS5VWnR5cy/4+UIp8Ei6
dPXOf6Z/m64b8BAg6APGXyOqUD6OlVTiJRUDFJXZfFg/IfReZo4wzZFeQiGaXzIG2sO5rwdl8558
nfzj9+i3Jim0a+QS1j+4PubAkRJJB1ZtwJR0jHJtIkHMTaCavuV7tkvH61px2B/zrHB+/v5Y57RF
JxKSo5/eKU5Xbg92Ke68DQF1pl9AVlHnw+MeIU/igB/WYTX1cJfRvsDE/Ph5Autr3eRyi2KSAJMx
AiCW8LMQRIfZl3DuTrQnjQVZZmeKxYeidQe0wecd5QwXgaHlOHz6JIhg1Jkjp2uTt0MeMkbFqep/
21elJNkY/NhevJeBIHq8NnV+Jz+Nz4SOI3Hi8Ny6iR5yYNAifI/9GggRXdnt32PlZ7mz9QnETqx0
5JKQ14rgvfOmiIPnR0aTC3UgiznCvZwCNt8YVMr1qNe+jXkgg5BpAs2efJJynu08hHfh8QUhT6dA
HDJtWp5uFfBhzPo1BU7BmRII3R9/cIhZIx1dZpLK2QkQcrmLh06nI97oCdPYhym2i1ZwaZsLhjBP
2n1AvC3ujAJH1AQzR8wAm0pfJP3l9VF7c57IXawA0JeMpx7fz/hc6cE4fbnxanqtEMKX6AM/zHfZ
gbGgZDOIaO8HpczPGpj1DXqBG3gQBjkum4q083Kgw8J59anRL11DOxhL/0LjhFWw3aMg46wYE32k
vTf31/b/RpWC0bWIMLksm6LJ+DP5AmDRnm3p+hCxofGE7v2zFMzJKhKCOSwNYjVcmq8fBf+URoWH
4B/QPONH4kmf4LUcfbwUdZOjPRPtQ8fRZqi5sD8NL/xTTEmBmTsRZqHD73n4o34MSXyIuPN/AXxJ
Kf8ZTiSHPg7X2qy1I//bjB+dVKM+dC0TrZWWfe2GUtmFo5Kw6K1tHaa4Zt0ym2cVd11lCD6E99sw
cICA3uCsPBimL5ZLJAkNx7S/1oqYWtxpATaGyVWh2Y5xAwdImIBdUvZvtnOXY4bB7j+AtOIBfEl7
No4+/HePu9c5etLHXvKROcl0GvU8xdG4r39AqlNgigwCaMHnQj8UKugmNWxyFZmpRWWWBUjTOWHc
55+idNf26QuPyWIY7uGZSRjEXV9RhaOrH5uuXqWFtFwfAtCpCmCPfKSQMdXq6XWv5Ay7pxtPpYJr
wLd4XTkSilEmaRkkVWRIMj0gUCOrREbMD+QLS4LlFKh547TWwImRRMIIZB9CW25yPVLoCD6JNGe9
Hje1JERjR89L5+jj1klyKwNkvJ3iWMRwr3glnDIRiAnP3cW7Mbhc8zWkVOMdayBM5M0ABlC3APFo
aGIOMiBsWjwJrzCt0cafnafsk32gDCZXIwb6R38RcyUGyTiHO+g5ujdy5vSPPbFdacQOcOkGysoL
UHi0/APh7ilnlXxAD2IUrPmKizWjzjiNI8lwxjZSjBpO9XPMst7uT6l0Lt6bdPNd46OkLa+ZQQUP
wMWDTzudfzGdW9Ks0N9OuP7ZhV68LMsdylVff7rQw0N5P+6L8RFrhx1s84wqT53O4lo60/3rVPoS
D0MX4OEwHEYA4kTzWlWqukqCYpXHqAetxsS8rHC6yRmMxJ+4b8P2CjeCAhPBUs831s4iVHeLMj0b
BjyIQRYiaxKJ4z34uSDuthqfW36wPXm46CcXc57/m8XJymewkiPBQtHqo9Mxi6/le7oruTj4NKSI
iisrA/s0AEAQt1uVqdAJSCJWMBmW0dLs8me9jOEtB+3bh9kFgOFt2PRKq2ETcQVzXWlJ3iElz5w3
5HxOlqDB4uoX8luO5VF01sMAvDarg6TpYVUliVSpUhhYjmZShZtSynDzxvULckQuIpWwf3c893su
xthi+ggiLGLqfxGpEq5q7mPoInboSgsBklFBAb8MQArQkHXz+CtYSK9R4mhM7vz3iuRTSpFK+o0P
nyoByWNb4T+ZnCYXUQY9fgvJilOIf/jHlGWXUQid6YyZeWbYuO/iGnIvfPyYNrTovly7y4MwHpgg
5Um98D2JjOOV2iBlEg2CmDgy/Q+RGDgPrVl0GI+0nbBIMYQd4TB/lQmIwN7qQW3sRTqsP3ekX+/i
B4/oV8U7r/quGU/fvFj82KsC9h9W5SwtKL65r5A9+QPGlC1kevapcHdfGc451pYpxc7OpGeB08J3
kpPgBIYlxTZ+PEC548RG7GdE+FZ0R+QRMbBvFQFaYb3wMgsMNdz7MnvY62iywsSUNK3td4NW5A0q
2OFNc8YfO5EzBYuoLSNOFJAZAQFFxIsn7bSlXXauH/g9fPliFE+rdK2j+OwvQuePG3P8oiKIl2uE
jjIuelRv9/U/gajPLxNN2yGrPa4fTjUcVTDFWfTSaaMJWypFpHxwN90R1HbIv/2kFhTzfLZMb/4z
LTDmpSGhrxuxS4wccvPkkVqo+uQ8fADWUbOV8vbdDya5JPD804gi0xPx1QpYpARt8Byx8ZXMOk91
n/0wbwUoNcuwQK3DaHt6aZuACCHGRIdRyBptOMZTcOkxr3O2MJOPSzjWM30vv6AGcnkO6IMWfVge
vkNtZT2UcrHleUQtkVD3kzEtb43KKSES5UaES1S9cDTgs9KlcD9wJ2KJW7f4B7vA5BJMOtt19Az2
3KcwkhAo39mzhfjD1JmaxnmGMDbAUuZqhLt/rImPTNh+FZadL4wjrl/gQx1hAgTb721/ERPjOFIt
ZUuidGrRHVsH1Y+BDyhFEPnDwQxt8ORVe5Tt/jAQ7iGZ7scXxlTiLtBTo0Qkj4zHXEdEuau6hutl
YxH0FVI7tqvLafM+3BQaLEFxdDNzOmNNMMPvlm9rfnMAJ7hwO4uwrfafwVeZS0bwotjumaWFT3mt
adcuhrlmg/Xa95RqgNN1Fvl90kbyQwa0TQtLc0qcbHqSe1P9jkHxns7TxDwwIB1TegLHoULab4Xl
fN/MZue9dqLWn3thhrXobraTVdbvNrozuVlXwhRRgdi8ihyFKYGMngu/8AlpqOhyHPg33mekSG9q
fSl+w5eMFtec4VFR4v0/HMjiWR+08DYqhe1hcTmnt7dYgNvIJrJSratcP0cKYXIhHSxd16fI8EWi
xNsKLINrmzvNddtEc/O7ABaQ4u99Py74dXHo0PH53M+cn4ZuAXlNG0GSSpVI0p1O50lpCZg5iF9G
pZRLz2ThTzM4MNh+P1CEwBSU4z2lJQ7n1cBzQ7eH7EnMGh5fYkthRvm+9Ft0auvVn6oxCIYbez1q
64m+INCV0/HlW09J5sbjRwml6p8vYaKJkKA9Rsb8G2ZSqKlR0q0lRyShf0z+WfZi92evvbwLDfi3
X5fgqgWRhEFQE2zpWqiQkbN8DWHlvLLbn9YWkKuSZTxwicwd2YLj6mTGxL1sr/XZgtIxi/hj97aE
9OYv4N+lDZZgTTkaNsnvfQKH8V3vcEErBvFy8gXlYq3wyFvDE/jNkASzcA2c+hxCjXdkoDmSqADh
fi9Wly6K9IOjnptbX9JHWgmsfezEKATJrifwwosnXrlERSNz0ln52k5kGxHdSbeCEr/paaedyN5b
z7zCJquLswa7dXDBzsMhQPA+tltkF/hHmxtLVRf7OFGOO1C5IdvaJxItful8BWl85YAUa40dfqwn
bcR+2rK/PybsJWhQV7oz2p/+UUsFA3oykj2ixFluG5zjCutiR9p333iD1GoKcsHkc+iYBYanxTHj
ogL1GXYqUzGSr5nQTw5qpDL7UBvAo1vaCzidysm/40pEWydN0G1Nw/ft3zoIH7Rk4PO+4nGkGIQ+
DonzMwLgQnTSraH4FpG1fw8vEKQDL0LScTSZ84e3BThDcCTihd9XDzrReHmoE7YeHhvHgeCxq6dC
GZm02ZBSRsKd5spyXYNzxrebRx5jePsrqdysg3nGdcbQyAvTg0CsbUx2oJ2SnBV2YwsCikV1q2+3
z4Dvk3/cDL5DmC3hQa2Kc1KkQemlFLwg7QupmSnGsJ/JO0zVBRXJ0FAnsJ4hNygmXYdRBJO2qEzR
RB/6NGSplpIMilukhOuhvNndFnZ8DnrM0aFZOH6DTUm9hLoPc0mRiQ6R4YQ7ObDxOAEtQMTuTmHT
e/ojK1BCymH/qTfnW2f19flSFaY++OZtsoCqSaVo0Vq3c6XQoTgF7+foRHzYQzcKoPdKPt9l77nZ
kxJKN8eySTvWI33anyJtoE1EB7JpDVeJlp2nRP8SEqoxf3+4VfGNM3y2I6vF3aDEhrpdRSJ20703
rT8HUGVNNQD+Jw6PiQtanBFq0TW4JlozJO1LIQtxevYXF8zj7BSMIc+tMp6W/BpAMcoOTo4hZ6UM
0eAiKnDT8uKauZAolx4+RtImzwd/Gu/drkXI1GxUZ27zZTLEmJ25mhsae7AVVVf8J9tOh+D5rus4
9YT+WHP5NYUAWwHY/waExPNLGp1BFs7eg6Mvhp2WAevwFpS1iRbHDqn1WilGQ71jvAcog8I5W/nG
HmKBzyDQKJEqKQfhHGjj0CrDWBPSR6Uanglumm8D5TJ3Y/dJ0v4rZcayWX8Gaq/QPHAFp/+nT+WP
J09goTp4xArfN7FWzzcaSWF4+vIPkEFGUidqFlHtGc4jLvFWgSYvba25uecluqCjqNJu2D3ZcorU
ZTMbBtGFBHYQ6GWcWPGjlITiKVn3jo9VLveVFHQ8hT1M7m/T7CoWo6SDWciDXDWK4hHrqH0Hg8Jn
QdrfgR+153Bbrt4449TDb7S1oOs1tzJGEnxAYjrUmT+BYkjSd8Yig1Zyb8d3HpvpKqIat0R1i+qP
utGwYf4J82iRZZGz6mdUoc+Q0qmRJg1O6UpSDGyDkFimxO8teLmSXlvTQOCwyfk4nSYvbpJm2cvF
yPdfP/9BxWT7Z9kVW13uwQbREh/MLZRTmsSogs5pyrggkhN/elMPi2pfqRHfZXKMXEO0RgBbgI7Q
kJX8RsKOm2U5MktMMSR7VZ5Cudx+1wg9j8TdAK5rtkPUk6c0U/v+Ifsz5euStZoFzH9WoUBOJQl4
bCl5nWiZ3I5uwctVGPxFOVYrSvZy4mrl30rccyohWn8uay6KRXYJ99+o/W9ItgxEi+Vbmc6umxx3
npMDwxyRtG+oz1xLMOjXU+DQM4Y/SfBpVqTvRSDGdRF51/Y7sS5c9DwXsUTfv5gF3+Ti7KeB+o63
lG/u/I1/WSCl2pOwp7ZOdwv8llnhohfW98kSo7VJ55XE9INzkUXPeoxXO6/exTtnFSnku3sIoAAV
VXjknJZ9yEvmC/pTG8saXCDCO38RPsbJQEVibWo08SLWGVLxP0oR3NHuKayWQB8hvdW86gxfOEv/
8yrJdpPNqQ5127yNk5OlQBWqQhb6YxOsjNj3jCeaEc6mAGKPF6/RR/h8PFrdAIN9vWOL886NP7uG
WiUP/3RXsHMKAyiAJKPfFBzKPAia3CAkCSlDMcbwRzQQ5p+5Z6yQ3ufOIjJp3kbMynU9MYqS9GyF
nXgM3AoW8zsUoxWGGr2DJuLcqtwEoTUGrTwNJnaAAfnzBDR6GBT0fMh1Xt7AIDTmUUOVD9Su9S1r
h8BTVsCIhttwO9My9HXxyizo9P9fQZfgHFdYt+1RODKZvgRgye3eXilltwd8yntUMhGo1mSd6fML
J+9wXF1fuJVUnIDyuD1Z7UvTY24FVagPBUz/oRcalimDNuxjlQfLCl6gm1hKfPSZGrA+y1iw3MoA
38CGiRCKCBvUjV4OLvK4034g0tMumqRzl3ZeieTNl183TLp5BxmamkdabWUp3EPM7pS5+d481QFx
KCHdCfCT1vmxaYr+kmdO06A48wAd92SxvCQhT+kGvSaVd87MvNcQO8GliFVmogrbbPYTp39ncQQR
DHhTAasXffbjyytHvCFnnLtpY3ePJltPyG8WHzSevlCIA+UMb/ggMpwyJ7LjnWklMXwojqIOdoIG
d52GbR8B4TMyWX8Tb1aIJmYAvEdv/j6BY4oo5JwATOFwdS0WgyfylF6TcO97nLrnfXSbPEHv5Nap
9mavUcWg0kQNcXwGW6b+UAB9MatV5H0amodde9THguFh+IKdyjUTjj0LsPmmsDJjGAym/WhWb758
bbZ8sYR84Xn4uVkKFez7gObh7aq53he5dqqw3D6Y0YmMbuPLDZ0130RdmSZQhWL0fAJq4gORRFvp
g5Hs+FAvJjDSYxnZbPizDrad3k94GPbJpNUJhGGC3LSkYM4eLwAVRaRVH3s+9vEuJXNyQ1TaJYGy
17o48WZ3haKahZK1MZ1NzvvRaGRNtyqzCMCS8hXdhMPhhIsK4CJioTBW3WVNnvRnfg5Q/mvvOAn/
/EFAm9hTVil341G6LdpUoOFb57rcxY/ZairhImj63nYk/xac+ByeVPUa/w9yCMP44KL+xIC1DNW3
eeatvMrEzbnS5w4pDiEgv3SYTzgXNrHzcEmWvJ/ICnqGs1wZtl/JbMhLFcdzTs5Z1/N4qhJTUGJQ
fK8xOourxiRzX45em8DU4pJHBXRMacZFsFLTkkpTf7oPeCwzxLoRXvI9CjM+vXQM2rr0BAkyLlUh
OsYH+yyZJpsgC/H1gvUzPDtnhzH8I8iLtISiTrP52Bk0Vq3bDvYOGAVmbvA8vEqt433eWqE6a+d8
vvK00juHqa1GMuOJZcOH3yxcKTkNw28C9lBWPiEB+lYUnwbrEEfYvUJWkrTCZqo9I6wPScCc0vI6
PHV/t/q2dmnqSxvizWx9AiFJEuvJXNFlArKd5tp+q/8xrBachr3t98Zgmol+gL1uJEXr5MXsi8aj
A9+tED+37GclnQ9JOv6NYCQLVwm6wOKOUw8lXcXTkHu1u+44LrVN2SiHUqOeQ8bWZNI8q1Tal156
KN8UzjU/fXAkslILb93gPGYPagfocJi2b5PR6OV2SsMTJwsTQTKKs/mNvUQ04PgWyr5ej8ojqGP0
Vwwba2BiUibZpstlmilTgdphsc3GjYXQoJ6qEbGQ1m/PPA0De3tzgY3h4eKKnUDU0Z/iGhNPiSeJ
qtE6/9O0T8tfeDWbVPuBKKWRYoH8Ty9askJE0Mx8bCJAnyicpNBEvyeELBrZfR5XcNVg+idgbVxJ
a4wDCbfV007GI3F3+SdTdVWwaJNnw0E4AkMc+kbpBKC8cgTboYG1xllP9r5aVt6g3xqElXcPaLXg
FvD4aNzbyIvoq5hYXHjSCOXLOAgMjdk0kwXPw7/xXpzFGuSnT0fZ/ZtkVSoHf88/LGmC3AVtgXDF
/sfoKmcU9UOJFPUFcdtE6fojtszmHGwzbSedwQiWFNoYWyzP5BJtKTrFJfKO0g/WF/Ed292ooWLm
fetPwuE8yTHJ+UCgesUTJwE8xNL190ZabTNItbDGHccRfSX2LcFB86okQNk5FGPE8U6VOqu+bcav
Jfv8tUIy5bAVtp7vzbWYrOJPLW0kz2xmeo/xOB7gLpKeVj2UQYs2Q2VNiEQo2xg6iFF96a72latp
pRWVWItelj8yY3R3LnCoqAaXfW9E9HE0jJgKR/tcSHyNl6F8sAaYUD0xjrEQoSA1JkRXuf7LvJWN
Ts+Da4gHVbirVIJ6TbKkkcOxeR3TW7oJEMrn4aQ4FJ2bpf1a1ptb7A05PZR0P+I1b/leW523f7k3
TDCcYMohzn3/iWPS/YXM+PQSj1jakuKCbTZ6dxZUfZ6qZgMysa8bepmGTpB4XpSwXhqAL3KxAkma
1KL4INmlO2CtWajJ8YkMUIxcDbh5+E6VqHyaDUHg2xxxodXlttz0mlHFu0llpG/xSqd0QYFTU/RX
A+tTt9BBtUsYjUXLhtsUWcvF1dTN6jQ02cL+JkvDZe6yzomw8lzBh5DCPIzksYHPI+uZctlLmhWU
gBiYvo0ZhU0afMcQDB+2sHupfmbwoncGnz/bAg4AqU5Rn2NfKEOvVns58yBcmD0aSL/NOeUyiEoQ
JQnVa/C1Yxp2d/qj5zYTeeRNcYZ0nmD78xSrJVmqzGKLrVimKhbQ706jZidj0oWI2VoBV9qNbDiF
S4j1b/eLKo8haHXaTVvN32MwIaDwYPl3JSQQr2ngnaAW/Ut0biZDATbZYfT0ibs9T93v50Nqrm5f
BR6vqNsa5VYJH8kr6lKL2S/s7nKHnloqBSXTvKZaQWyHPMb3b0BPaeVmNq30VYtkuzMRCodP/Z7N
MCkVLpY9BqmPbjRPnpYHphj2BJzdltpZ9XfibUd8Oi5se9iBwzSNJwMjCtG2QBMjScDW+7jUcau2
jHJKGgZ/DVRPnt1ZNJl3xEiE3NOjUHoE7XlDTYt6HcxmFkZfzzzKeMupjHgsgCosiBZkPoXfii/t
rzI+zTjZS8VYQoXRRu74Frx645/YHut3+oLOmGACoBsyX00M+dOahPD1arD4aXTA22mVXYwjK36h
bmHwo1v1g2JckzM7j6M06HqHTQCl/5/kuBXq1bni9vwhha3uMIImKZhvRUjS6vw35/sQk7GsVuhQ
AueVGLtn2nHwr4CpjCBWmC6teO7OTKdC17VqwxBNr9n8PwMrv+fo8BlotwS0DQBFkxEnHVn3KUJl
3TRivO14ltLClHe7K6y4wfOk0+DpImOmBbLsqZ6CU9DkWwQzplD6A0cxUEDbexZfsHOaT3VUpyoi
AjD/aHZHCGWou7rMbolGvFZXwEKxEbg0zUfzWmkplT/DE+2ARNM4zSSTY/TuriRACKYz6mD3h/vy
wJfgdEc3Nz2yRFaLxms815ou26DUUVNNarc968v74tfZXZZvlXbJGjakqwb0bAXr6TsYX/mK3yEK
9+lCl+IbeCOyjbjIM+4hoiI0qb4tKwQZOP4jPoAWt89WPC0tutTpoPNLBIfNhOWxpIQqUReoUUFq
6NdjlLSakRGiA5tzv9ifZ2wzMsCmtjwuR0NEVvNghFa0YHa+Mu5s8/GgFCvwMjPMtzkGUSR+XbFl
EuoDkkI2/qE/GssGJXEQlfl3wyJS4DMHQll4gPhyhpMeKJXRPDTZDsTlYT9nxqYQ0Vn5nGWUWB22
NNUshSEpF0xUwjNB4Ug7+N6HwCdX0pLnjsOyc8mXfPdASvDTcJtPTEOApnLHRcvoSzgBsZ0LOhRH
5f2zpLWzpZFSAPztICT3fkdZRaODid+bspobQG9IODh03He1jFZtTbmLkGI+ziJiGeENI1jJeggT
lZ/lkToqRGTZsMcw0lCSCHD1q5NFaB+pZZ8KhxdqaUHKTQ111s+U5qt+V0VMmkMARPRsLp9mPKyY
du18UjcyEEdtapy4ycSRIjmt5AV4AyYEXK8s1lekZw2zM/ar7HoyJs63yXuhu4ocYSMNSJYAQ8Vd
gn9CGy765nSwcxIVMsP3rPJ4BUzQoUi/4M2F2U6SEmiQtXO2K2Az7BTQp/a+X0DmvWzICIgkLq20
7EmyMyftR7TnIdPbGnvQKldctqiLboj7w20JPA3TaHdaSiWVr7PA2RQw5uq8o8e47NDk0TKya7cx
mUcBCymBTg85cKiXXabPA2cIxVlhUMipsMZaIPJgi5eiVuAlMYik17Ur18AG+dADLdxqQBoWaedu
+TcKeaPBIFiNZl8/Rk+wc2DguH3LbdRZ1GC/+QpO3tcobXRdWZvE6rvYH3L1tsiYOQcJgQu8FN33
dZLrVCtgoIKY8GZ60zCm75zFjXB+OMJ+chmyjmLvf7Betv6CtZRga7Ykvpd9Tliy/XfWJJ8AY2fQ
ugz0sJmArFLW0o1YHBQqc586QUO2xPg5kSmAOjmS5l55qq1RqpM7fUWgEXPXI8ZPWH2l0gbb+t65
fwjjX6FIP7LY1FNPjb8nB5mklpsqOZfmQEKEdHZQAnfpLL98iizJj149v+YYlsjDzjusPDifbOvI
+jIDz/4teEfa0KuUyyOeYr9NRIw9UJeOVSDWZ4CAlvIIfnR6+8y6SSyiWpKI64+7gwzvdLnkgkp/
axX/g5NGNyWatBkhPi8jiiMit7pVpCj4TGOhXuE1x1xdvivISrrEDn6eOxhPrnW4T0DTFCjCIOH/
MUXXyHOZm+ro1s61AYEjCbLJwCHcJuwWhApR8pboDGHhNtrM+KK/B6mCaS5XF1smV7ANqOMlRt48
nAiRkDccozKReshMjDGaCj+kuViimzUt6nmu1Bel6mScVn9teGVH5w40wXpFx5Ktdtzy9cCLkliZ
5cau8078xvDQuM1bjsTwMLt0nzpxj6NXfSE4A4s9nDV7MbmxsDTCOXAmO7QpQ9wkKSQbFBb5r3kw
pLHBqDnWNNjvXMSfknWr833StA6BvYK7i0EyaUygv16ukZAYKhDAE92SkLV3/709c4OSsDGUiL2N
Y7r0Wf9Mznn4X19dTUOf8cl4BegXtfewIBZEq0um2J23lx2aHfHXXy2OHt174kRDWjFbtvM9kaRs
QugF78o7S3Xdl8DIHyVBpoNW74x5lU1MEmeOq7ZeaB1/IsnOrtSq7ysf3mRxDfwQvJQ6cPS+vVbq
ePs7qWDxsYzO4PPUTW57tEeyyy3Eo/l38JTU3gL6MsuAA9IZG0RPajd9EHrUv8xF72RF+qLSYDia
aRQ96tYiI1RNL1j52UPgC+0HpNhbSTFuxlaoaQF5sh0g5/j8wMD9vpXRzLgM5n+EsTi1lRQM9XKb
UpE82atZ6TFGuasY4vT6TVDp9E0DKFn/ZExlDcOXyTkp4ox3+7Qs3jYcSVluEbtjxibCyHNL7YeH
5jbbnysHB6krs4Rqe76444m48MT0AQ9HC1BbcrFd2JJYm2A4fUh1/6/xcFHiKODnE7HbY1Zyz7vQ
JIu/N3o9ed4Zj4Kampw9TX/pkQepbjOZ5+UC595K7oIzNsiXN77fDx2oVowZhad5wkT3owntdNO8
sZl1ZkKLLrktKtKNlpmpuO9UQgCcIHNpubemfX5gDrr83pbUBzA+tratFnG47vj9lEuuRDX8Gefk
hii7X+nx5KhbzLAdtRM8FGnfQJcfX12j6MZECzhFFu96yD43e/BqdbPnor0X0zrgNj4qMwW9mY1G
37/kBxH4OUfVxUN8UJ2r7gg3JE8k+0oGkF/i5WI9zi3FGpy02ckwrxyXBDzR3NzWIdbaN8W9cIt5
VcIa4z4RwZPmutnHJrrhlvwu5md39Td47B73fwyEp7UBCMTzVQuyUk3mzLIyVuXEFtYxLrfdFoFF
9dbRB4mGtS6oLxA17akY8b6R6vxRWl0QiOjSQC+S5i0UuHOkYqSBMh+4HEr/yf1V/BoMoEKHRts6
pkEuQIJJL98iKU5KrECAVqWI+wurRIvkfiqZtHUUxdkY6RcEYo5MkoOgxLZQ+MFAyRv8YhnjUNL5
hfT5FHqT2tvhSyNer6LpM70DLwcSzR18gryWkNNRsp7lw29YykUdN7Zb/BEt6yGgYkkaLFj69nIp
e6rCDjrY78huWs9EaiD2VY5Zas9+Md5TxdfT6jRv8t0Fli7WkNYQHMOJEGw1r/a5+HnuTJcjJpdl
tJwtLrR1K6hbd4tqYHMiTRWWpUHahkwhZcSWp3Swwjc7g3duHZqE/SSZz5OA4CWtxRXgoOj+RuT1
yqggMLGZitQHHNf+JXcK4btSa30bFKWEhlqLnWIqDZnmVhJKzOn2h/M8FrZ9LFIggI9FqT6ICwEq
YLyiCs2JEzY0uuEf0sA6g3jAS2yQblfExTGCTGO2FJAfkl/M1W2hZl90bT4JdNP7gIBm8xLzMMMC
/aXyrdcpdrN74DampZnAtfqqWn7SfCw6ngU5mvs6dQBg7tDkjqiVokwvbPcOABRbXFflqXl0pJtZ
R+zj7Tcaz6h1KJ+ru52B1UDaAOx8UYg7W2yGNEfUN4zqNz57O7mAFFLJdE/gFnRvvNZVtztbBvUp
ezS0Z9GCbzSD+G/FEDcBNDe0MeSidamuYtf6N36TyKeToVWrLUN1bm989oE+a+F/UubT0kv7GPfK
m4YQ6Wvr68I3+fC+wVA7EPoNNbKTHOrbijGLR6K26PM8KkvR5Kjqi7lSGhBiZHBP8FAfGcEQQM5L
t4RAOh4ME1bE0fdvkrqzBcHGsPC5RgjwFAXRo0SxZQmfRB/EaRef9L7r2CgmkSHjuIC0qdOhzRvP
Wg0Mh5Cs769Ne42LBxDzUwYPbuXfOSAdz/elfWbDZgeAO75Zcaza5tzUjTAZr8tvNtSrDk+BwHbC
+N4+8d6YHr8/qI5OU+PVAPm3xE0PJGwYaX4GIEKnRKgfe746pb498cLJ85dJWnq4dAl8XugKuox6
09+iVlywIntm14CYwifJuch0tNdEap4tn6+PS/Wr7fKNGCCsyl4oXcEPlj5i/gIt371AomhcPqXG
9VGLVvtUQMBWpmZmH9NZ7ARp65+CiWAypyMrcyVhLI1waKLpxEwBlx6vCaC3CN8uhKsk3I6dA8nO
Jy1H3/UVso8GGsDYJlct8UNAo9g/ZUrYxdZ0zBbnB1pAkCTFDPqgX/bnAxO9ixt8OTJd28DnU8IZ
hIB6TWWz2G3OYelvt9PUQtwnnq+LLXkdHlbgSxaJLCChz1fkDPLSUs4FE9HmXekMamSqCCRyeOaw
A3hbs3LobR1W6cm7aLhCpAWyDIClmFHeglzDhl7+2w9trCAH08AbwHR8WbDb+OvHkEQoXO7YFEnn
QOi3o439VUzcr4pHbeJpXHmphGNaGq5oTo+UPenDPboGzW+V2OqsmXzku2LwuiKPaUJyfv22vG8r
qLNt0YvwTF4kR6lMhlPtv9vpfS/bKT/zjawLRB3txr2wJpuPyqOplgA9IH/HE/DMz1l7xTw6Y5AM
fiAl7ojntxBACxVuKBOL2wuvitNj7KGbyWoa5JOFEjOOIp2bwFirDwg28skvKQku/J1fAvGpExY3
4CQgHRaysDyh/cBwMQc4zqfBcweGtUNgirybnnzR1/RQtK3lcIyTHQxAUaaw3FaojJ9wYq/67IPw
QXBxcIl1PTFdxV1iQkcFxKTt5oPp9Dt8PPsh5mM7ha/gsDPkFfFZbefQ9DthinlqYN6EMFvQooQ5
YHCmFYL+gyq1TiTVyixcpoGhXemoKkPZa7GbmEo1aJ/o2s5/Gqbn8V2SyTef8xTxyF8fflPuxgva
Bd0wN0KtQtZaaCHA/4IU1bn9rbP4cEhH5WdhOR19OKVkbQAqaPCciB6r0oooLo/rk09PB/15z/CP
fv2RQJKPtTXZUTkG7gRTY1ddh4JbTzQRWmo70j5Mzjj9vt6+rQkgDcurT/lFMbuUrgXfKintPx4s
e+cJ7cW0kt4J0NTMlE75rGOnBoc86g3LDCXJHAXqtDl8p6G2y8VrLcXXySuoNNhGoT1y6/H4SL3t
mMyBcHj7g4C6O5fun6B4ZC2qQ6OHJ5SDS2nsR3Ty2ddtvMciVDtofnt0V3ExidXjmCwzL7+QQG7A
VPFgmXe1ikrT5nOmxOooE0gzgGQR9d/b70tLFOe8EO+dEVleThdFPNxzNgueiPAvnM6/IOTxHvTT
RR0USsA6lVbHb2DI+dxmh3gP+vwGSN9z3VNSg8gH2mu0usbXYjZqT9zn72r/jevPestdUvvpK4qY
THQYh+0hqaswOZuUTyfzXqQSinDhVTfRyQlV6JAfxCZT1vaYmuFxoi042KCUoxMeq/v04SWqom/i
JlgPpxaAgAunp7YEKcSZv28C711zuHzo6nvjWJHIKq5gtMnTJPnM0Lj26FgTN56Ecxl4bporVxCN
PYSVjwyktJtmTaYmWZebthSOpnn/tM8+u1ZvQS4Chm5N9Jf2ygOplR31UNEy7JNgnk/ES8C1Xhye
9zjPR3BeDBJmzRAqxqBVWOcOc/lALMzCJBnKe0vFuDCpvr3+vUoCaGMsWrxm+O2+s+eFwQGuCbGR
5p1px1y8efjW1Gz2MHV0Kue9qtArV0NWJmvwa+yGLsmR7xXAQ4DhEU0dS6FUlFeZAzhfEZfWF4/I
H52LLhII0qJgIdUVcMdXFubThOokdich2T20wS5CPmLArh08aePjs40Zgc2sDjPjfaH/OAadsxaJ
7bo2InF5QHHAOGtTKYO0fOyrs+qJysvXemJr7uawOf7tZWFDXJdNdWxo/zTQVsqSi3XVrYhTRhsC
HUA37zcKeKpkp8KTUA481WY436VzGkvH8TsZ8sWMN+5EjswCxL/xg8LZzFc3/3ns0Th7pfZeUtBJ
rA4loE8orXeREsaWLC5IlTpw8g155OwoY8ZT9hcC06O3tnVx0kvi1qwclOphGjPnxrDfA6GTly8K
vuJjRnLgjvaxBPIhMis7Cag21fstLusbv7v7/XWQFGCIBXFrZGu8qTlx4KHSFDaHRSK7Qj3tZRo2
cPVfVwSez3x7TmdbM6GwQ+Jo6+JfrHofj9vcbzTwXZjB/IsAZ66V2WUMvgeNWF/qA4l+29HHLI+8
Y512bLGRrBd1SQHB8s7FVxGdJTKNCsnj5VYuyC4O5ErJsLuqVVLoc8qLQW69mF/Dy0W3/h9zL1jj
D6ORsV1fJFRs5ZDQlxhBAiCwYP7sXeCYe+AcsjUPuPVn4rradVua65Qj10cqcDlICTCZxW3ztYJh
o142oRs5ra36FhgFRR4AjcwNy0a1IBYI8u0zV8Jj0Dk5QOpL7AntrdAc7SKWPepnQF3loapF7N1V
rPOd0Mf9DOOJr7kW1rQhMNzQ13joFUCEkuMzzjUj4yJscbIiu5KPEhWJPXeYw0irgQkSfKzSnFcq
YxsPS3T16eI98R45XybgCuNnRzTP5L1mDhRB767F2x8PDSgWPlb+dXiamsOExaperdkdDps3yXoL
lE8PkXnY9j01yIzkE1g6vfp70VISPNSxEwnL3vtAF/hFWkX8kZ86Qzxy1TmPHO/pdVXXbfSpSbSP
PZ3M90DXbfC+t5LA6PcInLGNB7dim/p6UyREPZpHqQYY6Bbv+7OthBUqBCTbbCEKZTnkRUSLZR69
V/7BvdDiiuCb1nb8rWnhvyctcXwcs4lbyuWUdb2FFnmmTjCFUgFaWlb66Z1pp8k61om1HdyAXYWO
0VCXIirXMzvbhufP7BkoyPJium/BdwTOFg8fdPGVv/aS+hZjGW9Fd9DI5+IA4cMCHGeN2eppf2zl
3DPxppVhC8oCM2MdOQ/NXCr/+tLmWaBbyr/dU0s95IWTGTFpZ5xXQISUIwW/NpdXZMXOy43EKqdi
HSxPimKJhqEOdPOOr87OLP3I+uJ2rWkQlZB7nVuhBBqKVdILHjSijY2Aendkcc96aOnlIw0D1AHL
S1SMurUwl7jT7bzGry/8V77DGIlb+FQu9yfAsXLEI4V7fTicFg39hebnc1O6Ij0owrHl7Hm08d0p
zy5ISd/mlrQruCIWYB5f3XUQ1pbj0jCwL7wS5y2Sy4jGAYtppUJf92U+Rwih8FW4oNuQeE824fIk
Nhj1GEqdHjMNSBUCmTbBwbk0gv3a+x6u4M3SK/QH7fc6OZ0nRPxbzAf7TQDPINHxanF69oGNvjsT
qSD+nVbJ9vtBxJb0jt5x0ZW2pa9HjaTT31/0Lk3tG9mGsad+UGJO1+QujRB23v0GxMxRJKf9tfZl
5n45Im0tMqf8UXoAHkAMX5rGVbZR1oxnZjhRibKlJrxMdCKCULs4xIxAdhiA5uIktjo5YxLS1AIh
tO3F4pjtDpHHlpOBl5dO6JOHbZqRHv/qvpk2IBE9q7J4zSksA1Zx0a0gAd77NUIwA8wBSVa519mx
cY+0HrEUtFi7Ot0DyQXVv8tFwf+rtcj/RO0HHIxCJaCnIRzuAxJGVcSVI/G3I6j6NcmOUuQvogCC
+KBAaNR2581FxoG6N7hvrrvxL+MRqoQQ37Jy4mgbcLQJMMt38jbHdTwD0Tz5gFsvAixkrlvTOXD8
tA/T9Bs1fKxhijICas5dOSZOzhSHSfUIj8wFcVtsqS0rX90d8OhrVgPFkwF5pJf/kPhDVYDq+cMP
IqhWOUC5J08Es6I1DQxKNsZUbgIo9Y/0KF364uAeW06Fb+xwY4DLcwCWsRpy73EI0GiVoUaquSS4
LUDR5uiqIg+U3kdxsYwvqt4P7b6dsx7A/zoR5dgMMAzBKnPkDou0kYQ/k0cYmjmPljvZn/MvHJhO
JccUHjg7rhEItw9IiY2k5ECRWyZYKOvddEBaXQ0T09z9SVpMXvsjHdmCaAvNc8To2vcsVqpCJqeC
NlzAJf6va3/5a2T6oMhzBozzbsKRj+DTyxzNBCsZEKDMCpnUeCrYa9Ou+cspqf213zcb9I5BoBO2
0J4vWZV4LPLhGrNUJMshtohZDxmtXNwYkqnP00lKZt5c+oo72aaUw1ELvkXTaOIhv9Zo5o/y9v+S
VJ4aE7a18X4N6pOIjik9NQOF9PKWWafmRCzUEVOL5ahVyViUBKUB3r8O64v8vY0yDU8DaTFmkdTI
cZSBnCOxL4v+F1UdtOhixPCuJC+xkZuLotXwpfozW5dzalGR+Enl6wvGW2P3j7ErkMC+UaEhxSdA
bjw9M+XTHTs8bi24VqF0K/XX4ABguJwkviGbnbAPFOIDB0D1eNhMFcZfTYVLhn8Y1ppk1u5KBFZw
9ZfIz0q60OK6HgO3/1yJaVx4nT235Jzb+OBhRgs5hWwYqmgBR2n5mNYoHWcWmrA6eSJYuE21IMZ0
yp/zpYqcxQ24NeWBXJUdXHpU8V5Z1Rqu4A24yUmWQgXElpeSLePQ5g4oYuFGutRQE3wOiq6Y6YkM
03Mbqk9GZDDpymTULY4R8g1wCqpl433r7fCM6NkvFXaxeN6t09W8BDl4YnL5MAAXT+U7WkYwYz0b
7I2s318H4ex70+JYFIGQkFmNUBDEHgHqUyqLVX1Gc9x0CSnFaEY9mXkjz0+otobGTUOLoHNyg8ew
0GfaBOirrrDya5+65bh69waTMoXXTJCCyXS6ht9oHSiB7kOhc+FwYb0sodFtJavTO5h2axzm6BLw
v/kLpTgwMOLI8mZn/iBbTn9iNbA6cbmcT1tUB1LNxw+1TgFeF+Iu08Hr/5CPeoWfIzHwKCRQKQ05
8Q6lrEcI2qOxiVk07U06zkcipHsbHYWFXy6zXMlhn6MZw8VFcc/6TfxUpqMfW5Y9OAZKX4QcHthS
5idZd0cv0w4rTOBDHXqaDTRH5RzRRvQs4Uz89yY6jF9Tttde+w3Sb1/Zy4Dhr0FKHQe7cNhkT4VB
lqWqxQUKEYbz5R50SNT8qoA4gPQHjp/ugPeHTG6EKzSZzV8yKDq78JuEwkSqmCa4P282zGDRiNhy
Xpv2yMaMSPFwHrkR+UT8HPsZPVYTcH6FsrqoaJa6sAcAPlPgOxa6wV4aEtcpmSEGSkmwIEbJMXxJ
GJFDGZ9efNyjrIDm/N4qYZWCcOZdzPrOQ4/qOYPC9/fj0RZ6aLR56cmt62+3KeNRzk70UlMUFKEd
DUOkGWKQWbU0v6f6tglyDUHru1fT9+c61nBAAyiICe4Sz6NSNi8+y1+wX2zXXXqiBEB78lLYiLvj
kiWd/BgZZtI0RVU9nW+xKMhUWRehD+BuI0IhiJJjqOnt9EwhkHgzfuadGRlu68jXCpiQwfR7Nvr7
uKBjZITgYpJx22KvUQkbVWwJfn6DZC/NGFKK8UI9IXxXqkGlAawyy3ksGRBSxOFh4bF36pgbk35z
R8upft4dxdrj8pcP3Hhrp8gmSFo9eqoxUr6tqMMFOPTi9eh959x2tDnY5/VwWnZXquW7scQsVWeE
lq8c0VGXbfbXLTZeWC3pj/ePPLDLbaniI0+Bx8Glch2NKuxtab7Wa449/IsUYrXaOh1bF1TSxHRO
YrCf/wFMm+OgLX+6akaPz4P023AHwM+gw0ecO8RKqF6zgEWFFOAg+6wQQ9OkBKXhM+nfSz4yOYHX
caj3i+ukluo/vQcfZc9S5burTw3Cw6pnT0OJPm8KToYDFHBWPz71NPqqBdT74wW9pVnUfb5QyzfX
nHKh3GcjvdSnNatzfgNTaj3qideAkTkNyIlIV2SOcMWc2XkoWTO7secVbUA6uOtEhpJIZZ6PMRuK
ADS0dedrnKoOJQ0UWY8/xLYLxCrIDk4AHN8Vuxe+Zxu6JAuSuE5huZirEcY+6efujfaY2OLAUOzc
3rS3w87zFh7/Dt6SCEIGmbsrsTRyFwkF8XzOExk7ASKcpQPGvnsMpjylMx/onKcXQ5t7S5zBEYGp
wFWYp3F1U1a3+m+5FXoPtblzcltdcFQ6c/s4GFjxReFZkHIHFEbWYbD8IM11j321maKbz/9PJVP6
JuzjoUgU8r1lPkUlAv8Zjws0GnWMJ789JlbrQHXWAZPr5qunXdogHsUMsg71LbddoTT3uq4bB5r5
ZQz432t0JecihspF/Q7GwasjvMYT+bUn3l28krxGNC07kkm6MvZjcmC/CI4V84kkFmfEDdKj/LoK
ckhE9TMawM3vgP58hoJlDTje8GcmCKmyl36vRXGkSh/aTo2SaPOy9emyNsTGlPLZbTlIqNFhjwkX
XVZW3uMAxWeOvWniDkAfEuXdbOaGe9Lh36FiTey/A++R6UF3UVnBFicnrAokAzr9jqa0+LUVfYF9
feQRKIxIPrtihmj19zWFaTK6XIhPFrjP7yYc2Sxtp4O/ot5dre3/C1hQRxpnWB9FyJR2EA3fkBSd
2LRThtPbN2jBGmdTX7dSZQKA2xOciK426S47BOeurqySlKL1XBK1p07PBAsz1XuQKIT8MmD/2Yxi
+UG5i1rSg2XMJayEtSL722y61AB7fjH8SnYPs041ZTFRoLIf5Zd3OAhvxcMYktq+phKnMiViixZp
a6yrLXMzNzOLJWdZBZI5Cs/X/K7R++P5oDWyjqjt/ZZLypXYR/98jTpkACtqfshtGQ9J7H3HAvrr
GxIKb/GGuYYWSZFWWnt5XwLi8gUEQJEjRrXR5Itd4QWxOVWsxzM26hFrIQ3HBeLFI/yWXwSmcHzs
kn+htaSYjw7NSrZMPjx9iiPBfQzniRI56eD05agiS0jPrB4DCKyE90ibOXTtqhsoQlqW7ZI58l3W
ONMb8ZWdBw/IcWj2HuxQF1DdOdfD2jEzAEcgsZJ1BEXOdMRpzQ5fXcvJ+psHS6slPnKghA2yM3tw
yzyOVJi/DKhd5gupiw4Pk/jHrKeX4AeAAOmcyfsAzBeHwIrtB64bnmblyOQ/RUSPBfAT8L8kRfXZ
ftLyDEDz+vkXlhG04XT/n/Drp0LzvFa0FApTHIUfUZPQsZXz63AOkIlvYREvX/UertpRVmivkoN8
K6Y3RGKONe/zVv+9nfJUp0MBHWxbSXE+/Q4CpZ67RrUw3G0f7T/bqKROprkc1N0Wo25G4rOvKyfg
sr/npMLfrsxs8gsDaEX295UTNRdR1vimCh4fDh7mdCcsvlxx9jYI7YEvtABUlv6f9kbAttyLlRvh
26R9Sbkcsq5WoV+eViBK0RxUh8Z1lB3Hv0thpbNlBfDfEkHhysx+hFhjxt7VUj7VF2ww5R8faOnC
ztPibm47XyNLYcEWFTuNaMgsFObG2OQzvY0JCwNMQUYHi8EnyhoF9VlSirRGdBanUiDnwuZ0T9XO
r47WPDawdL6ctMRialK6N11jk9kPgbdMi2oaLzW2Rpw7DkmPvOmwg0sfbLYqFw9dSyBRViDOFTF4
meCerEi91buJdWQGCdcDZdSpSy+183vqIRWczzK/zvX1UqPrSCDPSUJGH8o9/lEeD5YMfAxmsNj+
ThbE6tWQEY8hHjZi6jFxgyjc2hujP0IWhCy3gS+v8zMFXyHaHYw8eljdmH8SmmPnl3Qst/S7gyXQ
iQ3EfhFUKYn/ysXNhkf03aVuu0T3eQyUoltd5CjduifNHcC1GptH1KMw3+m2amPISaTnQ7fSjqPI
/h5VfnRA/srbFrz6KSFH7I7/wSjXhuZZtV28wu944j7WNeCvsxo6D0oR841lnj0XMOb5tgMskavh
z8p0wncqrmiaV08V7CoiGe1zznQg9OBV7t+Nthk+yF6UyPUKv4n2C7ydbB749FH7SiiMSOoqh7ph
LEHZ+9N7VUsN36zME9WZOAlWqez13UfEj2AKLyyRV60++v3LU5Q+CZ1q8ItMw6xgdOcg4umY3EoI
msWdIca2L68Y5ERRQ0faF2d+vuQcC1ZBu/058EJxBX19m+0xha3T0z511jIfGa3e+ZZbqXCe/m4b
1jqqhEY3V+Az441onV8H/5Z7cJPnBOMKWnM4jGVX1cbxWZqammif9oUuqy8ebbzp8MLq6RW9jWls
MBiExeEbsuRVx8+jRnOUoNoUihuTmm/PSV65Od0LA+QvLKymfjB/usBCXzvdmwFGfDFVvJLwKJx2
++p9OeGa4lbQTUgfp0mqFFZ+FwL12J6H2KeSCt4Ao/b24ugJg4t+p4SgMscMYYyqmOpDFIcz2qfH
coiQUl+cvDYo672T9kpsuKvWAhod0isjqSOmwGeMTN20K3WJs926m01/A9niR200uG0OsjS/PdrQ
d7/VntBzdic1BOUc13h+7QK7S1crZpoj9ppB25EIwhZBsFDEaX64dj8Mw4/lJOXDUj18KwglKlvN
i7CJ68kVqmpDPl0XtMXnsPD5n0pHQc8pQxcD1C80DOnm1Jv65cmfB1A+0WJ+Q6KL1SGuQg16WzQf
/oN7MyHj07aEFJzYy4YEjMgEd63pTe/0JAXHp1kR2gpezM8vyQuhkWFTtd0vSiXzss+whZe2UfQL
svGzGvy0tEzZY3FAd46m3WmpBsuRlbnw29NIonwFaKptWPZb4uXI5MhNacU+cAgXEdLV9ekaS7x8
KQh4bjiyi46Pd3XHwui8GXHbBhUXMBS88dRHZVCTGX0Igf0UxYzCfGHR9MMZoRqg9cG/UbG+e+oM
WUn7MYQBMTmAS1wpF5yAVhh4HDQCkmLbUYKrMg8oxw6kevggJ2tEnz4gxPT2hlrs198mm6eS2tm4
IvfgcVKWIEz0C+C022AnozMQ4o3RBJe6CF6bjQ1c2JrF6xX7eGy9WlQzo5yZhn4JGxJBhT7bglca
vWtpguiUa60H2EJhEB20nscv1a99ZW9sY1DK+Grhp0uct3lgRgV24exkGR8MgdBF3lmwLBZmQhCv
JC47rOv1XqygEoFsV3Y8+5bzvKfFbo+PPcOIyRBdKxR+fvhgbzGBX+duTU26wC3jg9Y9FBH01yEq
BUsb+JUbR9WY0BcxcgI5b2j5B1tokDQvkU2XFp1A+WVagz/W2C/dpX/I8p7HgphtgLMkKb60WObR
Zyu7MWgfvp0BPCQYfBtWr7jJiWti5LQDstnOPhwuPiGoIsgon8SZu4c8dF/ii7P/W5K5BmMHkPwu
kQod64jo1/z0P9B156m1iswdnGkVHLoC1UYgCSCiJ/EBcRQOxMrO9e8YF9Q2x14ChyEaNrbiXjWe
B8IsmsRYaKPV1lJ2rPU99Jbg71ZNBzamzgKs1oHPlaeWSkIN3vkpQkNB/WwCQnET+BLiTiw7dWNM
6LqePpmKjYuJz7nQi0ui2IHR0GinSIjiYw4DzzHJQoUsFWxJMdV1qxlSIlvZmVqSlBAqtMdonU7z
LKx7aZQUtMrMS4+9yeU6JwOLb+xDrupuNT8GRui3Gp5bOfvHg04Y0XZ/jqP8teNIpJbmhQuHm20o
IPyCA2Ef0D+/7ph+yWlrJLaOBXJkUhvCSIr2JDFtIt9uGNUE5U/94dK8DqsHB7hLuDtloqK3e/mY
7P7lpBUco5sEv6ke4XmyL7FWz/d1JFrQsY8pTBdBHafQLqDRLlMuF9fc1ujpCdN6E1MD1s4zUuFh
1EsbCrN1VqxUfE2uFIc2OJHoPxVPM5BUiKEnQkiA/glSg0QuSV5EUU2p9HuEgYsuvP1dP28DUpov
6rZbbNIIWGFSuTjJFDtKY+2xH7W8sMsq1G8fAvk+W1vvL/oCpQ3QLJJzzgG8a+eanG1llEy6qPfC
iLSqC9C6dC8XYwE4bZwonDBdzO12zkEYBsJVy7L4lOC/Ild7IYbWW7Jmh68WHyy428VjOTnp/iZO
OsArj9/T2sF36AX9kb48SfY+mrB9ix1kx4a0xvn8PLFELooHM0KghMruMimgSXy6oDT90Es2+2Th
OmXlltpUQ80UZalOOhdOI6c95YsZ21AsoZr/FT1WRqm8Bca+gneTx7vmIlG1GHgeHW1CVELDNoYl
UAlPMNGISeg8AknsgbMnh6+b4ATv0tvfnbG+aUGzHpvT4rq5O4yE++AlhIf8CPiWyZnYlDAUlDuQ
ZkRkgEluN5dUuSWFd3z6MVqbDPo+YS+UOzuB/n7L0RKLxQ4cnffVnW6tJVIpONdZAcUq+qAgVHzh
Im8Ty5dWf/GlJeJllPCz3r2/i+glAtZfeIcUf/ti2EQvJSFmI8p/zBq5jRyZXFhfazrb+h5zm1YK
F3YYe1wkVuzYGHKP/wl3dSMMukQvaGRe6yixOYyeZ92mgwVSJZlQwcNov+ohrBsml9ZDUqOGuMht
0d1cBnfb1gl4mBTkIUron/5ri6K+bscfcIGcPqt4PQvTJRAk9DG2QLxgHU/Hurd2zlItYgWs4L+q
fcNqpAeTem88e/Xv8Oz1QRA9lDUUfLvRafmPNghIkD7s7K0Rl5XkCZ3bAqq6zeXDK+Yg/Cb9IyHA
NzcDXWpdtovfg2cJP2GXRmPXPmFzXDunF33jbf8klETYFO08kr8Qq4i8U8hcWGGIrqN3OUUy7tPk
XhPBSWH3r6zggHOnaNw2BkDr04o9JfjfMqWwiUUhtaLgetZ4RBVulZQPsWeITlv3jsBiljO6E2/+
Pbf8vTsDhPPgIU2kx7t3ypp3uzGbeX8rRSqRLjWQxCbcMrNvV1YxMsdHLHId8dpMpIdYmXWF0lRU
uZ1c2ygZOkxA72Plbdd7e1lx3aW4ivQ7+rfe5ePYLY1pTeMk+mrvT5pqjs+xSce45+3LVp/9K7xt
kqk2nU2vv8njiCYzU4jhOnHe1jyr0q5ROD4JOzQuRUcs4NBSpvSUe/wCeLeds/wOT6OMacqyU9xr
vcZhsi4593FRn8F2xRptSxeM4Dq/pi+TS2X5sA0z6VSVDv5a+rY7OliUg/3KGrxjICvU0jOh7gQp
zp330YR37jTygeWsZ1ThuNjVCON9w7ZyWyAEIGN6u48URFGrcJHOLfuaqWKxqp7Ovxt6cgFctMq4
OxfGEybujT4tW68r8F0tEaVnGYuUikakPjgnCjqQIpAgxq0m2w9oB00tgWlp/LAPNYgWI7JFqRY8
TTGZY6zMlXIRUKtyRp1fgXM2LRGHnl2JS7T/MktbPs5vPzP9KM8pQ/v7/ANm/2ns7fjgqwf9cny/
QdDMpNNzb59dFWX6EZxu9SuJ0kFrsvj/1ohcVoBiiIwtXrDx/PhFm+Y6rKti8nZWdHDfldbYxXuz
OsW0tQIqDCQbMu96KksdDATuZS0OmDJzD6or4EgKCFE1GsdvwBXFtKxIgrWVAXusS8wmPseuz4rV
hy59vt+xYDiwd/0Na47mffb/d0OiN1mr2UVmIcz9lotcYJwNa+SUa7GhG/cpCioCiaJXxagEYWzi
GA2o49GUd50Y/dVydInAzK3P4sYDRImyCGogzsXpDtHYu/toHGFLdwd8V+H8RIxBqCCAdLX9hvKB
Uff2Vp9zXAmIJxOVf+vzxS9hphU05vG679VZ8Geo4ln7AUsZHlCBr1NpCkIGWCfjyyLzC5vhwdoJ
mrLDmOYfUs0aAYO5TL+mwMo6TPBIR7uAmpmBA0MFF2CVUnMn5D1Qof7Vwm3sKUwZUJGvtH0fRuGb
67Xe3zEIFiM841LgX8/OYgRW87ZQZ6y1289AdfKPgfUOxyneJgxKR2kqy0BI8RWL3v/Mrwh8csHb
UJEHD0Es1WlRqb2QVTYeX9XxwpLWY7NB9ruUvCIhWpRp8ObGOKnhWSU7UDwUNWEWNqOpzx+r/r3I
u+mdsEznib8ZeswR5W0sTTjaH2E/vBoO1SjARGgmtrl858rne/p70dN32+TD1HaxqFBw/0/VjhvI
5n2u2na5FYYGu5mbsZeLTaQxbGv8NkKO3GdVIIPTS1ruEmzObhs4pUj21zJcvD3h1uzr27qy+DvV
A6fx/jQZb8uQYk1HAPZGZSSkC+B4mgQ27jsh3W12D4b/KwXIbSCpkovcVhfcdhKia+KF81bvxoeY
sSduFtT6d21goGXRbhiR/KoBQFOvM/tK/iw2oEO23ZCDUQbJYcsERm4j8JtXY2FovISIr0YEcjQ5
OT76+wD2QoZAzIHEcCqOM+sooJahPgn8rWz3qlR+cqjDQ7wWZZWPVUz6xLRtjrKJ+NDU8YWWfLj7
rOVSWVSUE72yNIvjo+KUKLmzf5GgOtmMqicgkXFWlEm6vMNmiS64dSsbqrkMYJWS8poXfEN58r96
rvyc9ebXXPyfj6ZTRKteopKBcSfYrSHPmZLB/TeMekgpQFcisdmRnU2yDLrLLMkXGAMm7n23b0rj
1fNrQKjq0dywsHzoVXU9FdB6SEXL7d38oMQqpbues465f4KPfJqB6GQAeEv1WhOOJYsqnZQCbIBz
qrJTi0sB8DdweY4ikJ4vW4tmQHqr1vpWOS0223+rzTrTllbxtromKXDv+yemA3kkNSPQhqJAz5O9
E5JDETvJ1u3MNGNtP76go94N+buL5GkJQ6OtsT7/FmoN6XYoRddFlxVN79Iqfs/xHBxs68kdAgU6
Z1vryYRAC8jJodw0/IxoKgSAeuacIyD+PPRJj2PTn0EAtA9wVQkFxQfA3ktdyKs5Uu8mzFhrHnqd
0XxTSeIJHPC6Opow8VoJOAykDBaJQcZXvEuEbcPQirvPA7z/Ocoo0OZqdcsSe/Gv2HEIuY+fszcN
lRjoziWfHse6QE/Q7vf+MILR2OE4ghN9rake1m7HW5BaxkdkBhuRRfN4Ux3wmvo1yN2GCwHRnqB9
hOXsaVIyTPox3KFWaB/m9QNKPlKa0LXjKk+rMPsRwAjPvdVuYdJ8tAxddt2t09w8tucbgydV3CBB
HmtatCIT50P1EZngNd3cvVd/OtrsXE672VJHqEyyf7PhXmXGvQifuXyJBSXTeNCe0lva2sMa5k9V
kSP0augAljvXwYJQoG343nurL8KkCFReodx13HVXm14UqaVNfp+abzQ3mWN8B0iN2ROKMgAvogOQ
nkEac86Mkc2M7Te56DQVQR8DwsvUUHYibzo6c+UemZLVukb5VOLSkfGZwOWcUxePWuAre75hhjb6
/55DST3g+o5EPx8DSMw6R0JbtizqT8hM9KBX7NZ0e6dkc8zT8VQsoy7IT97SrEqAYyjD7ooEhr8L
YZWTYuYSPZvBt0mO/1BrBWMljMRKcIr4HfpqAWfGEt0y6rAfq0tyN0wpXZtE0tkO9uL8W28SwdwQ
7FLyu7t/I2oagbQ/1RIGmZinkKRnlrGcqiT88MqzFTqSSPR4cNQC3NB+bzsT8yU+wgJbMHdKmZCs
b41BKbcdAjc3uyMKJ26ojyCazHSrla2nLAtWo5POA2WmDdkNKuKyFMVthy7nQdc3MiGmuf2eK0qx
xMLfo0gwuVS1v3YM1jtU7CA/7IapNUU3wAcvls8xJzGE7BWqSKPcfLZsl4dEE2ISy7yuYxGCZSqz
H2EeKnebNgEyxYYYpmkr4lhhk+Yvi3bpmG9rOFfgvtprX/JrMSIHdj/UHIECMO0pc+05XelGBYMm
+XePVMvduiP9jV6wUZO3MCQKNchfNYyKsqlOu/+SRx3XDCucq3/DqiSfq45SCIyzXspCswG8eVgL
8kXDSrBC2WG2CcbZVE9ufSHYtJHrDc8dG6594NySH6HxHU1qWB8cKa91ry360k0pgmrUzkQJYCGU
5QninFbGqUc595RWnu9zhDtjb66k/fQYdKzq1GRrvgkMv/LuFudaTEjhQxLFROain4AnJDPb/cf5
DwvZ1B2IVJQ6TB5f/t+YsjtKY/TztaRLRYK8AGu3CmRzsiffnUhtI9UMibzlGXFvedy3MwHPgiPa
51uZmW+SYn44pZJNmv34TJG36sr/P+2hUiNeXm4cOFgxYl1YrbI6UCWZP53+4TcCrpk/+QuXP3uR
C6L1kHkZCYHQMRZluEc6ZFajkR1MxBFA0M2rUBlQVqmKXzo+kGaWlw7PFVkJOGW5maeumROZKTpP
YzOqdtYQWnRpWSAz0NMgX4xP5/UHIfVBc+z3E99I1vjF22sK9fOqrXBj7sKWl5XNgVR8t9asCKZW
7lnoV9FVNeZ3+ZdJ08JLy56dpBTQF39iqm5Pf/aiUxNrvxJGaqrqpuvHS/4D/DcGenwvDPL5XkGJ
bbNnacqS07lqW5F5t4GPUyQyK03F5yumHd3lKyYDwlS02kHltxzqmzZhCiiGPRx/SvM3NfMM0wLc
86Wp5mo70lc4sGcmnfcdQcqGZXTXD9SjjL5Znn4HmnyFb2F0Zsfkkb9CNDsMl6HO6hC2odnEj8Q/
i6o8IuJeaZpIEuG4741g6OZDBlL+cgT5A0zelLX3Pqu5bx2gifuC0xgQtp6Ye8ThZkl+1oJ5YMzI
Pg9ZiG0Lsf8tJWBqzfN4O9rNwIJPE9lIY12Zu2Ci0ZVm7T/jJwUu+C5okQ+S6kKVpEwgR8ADNOOV
yjqyK488yW95xuZIWwoeJKv69n81kar7e2jN3ip1aPmlS0/8kKEs7teDJEpOrggz/gMAbGzewx/I
7fVWfVuSf+n7JCKeL9uoJ9nElYZSC4106UHmvQebkbUMSiKfilyVjvImsYHQtww0YS/u+qEvAgQZ
14D0IFDyG/y1t3a41WsYUIIYQzJurDVkEOmiAenrC6nUW630YSLkEnXphXt5OIUaOzUrlS2lNggV
Q4g9IyNtvweTIJNmRk6PE6Na8KQyAcQVggR5IqSwBjoMGz5qxIiIy1Mauy5l3dCSRiluHyTmCc75
OcZa8YZrSv8NzJrvbO+sW7B6tFGmKBGYyuLzQbjytBhjBG560dl8lfQ3NZJz62HqZc4uYM5P1sDF
H0Qf2ZnzRsWsN9y783YNDSHb/EdzdaK/RX2OVonznLxcR9El9UJyZR8HMELn1r7CiYz5KSk22845
uBiVQft52fMsXLgMwjpdCzEC9uhgo+9f65CABg9ogUBZtL4Tyj2rexPaUzppi+fetaHfa5wxSHZ9
OupUHDYw8ImSRAshjT61XFAVGhJTKP8SiRer9EbCuK+/8FMuTXj3FtgR3DqhKy/I2Ybwn3i1PjcQ
+bsJo8KNhVA2rCT+O4TV9CKl4nBO8tKYRanK+GQLm53AGfTuKN9F93dHYab8leGWdHL8PWrlV2B+
qEenPLGJHBk2e+MlkAw2Q7xmlvsqyGoNI3llOB5XkbWjX+xugaZ9HvMPsosT90ETdabkl8uZg6xf
o/U4KSL7imhaHBqls2EQAC0jm2YC+wQCAJgf/EVz3b2Fb3Nc4xuYHXPhWFII9bPAC9akGy5ib8oA
nDceKUDOVn6VBkmwKAYexl2Ieoqf7ZZiPU2dSKeAFwQM/RiKnaOEPsUFhk+bGHOR8dFjjCbpSXq1
aUlcizDD9gu43daZLI48x5XUDe3djCkPouuUL88wB5g6JSg9bDoPZ4suSskRwIRP/grrgCf5NbTt
MHdAZXoGBaq6yKkEPQs2sxXIfcnZHd6TfqWYhW462HG1hWUlPa3vIWrxrqyNxvnaB6gVvH+GK30U
D8m816Y1ug82wT75hafMdUQ35CEiFnaAwdBr7FNux4T5+uBNhGANaANjkTe0hJwvQQGxb/MIghly
nLdmgeLbK6tziKYJxd31ApSQD9sz2jkhF4znf75dYIDH8DIteiLojddMdhJjuyGRpz8pLS86+ssY
42sOKOrzmiWFMcLc+vmShOpggxU+ep+DfYS7CG3YW+UD5FWRLsfntsp583/xrNi4xsGZhmlS1RUU
aWKdUXa3nXZ71gEeNiKFTPmAvuVF2+QftHb3kpHxAQY4RoSikKKtiZscEichIo8WY9Abg5zaQcVV
OzsTUaaEZjWt7PD0xGbkMJPVH7KyaBZOhgdHhjcOe4FMigDFLG2OGg4iIhgyq1d5E9OkVfCmN31s
bGvyMQ5JiBy0bEMLBHMg/Yz2MxQ5aaQBQPjWVazKXvSIOvD1rpuRMIDNhcHL3JiWpLDQm4bv6hF/
ye6fZBdcbl47ssjJh5YS5y1t6TGhh6xz3rLMsL4FnxiPAoDJlKudRUp5AcP0JBuvequ5cKsT98TJ
5oavRhLr5WHx/F08ktSmgtjmUqkZevJkPxqwdKXc+oFQ1eBGDtXWRy1hivf4On1wBOLwMM3iNcv7
3JmJqyAzlx5GXAAlj7ve1Dp308o9mHftxkfnr6JnhR3tcnI9NKuEM/vwixryrKBno08jc7SIFd0J
12FERqRSJxQKkjIIzJ0G8LCQRMwNXO4EoSxub21ddIw3Kt/kpRrhL1H4y8VjuykU/jgvLqCgnyQI
Livoj9D3TRQbv1lwaWjfOAQKBWzDX+rA3uXgjQMhYiZYZ8VG0QcgMNaXpC2VA2BOklTCVytNg8wy
4vc3GAWEbk0pVsTYWFo6uI5aZBKJTByv1RWOYc79FuIVE+R5j5MaNiqYVmidbn0p1GkLDTw/17o2
kEWk4ydWdOW/JhnYjv5BoPOCzrQD9o/yHheSgadiMpjqrskvV8orYhZgLCV+5K3sYX4VkS8UQAkx
Qt01ZeCJRzZW45S8p309IJccVZRbscLq5CWfUFp755J5EL5ka75vBoNi3Oy0g6XGIP44bVzkCMYi
/TYBzmYcrcyhdbUEcZv+StrHUbHFikC/wODJxdpKG7I0y9YnS/vFfSxaSXYjWu2HwjGiSOuxbZs9
eSU7dwyzmnbYvkICp32xoAHkP/9/j51EJMFjSiqOUMG9WnsT/v/W3nAq//dn4p4AMucZW50CDk0+
asVJTQnJBbHBd1oo7/AE0oKrIy0XHntHByZE/cBGHMQM2mtRLQnN4dbaRxdE6a/F6G/sp28mKIPW
/UQzo+jVK1tmsjrhFoqyK3A0FroKFP9obqFQh84FPUYbtwjFRp8F9Z9/pFZhylBOSKRomNqA3dtm
4mVHdt+ZzpaxbIKKEy0A/KHZubf3A/Skp2ihVP0fq8plU4NUffZm/QTPv1ZOkx3PhvpAPXIYWIC1
DE4TmyEWfZg+AwhY/J+hHPVTLfLxfAhoXlnLB3q3fRbbZVzoFlXxJgtdqnZoI+AuYslw/AJeF3+b
EEi27bbh61qDdSCSfG9fV2DAjASLwjDr6QTQ0r3WegmF6A9jsZAtXNoJCjBPls9ZjEvk/fsndGNa
3yTLrb3bHlVgDQfN1nX0OwlKjgGfmZTy8byrx+lMr5PM7w+OpkHaBb7msmi1MvPqyjgusacgg3EI
BooGjRFC5AfBg0FPKpGneXPd1SwiR+6w/6kqsTDPDKRyDsR7nuhm3jPJid4is5tmHosbW1o1pbXn
QzuTFzoxoEz1W40MQxZX1wQVDs6uAniHUTnULaCsTL1KSAhkXAZykAFs6fpFhDahALFSibjc7xMw
DxzGJExhtH6ts+XKJd1Jp6flG/nwXYLGU8V7S54yBiLCMmUx2rLRzC/5yzlnopPDK2ATH7qrflhz
m622x7Lm/xC2mm0iWju+P35PnT+/Gs+JEEeqhaLNCY0dYEOSJmt8RxWf1TvLorGa7uqnrh9SNy/u
Y3P4EA038paAHVTdm8xW4FD+Q4ZBAcfM2m3tRvG9o240mn1GW+cx4OZ9lnCnBlHFvev6V7KhaXFC
yxdljt++PVzelCE9r+uhmQ5nKvpEiIvCaZNW4B/wLgjQVGSXhwJgv+abFCfhoERAVGtpxeQn92XR
meU8fXkSxtV3pCs18rVGOjtR08d37sCuobaGsrJfSI4T1o3gbtdhpiIzSFVN6162kKeiFK2+iW29
Kp757YIeO1ietpk1YgL5EnbO79MKdo0/nj7tP+PTfq5M5AiTucQrC4Tiid41sePQUmjlFutnrJdp
FoL+qu/xf/QXMweKdQfRjBNRjlnhUx4O6nwCDEs/CDorOixt1wqGapXb8BVvHch8fcIQLjEwcEMZ
RE7ePHhnIx7+U+VbPSBO1OsETwHzW4ScNGr2VjSrGvxU6IE0VuHCPEkchTbsT8vdx3JhLgBXCi+w
S+KwYBPLeFlgzJg29FT73siVTI0MljNcr6ws6TuKDMXoJ8Ixa6xsaRfwJmv+BGJfhRQIETMAx6f8
Jb1747z1oDxFXCykEJStnw4vcHtiLadeQj27XntCwYM5fYyHexPgSqSOczvg2MQSpAwOpwxcT+U/
j4fS+ZP2+hC6h7fB3q9mLHs7v2K0UtR6a4nAbNHMXNbFJh/cPcXkZ4P03+AxcaByORkPdcQJbpy2
DbnDzhJFJXSpHn192T9IjaNj6TLwvkbQO39F4eLG70BwvrUGENkPssVJN/s3uWCbFfQaCbUWbgse
ro72AAti+YxOH+y9GUZ821ERgNeqILNuhNUS3QdDtG+QkjR9RMhhw0e3UBLP8EPkkrhUURUxG1yu
gyMPGMlE+HguYAwD67HPo498IPu+S3xFWehVS1vxgjsbGFWJUqlFSP6eVZ0zWAWe5Ppct02y/oQ5
yMfGKmlRSjroVXzM2SWI+JF0BAI8Iwd1XI+THGYIZ+TC6g7lrBawua3wyDSQuVvaaRTAiBoVWcIo
HdbXFp1nrCoPH2O788nsg3LPCq2NFGaG1CuFiZiF0mdQnVapWLy2/JHqZNYXfpP3h5bl9qcFmmix
k0PuGEX0vC1l5r4lrkL0yRpxise9IricIlfJbCwy89O0oiZv3FdT3TijA9yV6WaDI5HdhSrnUg7q
tu6be7g/BfDymnPdg/IPiYpCgHDq7Ln48d0MF5pFcJFCvXQLxM5kXmPMhouzZQwDnfoxcOFd+WCR
rzNQUxH9wWrfn4i3by7k/lbjnIq/9Bq7WKlc9uy0sKu9YW2DOExCsgc49qBxTKuhoLSNuq3PXCGO
wtuXiryagiaNZV19yKLUwMKmd7RhdrrXnL1X86roxC8+Qgwv2ldDm5XpLzSO7g2KswAgE2EgQLX6
EGvit1vemBXv4fQ6Th1HyARmJwsVSMpy/FFVwlTKsiNDPonOAxJaAPh5iUlFHxvb3H7aNzZoR2P3
yT31jy6A47veHlvBV8UNsY82I3oaAljYHF0JPkAEGcYJjcTH3kynQVVeJS7vzibj7IeYV9dQKr9r
xegNR91cdy5y6p4ZCoV1ABXcf5wTRTJaCL1zhkSjbJTH+NiaRz5atitNZJRZu0LFnhxXFZH9VRoq
kxWlrt9+d2hktCv+ApUWQ708Gi1TDV62WY7iTo5VnWeUIYcOB599HkQmwcDocRAFlHRn2etre3/a
l6cc0WvZwkmvbKETKxCI/JJsFPYKHLeM3GkkMIG/JPHh1lCltmeXNBt6RHd529EsDlhq3x3jFGA3
uV4SuRxkuw5XqAwt5mP6evLCGfWGIoDp6TtRa4UMPUJxuCJGXJlJ4K96CWFvDF6MnokE0vcs6rer
SN9SpZ/CADnAsVs0dKTi8MX+icLZoVO9L2hO/Wwu9AOKx3Q31xtvsS7yCuTs2viuM0DXQNHnZgmE
OHvA7ni9m/4x97sa65OrcIHAwR5s40ge4at/KEM7k3ykPWecVufj0tzESE+bX9uaUtNNZLtnJXFq
ojfTIByqs3vxKuXEjz/7eCpb+EtCUj9az6MCynnhRVErWMh45PzPvbMgkdfKMK5MpaIASKqRmrzP
7Pa4NUrv4F8CtweiInr0HSrYpr5ELUsTMtvfczFwRCvCW/h82FXHILyodWGW2Rh2e3G3OBNQo0CX
mJgcLJvJHiHolJzID8SvXvntrID6gNoU452U4Yqb/AfPgzQWVciZfMGJvarDHKi+SDK/AMu9xvRD
weGHSBbkZ/O2f8R+5jhmv24oyOU1s0s/UTHugEDLViA4Lou1AbUyYo/SHuaJ2vfRUVAKP/EXA7Oy
tet1RuYPXUQ/TYqacyNcA7ipFouMoWCiDUi/EZhqFSZzUeSUJyuLPlKj2i1zy7Tuq6A5LfAdMqN/
Ssz2sWUxGZqsYLRoNNDbpble+3UGOBEiMcrJPsdrnU/9ZfCvWiSmc4w3/rGZNWISmgT05RtLdjMY
t7//F6NfDZc1FYtMTZGj4+k0uCPENazOLi+7lNmSRWIV7MnM36z/qw3zgCDxCPTSOneBkdioQGSJ
ggpGTcERWIETzvFaiKTETfmpxKjUVbFfkm1C4SvoNSyUhNymo5y3E4ZnTu9BesVA7LXELSRQ5tNA
x+pf5CcbSmFnI+qgb51GeTSXBQqFo1jYf/knsABu11HepTdipGt8M5FdpOrsFaXEWcGFu4ZB3wOi
oehFj16LSOWBgrRNaR0hCA/k6qqeS/6oi8tYG3asuem8HLTxQ7ujKIOd2osngtZHnILOJ5KlGpq2
xyA+sL1mP0bcUTw2hVcGX3yzeRVbU8FyOM0sAWR4Zwp5JPJVo050P95NvcSGt9atp5R+wjeihjGy
lK2f4KxviW8OOOwVKD66CcvsnHYGbm9z6UD45rSQSuKlhLkMYQ5uXTWb0urH82v0xHZK8CcoOYTJ
YqfA/xYdC88R6PvUxtK9H67qIbw4qoK75+xJp3tr4n4YRiHokZ/WUEI9RQQ1nh4hTpcQWoEFO8yj
jTppyisz47o6ewSYeZj5Q2SjDB+GpzEU07V1m78y/JdfpyuFzqGtCQZ5WG3Of1uEpRVEfJhcrkUC
xrTOBoOclwzTFZutHG7RUvp4ERbLxMs/DxPEkNn9as7yHWkipGCmsJ1LSrltV3aohz92c8rfTZdt
jPY8we2jl0y9cHZ4UKpfKfZh1Nu0nHLOoPD0iHk/sU3u6at+ISsKbBLgzuIYQNgSo4yMzzXaHTx9
TkTul4xVTP3lmD8gMKYL1uPpXqHHsxY+HWMUMD84LYjbxe/M58jlQpmva2CQQfxRnfi6NonsN1Ox
sN8DoGHhmYIkY5desZ9LNSiGX/BZD12TlVlKRQ4nuJj4NtKlWcsYbNyBwLgGhVq3rTTzVKLmvVaI
3/A525DuQ5qYJWm2snrg0fBPiuj6Wd4a9Ec+ZcOKm/6xJonl6bCkUC9+fNeE0w0QIILSmIWxScO4
UbA3ieLqclXzM1xXugaawnuyUNaa/aacRo5PbrRpqfObBKfrk9DWr+c5cMZmBpqXnuTenluG8ix+
Av1gXbzv1Rg3rAQn+If06aEbCnF3OHWVIbHYM9H0H8qp473U4pcdHC7sdMeMLZQ3gKGLvPSOqEsh
0mvMhUSNpHYzWU7NH0GlxzA2h2stjRq8v0oGeM8X553W3CPrPL/aOG8fAliOhyrMiHPr8bM5QnDl
jza//OwzT2WMYCo7X7fhOB4PQPkcqNIk2PbnqVGh0rVdVzVbm6rZdgacUMcKdrIzePkNZtxKsKq/
MBWffvhDOIvhV2JdY5QxmROyyYlwtjUsMBEiS6cgDxrLfVoKYzfIR6RY1rNI6dLApqitUTKmvaUY
3ZCr37sUdLwhJR4MP7rpD2eWH+3PPCPWT0L7x6twd2l6F6Dz1W4FMrnjjrrMxqnMitg4NNAtAqvF
PrMBcEMWXiB+j+ahzfbsDbFw5tBaWfEqq9k1Bza0FmBjtTnz8jb6jSa9vsnw11heYVA9NUWJJ086
JcZujwQFU450vwqgEmKBRhXngfXmrj7CSYcMUt6f6YftPSdrrHiCIKwZGwnE0Tcqoc1KQavIEmF3
2hoh49LY8GNtFiMeytHOAeL8tQLzVQdyCUZt7qy00kG5gP+mnsZBxU2P1NbWvHnVJv+/QWCIIUmb
2AZzEVaiQbcZoqAVoU6B0wiCIdWhIqCFi4AeL8CgDw+SAXYGMI/CjoO/kNSHmYCag4hSTgsm0wSP
o85jhiPkkTjHECKuE0fHKwY/cy0i4cnj505dgHW90DpgYsxVt/jYMq86xU+mYmNni/SIklxq3meB
NgDz/GhX5M79TiRQnGxHMp9DtjUl8fP+0nSDiBKiC6Do4TPDpko2gbM2uBBk3uajZEQCKUxWRkRo
ifH8+ZG1RXaRSWvrRm+nxMBfl4ZMaIe5VIojRufw3W/qcWvLhc+5uevNEQ81b9Wn6U9d/ZvB1bbH
xP4wzsluwBw3mjF654f6MCjA46YXJ+JIJPs4mwOavHpi/in7nX8Gsrd2+EbiWzxMfu0QeJqroGtx
Q314wgoaIePlV4hgeOWu87g12fZtcSa46VUms7Vl/+KwwFt904pjE0WIEYDhGxspsW439hoCt2mS
VW+05eySOqzCqN8r9GgS0O8jToM4+A+ZlwHrJuXxlLVk15aZP8BL4crkFq24Cmcq8doeIIh5LhId
HWbOgfPCpa/iOJ5jLwbNC5oR7tbMMXNI6EgKVSW9gseGmnX05ZFGqWCyhL37evW6evwqHDhX8q+J
xFTDl8bnx3IH+HA++QS4Xldk0exdJIF56OIk26Y6PfOcb74XPUU2qItRfbV1Sgy8KYIr58TuqLe/
T2g+bbkbSR/j/wocbSLx5RHKr1OrcZ4RizbE0uZSHc8yQkYvd7rmmxbJDMDn7XfCwiXNTY/t4Ly1
VGVepg1RYYbdfsdsFymLjesGrGSFclri/sm+iDHnfVB/JuS/WCbjZGvio2e6WEJjog+XqrxwQaYu
PVOtG8HTeVCglkrg4y5YWWiVNlcgZID5KRKbvCiRLMT4YfQrlZ4tymY7cUlMQ8k9BIvZV2+93obn
pT00Bk2gNX0dH9u1IRng2+0J/1Vqx0fgDOYL32nYB0ZtcB+LsFKEr2T9lzuXzk02ufrog7hE9HUG
zeBoZCMMP3cLbTB7nfhHoVbh2O1TF6P+2x78kCffoxsfHMZ7wGk/Bmmz9cAn/+frbiTyK5x5bx0i
qNyuVjoU9+5gSQhag1mpogcT2sdsmhjX6XDs89rVVnl5yFNo/pNUG7U6NTJv3Sx918sT4auW5/64
mFoS9fZBHZBJjTS2APxdP4X2Owig8IZrf4hGlaHU7cs6JiiBA1+aiMXsS1Vec4/qxXFjDv6ow46v
EL9pxewDhwDxtuCOYab4RGKy9jhT5df05X2GzQwmWQI9wY9YozIwJzytxEm/nUH7z6jg0MC9HrQ0
iJpmE5G48gxqL9+ndQBgyYQZiuBqSHaTRoU1+LobsLBVkkyYuaHJPkSYW6ujEPb3XWXlNhfjQTSd
7+dr3FiR1B0lCS4wfCG73ZPkZzMmJMwfrWk6k7HKeKYmpAzbxNSyeHii6TcYBgekG76pDAGdjKjo
e3jNcyJs6Njbr1bugHAn7/Ji+c+WFNXiWkwYXJOb425CCeEdKJquDEOXUSViQL2WslU6CYQVDZ3t
7lgsk0H0JUUZpuL08WcMMjpLt4QqIr/xbG33sVIONFBbPsDGB8LbFuttugTYs7a3kZ1MMzsGotxA
v6v4DUx6KBC850gL2G6Ks3/ecndQ/eE/SMMt62F5alwhQoHpinQN0TxIn9driMsILwrnCPYE6NEP
JUToYKfZ+XyhWOgTV4kNeIWFKhwd1JOpjmEQ+cT6YjKg3ApZYl1C3FuQHA1Qpd++y7QQOT6Y/fWx
0r0JvF86v1ji0EP6rXi/AKkmPqgoQDkv3SXEioBW1AaVy2azX2kNt+sVs4Nw01C92kAlMUQNd54E
HAZBB4Xykkr47V9WtAV5r/oQ9nHdbJQjeRnNLBZAhJhcXk/IN8XryZy+7nwDa/7lE4KCcTGuRzdw
nQYQXsZ3jpHDMWquH/QQXr8SOxUDSvp5g9/KvSR7XwDl7Lp0GNn0SLOJzEU8b+qddeFJkxUwdZye
bpTXeNP/ldvDR2hrdG+DGYCdAchAE0ZnXYXQQsNgzkD6uZIDD6T7EPQtmwa4mk/uuYVgch8OJn8G
/cC6lMLnAnwlfaAEXn+CsXap9CtbhJTjMCPdzlfcJXrMFZycIaWBL9T4dJ4d7uq87Z6Zh476rtjd
i/ZWeaJJigi8DTbcP902LtSBWxRxlEtpRWQhb3LjKjr6P2Y3k1YX1nOZToYvm1QCfyXL8pKyntB6
xht8j8EQHRNwbgOfxyrqdkA0GEmfZ6tpcQdIzak2plkDMLFBEI8jQRUEunMdu9V7TSETDQp6zYxd
g/AEW/ljWXVMBjZG0CX74c45LmGibUIWP8pQ/jVwd798SSgYlheZwFFaqJTlsMZNhiJBEn94fCAV
8wuRve98xD7GEhDKRNFrx1MdS7c4dhqYSWW2favGym+t94t6SM31bJlEjMytWAOcuxnUAde7+aPf
XLm5y4/efn/hPqQyW/wnDea6cs1r2hM/csPboPEV0MN6jTINa56Cbkx5LuYDqA0c6RBUW6R0XIRI
s1Hj+rAX+f8kmUg5+OXrNvXYyf8hDgtiTxOBtC2MhllCYk3dWGWWCiIh+VkyaaRPYoOckoQVudZD
wd5XMt0Aw/YhcPLwshh9S2dGlULXMp67uIfut5vfTnFDsSJIkF3F4aUe3wfLlWP00mWxXxAwrm5F
bnJ6kpi0D8nm4XABprgYCkPlhMPGaRmWtQ39DeEZPCxvTzetlksBe6aXKGcBYhLiJ6u3qLFIBqZm
WcJTAUEuQfOoZmM4vy2gxPpgQd1uby6AywsXj6OXgnpMSYG5ygU6TfDEV4+yXDUaBB+VVUVGSwYO
Ct2Gey0x7T/F5hL8H5j5gf61DYDXaGpBroK2cPYha3xxAICNRO/eWijBI0nS6BBfTo2TDEG66UYv
Tfw7uv6fDcVNCIIUxTNiqzD03fSVx+s4tC2CYMQiIvdPPrcZp2XSo8p2Om0JLDpbuCdk7ykKUD/T
hGJaAdZMudpU6+KCshaRgh6vaqTX3wlELCIq2vay/P07sstBiMOgTQDRMkUorxn4HJXBwQtnmD/v
LpNopozaPJRHCAMLxWH6qlxq0K7fxOxHfoz9L22LNmaiCdoSI9gpYYUY7/EX3dMbsXdqMd/SoSIR
Hdqytide8MYan7Ha4u5ZWLNdOiBiG7WlF6dRZ++lkX7SxSwfHpm6r7zmyT600JmPc7fF3OAm5fxI
pr7AoXOPzjC2njsAXlYfUeqzKPleRJwpyg/2txaa54VeeQYzsKWbHvFh7bseEVsbTeZMVqsS2UNJ
Z7l6LgPO0jv23jt0SIgGTXqawOpYpx8m6rAF4rO/qtFrnvI0RmOVnVE1iSPLJxsSfTRWPa4Ba7nm
U4WYoGsPEXm7NslDXlo2mWzqO/cbw/puz4+iFn0OBgJJR+0uTL+4pJixi6bl/fP7aONoKZwwgPIV
0ShlC39cm+eoW9luQ6bUrmJCykC+TUnoXWCG3ZApC16sNxB0cWzS0xrIBXaXtOiLWMhWqzgoUsN4
drjNtbSG3zkp6ZGmWL7cp8TGCYFIF7cH8J3p+6eTBdLc8iLTELGsYFo6ftJLRBWT6cKY1au37Re1
BWvG7m8zp1bYuml89nrGxypQKtaxlUb4H+MI9pq3VRq3W+AO768gpJ3WKyZ9ajnmcdp/a7lkbVYq
DGUt1AgAqmoYteMosAQThz5slsxPwyARpzOkWh5LWBHBrvT7M8BJL2rUtK6lFDCJy1z/SjYPZQZz
gx+ZdP+jjedI4s4Jt/Sy5dxAVig2CRB0LUx83aeoqzoH/J0kVPZ/PUrObcF6zy45fv1GYY1JmXLR
PImkvYewlr/Hy1D7TYVy4vhI7gBBWDhcOBPXFySidagQuETZJ2L1BLZQh7NZgouHKeHnAnbHYhSU
3KkMASCie6RiSclZVopJdjuB+PHy/yZzvNRB1Qp1oYroFrZEixvfiCRVfVnjfnKZ7D//ClmCn+Df
WQtf7ubfsXI+D/Q72wRXySSgdsCs79N5Jb/blHh+Yp/gD90bnN65V1FtU5EM8QPoBqxMgxn3i6fe
wKPLikaUGXVaHt61gxcQKaHc6eaCbxivcaYPnWtM/bv3HAlnP2j1UffzkIuZwM923QKBhf9HI0fM
0kDalcDFws+cdhq5e1JE1gCXhjHpbgiNxNB9/iWO2InimSiJdZuhRdGO8RcQ+6YzzfJGdnHTTdjy
cmH9W8zvwAZ3h6eVtc15j7X5+ebkUDx0KoUOMqAVsEiQtMwbiY4GjFWVZD0YweLi80v9fG3au2aF
bcmOdfjJRu6z8rM2Y+iRLoGVY0QmakFO3fxTCoit5lfAqoWrQq03td+c8/YfFrerx/zCKTbofABt
KhTBv18xH9qMth43TBTLW+K18GjYzbqkimvtqxS/uF8y91SFM4g+/KQtmKQH4IceDz74G3tuaTjO
7Ob7dTak+gRHmIrx3SYwc7Gtq30rX8qu39XXMCXv7ArF1EkC5v1yXabn4bnIOr0WTSmMQLVEtJkB
PoFiY4VpTbSrJ+2yAgTcENNvTXaSKSKgteVE6Rmn2cdXdTVh5JjFfwV9Kp7Wu/m62lannaeIOo9P
ocQFD6W8iUKwgKL9DloJNNSwXQrnrIRPgdBvFPmYP8QHfT6df+mrSjpLUaUVC7rM9j5JwYqOKh1z
8gjnSuKHD8OgiUW9/aNnjqj7VoqAxI3vc+oHNn3l6HFb5BU12QRTpbe/eF7PtYoh/M8tdQN6EZff
TG5uvB+jk4iGiflHImFBbuLAXSIwNYz0fEeUR1LEfs5woQTIJ/pLGIxbE5HY3WU42BmvQGYINJoa
+uKe1TxKROKqbRaahm+cUpt12aI4dwuQTvgcRPfjN8/tkdtQTxENaZuJ0UPT+yBdoBNnjpTlimOF
J6jktXK3cOAqD7CbKTiXf6wFm8b3vWdIE8EXNTSDqKx8vwDz6LRCsraT4OJfDeGVyDSkcJx0cOKf
HnE4sJ8ARzx0lbbyPeLhJSs2C+fAzGcVt4kSqrB0Nzex9XHrL+LbTdce6Kr22gDOhdB1MtK0XZ82
AOtu5gsGuQShHWdTpByZvqIegEpj6/C60XUVJtz6QpYrs75C+KkPNIwSnqioP9sr12zmGUApVJMB
Ju+nwRGoHdyKDbjRxgntUNJdynmgFe6kcT1QlVFWPlHjMjn/yU0x65Vzhb8rYoOQqf7f3MS2gEBa
F70i+OJJIOnPhtm3FvIT7aOdBmeT7A5zajJU/qHqUn86BwmeDDK5S41NWAR0uVFuzixCOMdW6Avm
1cxjh+eGmZdfPggRdBDhj3F3JLu5bJBWSSiNruhPbv+S/i/emruVSXFFKUBSX76JU6MXam4oMpdH
6swk9HDQz2ZMAKuoO+2TKxmX56WFJsNj4P9JGcdkg37UUE9gUSBm/OH55hry+WmEUebQOo2mGbLI
lNzuxK1c7l6h7h3C3wFWdkh8usV/y/h6AYVdetiWvB6mT8kEIA8Ri6wkaSp8TrJ0icCyd+Z5oBxU
B09bxGKQ34bd8wVH7Yw0Ofmz0dPXLrF66hG6LT8dINKTGrDn6fmWEb/Fm0ilmw4Vby561y537pC/
k+26F7MsLEU894izBa+vbb94J5gQ2dLrX1KMnHt/sGx6lWFc+OWF1aMl+TCAzEJix/0cykF7zrUQ
y1PD+9Wa4U7DO4tetXn4ys9wxBRwunECaikn55QpPy3eVb0cXWhkUN2pFpMF9KwHzUCmCFxYHfo6
67JGOCMgc5gMel9TaqyHZ1vNcXdaqMGX2yDp9Mfds8N0FJ42i7dgQqVqB4kHXOj021Tpvb0674Rd
cN+ba2tuT27guvqetD+E+MybXRgNkZ131X1S1HrtKJNG5RwCti7HqH+Ld6JEbZ4rKBsZAL5kaNcA
4jjeamDvr9u+pQT9AGIvgzIT24S+Aj8DPQOybU35SVfRArNcGjiIMrWWWZHSwXpqnhZnFfNQCuXM
Y8xUrCixdt5dtK88aQXyqtJ4gsXTszTB+spZMbUEEqbmMLNKnH2efwtOln2wiQz53TgvGKjIeBvz
orN2LAE9uYcU6ppnCdkvS3gvXmdErb1wp5oT2MC+hMCy1tk7wRbZqOI7W0YYNf9yogRyjFrG2LBC
2k18P+t2fD1afDVfsGrxBElC9i7F9PgMtbD72+BKDjZUR7bvSXBGjQzhJ5fVUwWxNp89+OWcfXTY
IcGyFEVziBFmNfq2O4JeUTlHl6x3Idd0bQoUB3IPbeHjxixHnZO0D0n3tZlbOLw7iCvFK/HYdoIz
NXzkZ02jmttB9SFY98ToGKT06y32Su88M4dILGV3RZO9+BAWtEQOivHyPmMcjRSoWShqvIwDlPLX
cp3KwRt4p9qyfp4CYMwArl2jYYVoTOk5ugGufRG1XuLSw1zKA4rTUJ60m1rHvJ39CPyKmfa8qg4H
VOsGGMsGUrKkA0NVc292OIz3xUglfELFFQDhXQl8FjOLmHGkD8/83kWCgy59o7M3ZrS6HrZ/8KsI
0O3yOFrzz3Wh3n9AftuvAc4eaPNQESzZc3cpsw4xcR8KB4/PTA5Xz+yyp5DEFkqJY4rF5EMIstgG
jXcBpCtZ/DUMukDEvYjrwsVPsrUsSBcmZbfLqr00uXOs30/4bRYGnPd3dyZNRlpxZ0hRvhS9hziD
3xwyBgN+Offq+1j+2xOXTCevUkP/b2Wosnv+vv43FEtSbulYiRP8vc1Ws0oXq65UAkJOUMJrWpjV
tAKl9pdGhDAxuXPBEwJqLmpU9+nDIzULAzw0SvLf+cV9xKXjTjpg8gcq1kZSPue+3roCJ3yFGjA1
Rz/v29Lzw0vZKvJ/C6kKRRdvxvWM5Wu3rwdCfekjlXutRWLqBR75UCN24K9GfGAd44rp8vYwoLjc
TFAZrbXHbEWmVxmzoYyI6+sctn3ydOEBN7FDwbvdSAsrDQYJn9/vqy+mJUu8MniMOpbOovgz+fLa
v50v4JimG1c3m0ntEgcjfJRrFf59a/eU6FqHEFfzPDoKFKWtqjPtZlBMFGCGQD3FulvoSgVzdf1K
EY20YM7JrsbqZztHE5etXCN+gnL7uOgz/2LCKCZuYz9xUELdOYFx2o6UBdwMj5aPrG+Zc1CwwUyQ
csZzRNG/Yccz4XD1T2+mVKSIDg/tTpz3eJVLr5PVtVFNkQXV2y0FR9rIB90TBVuRXkMwBjSKrkJe
vqNW2qUP6b03gZse8L/peG2gBf5z8KwHAtP74DX2rOk1QxiPzdKUTzXSfxA0LxPYi6+z41gr/bhu
W0Hi0zy0l/aqY0UafpDHZc05bcMdCnivoPoUYaBK6FhBfV6pIuCP3qrHUogYVsniaPJjRyJATxBk
Od2VNSeYABqSc2drOMSWQ7+owFbVm3O/Wfok9RiHdmDB8eHHeYAexCQ4yKEXsqW1QZL8WVNiCxWl
mTYrBtcPtycoNKcgZCRyswXNjR8p7RUvfjj6qc20UXiiZDQULVvxGLOnu8dCxHfJzdLSCC8KrDI5
QBh086NVfJmwST5zSJFufV2kCYzhyQmUXZxOKM1VHKpaqBJew0i/qvLbLEE2U1RzXx/Ok8t7PUYU
GRhblir/fR6lcshaQpfvgj84pBDBtJo/WQFrPVnphTE2cQwK4zDOnygaFGxmmosxROWGpx59k67R
CGP7pbLgKhbygwDroNzzwiVGdEmpkAy/HDK8XFKXl2JdszErVy1/LK0tapTKyn9Cy4HdO/ywDEv3
j/fW5sX3QWGU/8LfXbxTZ6FnqxT3gElGQYz/o2uWJXIn3YhY4lfMfzGNK1rHC1m+dly9A3o+UFCg
/TmT2lEf5uEZEECYVD4M738SZqCf8Lr3DfBa2E9rect1pupzws4LYs7+rvifb7ShhHj4z+P94ux4
CpqEoDl5YaA9wGR9bmIboLuGMsSd71Fp1pHIc0T6yQXbLJWZQI3jnkrzGObAJH1YTVzeiYgjWoRd
Yc+Dwdm5D07nf2TieVhqXuTiDO+WAVYnn38ew5rUVrGQqdKfv1CGSx5ng6apHfUwXrfOiHZp5gva
M+HYFSO3apjdTwWD6HChh4Dba+uVnIB82vVoBQJtjGE4Sexc+tqlz0ItYOrG7fKA2M9/WCteEroS
ynJOq+P2NLAudwj0ICnSUpKA0323GhR93X+DEq00s8xZYBUJVhvDQAHIP//ObYX0DeWnUgXCpH69
GUjASN53yO0e+5NgXiT+o4/B7sFVhf2Ll9YFI+7XVhJ5AjlFErfacKoHzwUgRZT8ceczVN7AW5Jn
Hp5sdlqA1hnDs2n1dmMuSll/0IIHmiUnm7b/TbqciLyo/fuwRPbCgHRqp5+ONm+UbJhjXReX665e
jGRD/l5bFvUtWNpVYjy1prAjy587PFb+7Tfv87FKr0dQCBG6Se2aZYAyGHnHeJ3d2s6HVivYd/7C
HHnytqxLP11TOZvPRzlbAcMmOL7+E1k/uqRuOGDv9Ka3FHpOUpX0JjXkxIqjs5REaoEjijtLxgTN
z3U+ZiIYCQayKH/Q6B470Q+tFvBj6lycrOeh4dOIwccmFf/lw9BeN8BPyOHZwbUg8taROGayTmHi
XCD+7Gw7JrZREZfHJmFuH01U3xugO3R7w8anH+1scc+f2ftSklIoTu6l7w7yAWGTomVQ0VjtNtiz
J25kv2/XUL3Yc9C37a74SoV87OVnvOv92nXCi5UdrYqhUtevXqLiaIkJDQjoXja8zhftx2kZtTNp
DJlMp15gbB/VNYT/gDNXb+u7OrpVKDSUjFIMRHEzV8hKwLVod82ZpDpBBB9C3EOh//90rZhscet8
kaRLGLQFB1DBfKiw+9x7zJFv09MN7b2/N1zbM6JgAh80j1/do7ckSPcyt+qzmHPrkCT+OrFSVTJa
Emp1q7nzjSXMt9S6W8XQ05wzvZQdaW5f/m5Yat9msbKwUy6Acq2ckthXF61sOCY5CXXGkuMM5OGx
M/vLdOfH7v1WXp/vsjywkaw2GoUFQsQswg0Lvm2XvBVDevAkO9yIPXiYRDQQjQgXMWI/gxxXhkP5
ZoRuAP9wltosM58VFlqVcNXkoX4488rK+iVu/0pOtmpYAzPNtRuYR281llGGPEXgXxL5gOFgvzSc
ivCLS32tFscgygkMX2W4tawuL5huyiWer56SgAaZKDsak/z4x+0Sl6BgElEyTmefofNs8A84AFv6
Vpvlan5jv9oTxdcrL/jTAqZjo4nop+JUT+JocrHIk6cqQ9hcrI+If64bqf/1vafPJvbHl5AAHCdj
MiA2CBgoRTii3rCqziBkgwf+bPd37o01VKKCai8nSRQmouYCwdTHE4kDC5DFlGSU7YVLeYwCPPXM
MrgxvGULAO3DXf7uyZEYVhIZJzxvavPjkTlHapfHRQIl0yhji44H8Jjwx2aE5F2NsuDogXR6rv3j
ZB6PS0atnz4Hwlp381hhGkH9EpEdnwq+0ovqZar/TiSB5oPMgzi8+BjS2qpG61qOKtyPdV62o2sS
DziqS/RaecZhnVjvC1YIbderXGvWbJswLQGaRaVmG8nvEIbF3+vmbXGvpzwcZuJ+nKM+usON3sg7
cY35pss9v68LvhP8/peMf2uF6RxOsr7s4zhCN/EEWp+hOKJTqwSljqd7Iy77yQ4r57lEpqK9hWhr
hRVsymddjFPI+FlPNa45pkvq60Kdfn992ue0vYcVqINNAd0p1Kiu4ucG77qcTF0CrLrsLVOWlCC0
rLsMTIq0e/MFQKbMwosmvrdMQ+SNBrx6jmQOn+bV3kUT+yUAVcgnYoSapMI+rU1l+L2KH8CjXnkC
gJ4eJ7OckCm5l0NX43NDlqYzIRRFyx48RAl/aor5+knm16ReYxbBSWMsBRV0h0DjYM76iPf/FIoy
6urmZsIXsjpz3soq70NPK53ELI9jcuyzHZFFFi/22NioxMkJ8ZTVzA0YSVr7Frk5c//IxiaMiazJ
TjBYfi2AJ+3U6DQ3mGW6l3sZfpGp59d0k7juj34GenrOixynOcMW0acd3Bj/Tr2vScNgb6wm/fHf
TAXLXqt3jJDuDXJO+36tPxwts6TqfpXqy6fbASttEvRGmDtS8eJ2taZ5Wc0RKw80PAYKHlZqT9GF
6PfdsAlqc/y+2TC6/qmlzUy4oPEwqiaDnJEKwtnoQ2gjR6YxA5G8jPDUaqkfwdzoGleKUv5sZCfX
WNoOpAalJhhhH6P+wOtKztCZ/70XQKc50DGxj0OwaA2UggZm8oXNiwSssWEzowlTGT+v74yK2qpk
z04PpnnSp4YyXFCTgE2fqT+RTRMHwxFGnRA8qZWO7RSCLKy9erte4IK8YrPEei4wcE7vtr59ECcU
zWog1Sp/IUP22MkHC8UsdW5vITzRcdrezHtS9ZRAZqbwh+b6qsZ+j6lz0Yi+is2RtlUtreDLZVh/
iqmA9LMgZIDQea3TDPPKu+wS+Avx76h9bTo8C3bLS0teL0WFkhzG8RYChZKE4g2EfCrBGzGtJNO/
TgCLf+NUDQLtDelLJKkkK+yi4Skc0OaHHCkb4MjpOrLWXiJDT5glZ1fyhE3eVB5SvrA7idB4Qio1
NqinZ3hqCNS6gyvGqBkZYHKmTB1rJuDI4FCvAeUfWVccjaHSFSldGMNy5a/MvkE+9/wV/3v1obN2
khjCUpfpF3/VZjgsgMwrus68hC96xOKAyAnN/B+2SV+zfSHXaUDZN7c9uiHjf5c/UlPZGKBeXuIK
vo1kTGGP5ASDTQbi5hAZoXvDLmXIqqnKXnYQLqMbZ46RUSr5B6ojPLb/cjWNncDxBcaLxUE1Wn32
pQOdfhb06LbzSxWlwcaYenPzyN2GCEnefAt3jUkPjsMRW+F9xwb6i+rtlS5msFgdCKKOJriRm9fz
wLrdi54zZK7eUKBbubRKXrnldk/m2V9of41I+jnwhO0H/PJ+eP2KujO+/TyTsN9/tid0q+wvowOF
PaS795cj42U4EiyH6V+grND4gtx8ne2iW1D8K9tZkro1tt3nyNhyUorHdgdZCweN5hC1e7PgFWzK
jVIaybrVgGpCYZw8ZJw2JjZ/b71kn358eLsaVDfIAmL2vAiMmSn5tbKvu4XRmhzEE0AKUviS+WJ8
bZNeRg3KwNiH7eHr4JdK6IS3n1ehuZrQAhBLw1fDjVnPcSKww1n+h7dAsDI0czzcWcOQqcNmlE4+
HtF+nGdcjT5kOovquCoEYIlX7knKphIq2QoespELElMlH+iYfEY3NOcG9XWLIt+VkAco3fw7J1dU
cQTZ/VkRG3o0vvOMH9JvMRSYWeJJDp2C5IqmFovPP1ovCIEkfnkPQ3zh0+Eg3hNqjjde0cRolLyT
8C1dfYTGVByno/XefW3wu85yKhmYOi0qMuNVcBXkFvqc/QzSyPdaKEy6eYGTLS6QP/aQ7m1s7Fb6
w7mXMwdZuUz67OQG2JspA65Gv80uBULEwZLTrnOA+a8ehADAEDjj4TvYBJZmidNpFloz7vyV71ZT
yK2K1ZsntK/bKOj3gij45TZvykM8Q7QJDvlvbEN7piB9lkX98fuFcMqF9CwldQm3BvcyetjjY28n
xGizSffeEPNlgn57DTFLDebK7SJ/iPhnw5vXFRrp7CDHpNjiYic6CwxnSJyYHCKAp/TtnwQHTKPv
iEzoURXxXDYkDx47Xvj3JckFO5hAyWH42lllPGD13aym4wG8u/TG70FP9vBXI6yJiainL+SSJOEZ
PsyFxxwjMEnUP+3TDEbCk1D5o4LEv3g58Nvpk3a2ZuNNI2IBinhe2o32N/2/L2VpA4k8M5iCMj0g
CCXqDESThli3oU28AHeRpRF6mboM0007+lDW7EZz1M3tQHJQdjUApVIwLPNWSANWIAf2N2g4YjBT
jVUBa4JrSIkz14HJ5tfePamyrFQF2wBDYzuOA8z2Wdy+m0n61smftuydsScmarLDXaL0o75N2gE4
JH9XlYM8fBaO+t1P0GZYPMkNy33eGYdpu3OnHNH24kLrd0IonYoIAyeXk8Mm7RRLEJ8Mk6U9/ozQ
/Cjk5KTwyfgTXE3J20HspdWpAiWuR7h32DtMk9OkkkXCZH0SFxA9V3Rgw5q98suVM4QlcRiK01Xm
WHgMtr2QRsHkhcAl8ThDolsWabWx4DuolDMESepQ7cgociNTeSvfxP/8/ytD1hgUWs8CM5pC2o7l
KoiIWNZ6id5/VD8P2MPeRtyBuwWbKaqqr8QrzBv1NCdK0mWXh3M37sTiSpjVqPTd8Qh5kVqbp3Ko
d8J2MmxN4qOudIJPajy1RvSBWiIeKTvjCf1e6+k/+7Ac74/uXlp1rm0cB77mSOq+G8LRZvGAKNQS
9kNv364TxWL21+ql0SXj2IigYAH9b1wAb3NcBV7siRHeXNegVgIzI4ZYNlrck2AQ2yC5rkBIylcj
bJT15KMUnZLYVZeBfvGtWvpN+BuCr7tpsku94Zji0vCi1wfBIuPvZZlkOkgYkXFaIPblxuWYvYUv
S0bECs1p5LJM/QpaaPc39p+OozPBRvpSyTKcY0uBi+OB0rpqcjOqbq1YQi7h76Dv3+j1X+YmUAHc
yRjHgGUg0obxX2hsgj/u9nNxiK+1HLBxDlxhErla+XzyhB6xq+4rHWTcN926/s2oE6zFA/2P3/Rz
owLe70hRB04+6wMcjA8gtOmsPT61uhZQjLvmKmzzehmV0K/yVlo0VaxgyTcW1ryawVjO15A/iOgH
rdbhiAuKHvMq5NeMnWgrGCLpdfuF/jdQjoY7/pJJR+OjdVIcMOav9ZPZV8NOGauTZXjLJCrGSMId
7g3EYOK/jsfm6wMJdmcaNzLcRA+8SNeX32i93v3ZMXOP6bDj8wgnO457oYO48PSY07soCP9BKF21
XKeHY2+cxl+fC5uvmGlI8uB6HBsB3O8EQUrtBWQT0RFxjJ7vXGIz+w3TWYnkgMPbrR5MrN7dM6dw
FeUm1FzkdLaI297/0z7SYvhSsRL3/D0VwhwzuaSEYC/w9kI5S5nGhye+P5BIVf/zlc5dOUP/WgmO
9qxnb51F1FATAFcABsmoYds4vWJEJaLJus+lDrGXgRmVFaRA+zmZtWTPA5Tz9+prhBxX0SWLFc/K
pjhU0pKdF/wq32m6BAFw7kZgxJSMofNo5cHj1XMbVn7On80d/nyvFN8ocsfwxnl/0O7yJABo/1gH
gp5WIZdWWZHG7s6kRBTdGJVGbjiIhTGKOJRo5VRf7qze01cHtbM83H7c9IkwNg/2JzbbMFKPsVNw
uoPaNWbss3NQD1r1tErmhoOQbZ5++Z1vaGwEtvJ2Aecrzc5Z0xofvtf+ePHGLxoGgCrvrevhZzYJ
ojeyCkQV9WGKMsqE49Y4HfegHs+NDlo2TQGDNwibBlxfCJANeK+7ZHnwllhxXIq7x9baCdBUOPaF
y5+HRcXS/g+UVLRNSzQQoNQQVWxQD3WJP4eD83jLMhsnZUXruEOiC7BTCkgZ30ZkmpRVHm+I+Fbd
ECWSW6+eO89Dd4Mk6rdP8IHNje/mW8dcizk/diV79MVWZHcDUki4zmmwVTneestmAcWteRp7Ro0x
DDfX3Y++cv3kRf84wYgeseUjaBi57lurKQEBr2P1EuF42v/7Y338MUusmW/l1KiFl1pUFhteKnhp
s5n8Cvdd2pVlD97IoO9gehm2f8/CoG0FzsaWPhmCknQAdo20IPLQxqsjexfFWlDhKe3/THp/AtrN
PiR64C7LljWy4B1h9P9q53YbrbHZJTTULZrk4flFqA/wCacrChjrwxohG4hdbgoWYvspXvmrEFdO
LF5qitZQyazVlvKiVImlELxaQco3ky+u2wQbWc1hDeVmQls9Gvp9L/bNDebzH6QVEcWHc6IP8yo3
cY4UXGFTWsHlw8PM6e1JDB5YcbpN4Wc1e5865iqTtExek5Ovb8IjgEaiRJHQ6ZL2JZjPRlQs78UF
i+Pied9we/2Awr1MeEQSdbVL2iSvSW3FBJVb7gSHbMXPggIfUlGxAEjcisavRCBoXwQjmbKhf3jY
azCXYIXgdHKh8C8FgXsJgWk1cr4GYBFNNvDnQP9E0AI9+8py4wS+eRtqSgx6SBlaYRi31oij7NEv
XUJSEuRTQfetqxsu9pG/KWb/eHYeWmP9my4bLFkO9/iYT57uArBcbrEc8nc23CyAAyX0G+Upbprc
swt84BvGk0WW7KuASaHLVqNmTtidyv7VJHn1HLohTMyabjdmvSqNPVEkA5G9FKduM0XaF3fXJW1o
wCUaruP9v6i6KddettII4upd0emgjZ2baYf8pzxxwjYlUS15jp2Ihk74HOwyJk1whzfrt04128lZ
SZcllYoNM8i6fBtorMojd8ssLPVvsT/KeglgRB16O4pZmFeSc0STdioh9vLSWFoo72FERHfKS8M5
7QLpjAGVNMFaTWkDIv615GARYLxVqQRHXt6RtrRcENDcZePoqlZMvz0K43d2115AnWwKzMyZkHJb
tW1XRf+XGInEH8x+jTU7mCKhGFxhmjbORUlQukuKENBemYouUfEsg0P7nL4fwjEJL2i3rXimoda/
0iGcsVRyxIJ6f4OQuRq2Z1xXiQBeszV3exmGlC9MADlRlS1dGiMLzuZyGSQtmBsvXfJHZZ9H8jcs
v2hfynM18XnNUr5OavarjfpVDJ0Ja3v9CkuIjHy+MQiwqYmGpThJ3WdyLd9ZsjHmGv9jw0qpWfNh
HLWhz34qVH3NmeXSZX+xwabuZNRHExI/BXvbAdatwvALtOPvdf1F9bxoAqbylJoVemJCR57Kdq4t
zUWuVOI3D9pe6TtHxHW/ZGX7XMmoNxMrexygY4sHxORwijruB1cCaZpZTMA8YL2yxYmDnZ2jgTMJ
KljlkpPNiff0aTMXtq2vY6tX/TKApcPyqQsjSKJP9TaosFMj14n2O091dUGoQY52gP2PJ56Rnanw
w8ea7iMPK5DVYIzW7HycWGopEC/etmgcdygNxsTykPGiI4eTSjgqKzFE0XJkM6I5yMad4IVjSujY
pEe4jnptfaCF6IKCur7O/41E8TRy+ksEO0rznLX/yJvwJY9nemzWUl1WYh/AsCESbtB9I1+svSkr
Ztx6B3ZRcM80yF1JdNBbHssXxWGorjWiemJGf9LeirSPiNun1BKR/rVKY/78DaMOCroncRCaKsZ8
jQzMy4rJUC1nMlCayPiQBLV4vpzH/WSmcYQNwis1H5DyTa7PiJO/a6GZ4LvrAKlCnIVGUwtYg+8x
7kvG9sdI0QkRJ8EcLls2VXSZqLv7xelE++50zqNQy2NJvGi+bePp78MDv5sdU74zDdny4VZGURHJ
/8xvjFBkYIZzuXQ5594uzO2icr1FvBdBTp3Qr0+r/LdhQjgtHlTJ1v+9ZJCG3Wtr5bldto47651A
72cUIUMPNJlHqYUPGJPI70JWsAU7hVYeuMP5S3r85plrbRSpsOusdnrNTQcegmxxJ9QaEmCHmuAe
zI/AvUwz5pVeacrGgeMt7uuPw8WMFFRoejcUc7lWDN6v+b3kPnKLeAtmu+TG2RWqWIxc1gA3Jul6
Q+gf62A0zdkNUy1MZzB/iJTRMGrsczWTwWHmCoGMMBVCHqpNx3oV/XtIdU4GZsuG6xwsmub4/5vv
yfql/y+LTCkQTyNNSC3PRvWHxDPFGA88fr5yKPs6g8yTh5yiwbyzs5lpALvXPP5cjBpl9EdPkWHs
ju04LlJvVB9FZGIVg5P30Tl0jqXy2HLxtbgXQGWYk1r2I0Hi2mmuQf+ea9Ofw43uYRu5TwB0VahX
k/YMYlPnW7iP/3BqAlv4yo3DCRsN7PCUXt7jfIDC/rqadlY+vLeGhezfTw8r19LL9cjUx1ntDuia
tnwDM7CoHrPOajNb0RtGKNZgZbcgtNOtM68jmYZsb2A7Z9Uagw+YpLsX7FFgODN5wdWcBlJXzgZ+
hVsvWA1AYV/rtfw+TV2o+v45Rcnyvb0Ttajpe4k+7xi7/YlKtAZ22+/m9yJ5si35LZW/t/Grtcnf
2WsvxNS3rdxykQibY3Ljw5ouRlzEScyGNbe/qh8P2QisPc+IYRzZTpvxRHrV8g0VPZLGyqAf1keB
0jMqAKe9Tvae096Cu49YYDrVg6bcXvQ9fwpn31RMdc69Si0kphqi1RnRjUSo20Vjn5WhR0HDsJVy
+J4REG+Uzmib+qRx0Z3B0rWTUgZ+uPiNpCAbziVUlL81tTR8+KeZp9ZUCq+Wr+OENy3z3EbjuUFP
Sj/uqQOm2YtuU7Y4YigLA4ydPrb7NU0NTvKi3+upD0/mdOMVxzczNZtxDSUkwLr7sRFdDaoLogbh
9Gxme7cyUTot7jr4y2gTaBLWiuKwY2SnRvcfrdNYdLopXAUuGGY+I8CF+Yms72dSfqpgTBVyDG7T
UsBGo0OYcOEJzso+QPp9o3XYB6KKJxu7me5vHURpiTYr/rDhHMjSD43oIFNidTBxJY7RWGjKnNOS
eoAMOSs6UvvY97rGpA1Cy+EnHCEk9WEhzVaZ5PN4QcFoit1DvyqUVPxijRvFrWydxbIPvIlsc6RB
sXkukfKz7faA/MURNcXHhcw4y37E6JgHb/aux9S06SPX7/P2wth+Sgr360yfwmLGW3xtrb9tjs7S
cOdtjJ/dGp1TPm86ORZS430ShUikVw5Hh9W3vDtA5YTHP7jwMqIclqaAaMMK2AkkV7T/umW8030W
afUOH/IG64jLubduu35GHLGsTbrI5dVJ8DKV9ryU3yF/MRugr6Pou4WirmomU2sTeJFTZxd7sSB3
xqX8tXcEcg3PglfI8i3ZEuQzDTiU/CYVhffAkO6CjSQv7wconiKSDgapghxzv8s1ARDEH6AKAh0O
3tWC0VIIGmrpA2PB042Lujt6DVxmrb+UTnm6RfA8tQiwIg+DU2yxrdwa8xRdZhyOl15H3owPnRRI
WGaNFmKbXAP7ipxfZKK9VrwfDxtRHDpOYXN1LwYQFhNDlPQ3bDk1w4syr75PlLrFqUU3nxvPUY8c
fGg6asbeIpFEHdOeOWz8QZ+q/5uOCVPA4p08P/9aU+6CmYxQdRaN1rH4Y7HlqwRVDsRXm5A9DYUo
DF6gGjBc+xr5lyJ0Hm+I5M04w0Zmsdawn01PM/FKXCOStqfWqsOMfeFqHiTIGoFq7z8Lxis7cQGC
WO5MIVt2x3m17A51xXkQ5p6YZv52zkRUsnQmIywa3gOAZT2dxTPdj92Mknlc40ze1ksSnX7bDqd8
syEhNjCRw8bl3JjOtsioG42lIP5neXNV5BJ+y+ShibBj7b/92+9Rw5fCrs4t9p+fkgsCzln4jFvo
hMIUCH0W6DpHLBpemETk7t5jKeA7c1n/7RT5eaNZ/sMIVCOdGslKoe9iMnjHPS23+DTciuQ/k1E1
eUsPfi0matdSMa0V414Rb/xj05m5LDCrOVd0TuV3HdpaTsUpRqgzBpOySDlHmyehviN6g+HXKWoJ
SheEY66d+NtAmreEEaF5HfBYpYXb4xp44UoIjh3uYyexdalXiFNqXeg19jsS7Kwu9a/c/YAMO7ND
/KDdrJrygDYd725OGnVIV+218YYG1FpPfHfUJz7/LvJC4WBtqqCNX1VFS0BweR164VsnZDMZEeJr
hdXDfM8z5lV9r5AA5I8qtnovf0dqhkzAyl4pcwQXgfMAaj98mOwMXLJGW5VW11trcivVrDAT1Ltt
mmIHdbGO0FFj3e1ALbDTCwyRP1P0ni9pG/yGthJxXyiXseGji6NZ2+dC/aA6/L1uoWyXYMUU1hQa
UJg7Xc2YgVoHvmIOu++WKcG5S9aT05D+nZtNUVU450jeHvSGXcIz7YTOoiJE7sel9chVRixt+a0b
eBGQjyr0Glb8Lz8u2k+4EQ5Eqh3aGv/c2cjbO7TbWcMmKpElm1xLBoFEfrWGFlzk6PFoKNxqFd2m
aCDPfmbSN0I2QLdXq+9Yt/jDmbVg41iyKJKBO4Gza0JUZzdIYjOcN1qquREoNA7LNELln/mHFKYj
wyvxVPx4qICFJJ+PnjkLrzqV9qMUL/BesD607gaHYHwqN9oUsTPLPaWjoJ1WWtku+z0mtpsfbZQv
/dz/BzRcfYB/0/7VBmsK/QfO7+tDGQC5Aik6N2CihogQ00W1T/BiLGOxHdCSdsbP25LFFWZEcNhQ
md+46arnGZdsCVd+JHj84Q88n+OvMOrNNMIXgEvq1Knd1HmpcvoJ3Dk6fn1AVYKt3pZt9rFJKG3X
/FMc26pUrOAqGSjGLqeKnDe7J1bPX8+MX5WTokfeVH0JIX+mHtsRD8z0TSSvsblcSA8iFH4xl5f6
Ll1GWRlRmi66laxPTRydYg09cz0SSse0LwjQ2dvUaxo+YgClQrRXAYayNQ5VJZIxCoAQD0TnZDGG
ebjxqTMmcN+sFZzBIvg9Q9ol4X3sEDy5UQ6NxgkkX8muRSDmywtd+lGCwM2r08RE8BOLuk8LkNVO
LHekjBMQ1QcdZnsmne2B14NhE9Sxl2hb42zajRsxqGyecQAqXGCllT+IyUdCW0dyjTmaHktuazly
N6UJhL96Ias8JaJXTRsdxTj+oH4jozF6OQJBM6y8/kX23K/B1P7XLxSPOPv/UGs+JC449tO6RLfn
6kgHT8Ylh0l9pbc9yS80t8tppHjlznxsWuqCYAna87PcW0Y6uNFdAKyqDyM+yYJDre3ClBcBURFb
uQtlmYNbhGSyqtQpflMJGHd1aWyHptueWSx8z/syLZ1LOKRBekIV7Kj4NsusSLk7Fpt8WuYxeVbP
ewZ2bfaLWNGiTGe1EV57hsk+bEgM6oG+/64r79+oaUdUje4HsKCksswCfe2K9qI294bB3ojMOq3f
+TSLyGrYPugejXmBFhu8KVo0rIHA1k04KIccshMthQIPoIFjVcAXE3BRc/NmBUBPD2AvVcKV0tKN
NGkR1eN3gO0eiv4J90Ke2aUimDNUpvdna3fYdNFvn5eYiurNabgGB/wW45V4uSdJ2dY7yQtc0VwA
YqvIVCZ1PPfbjHh/8RwE8Y5HiDQsRBBmFkkFhYPplKMZVV0jrYRi/5syJiYTdEedo228n2M0TAUM
1v8zG3bQCnb95J26TNvJLmkaWN/A+JAJXdJNeT2ldbbutsuPKoDv6s61oPJagGnhGNOCGHe7tm1P
mv8nCgGwHu5XyQMVUYeyd9+hiUnP8HN1bqa3gT4Ia+xB8wv+BQubNFaBoVNo7/xIHJME/xNuVg5i
BUoCeYTPB3DSNf/DkpGU2Xn/6AEbQKgvuXVy0OjGkO/5g7ic4aeXD3buyTzbLj843IrP7wU4YVeC
U0P6OLHTLFjnc+wW6O53bTvdkMcnUGTiGJsikW5szOFoU9Ahfp8liigBoz5gHB1zsw2vCACiCZfA
SYPEPQnI5AEw2l1Lv1VnWD+GUO7opGpB8glM1RwyKkZzfBJOO9CbsuWJVsg2E+I2wQB8lBoUGnIl
fe3t+JXuNM3NMz1qVkQv2LGmvYu4KEnntrMChD3ZPUmA+Cf7eaAo6nO7+VjsoaZxCFst7otEEqJR
Ch9gRiajVRsP3Nr9Ymugmh1Nw4LpH8gg26TFZhBCGQ5nOvtIoYaptrmyteg5npXJHLlPwCukixPh
Gcc8dVGj+55OneZ3aA/1urUZS01PrrwzcvtpC5ny3RxRZD1oPj3S6PX8ghvnLNDsTudPaP3XJriW
jI3ry8rFrYeKzudgGwcZz2QT95c03SGnVz92csTsbhYG98qXti7OWfvs+dlO6KROztoi+PTEGfye
MAfOefGdAlQ7IDodZCXncEp9VwA3AUpZAYPnU+car3w/g1pBxA/EJLOM1a47MAXBFC7hGTpF4DAP
JIqcWuCxKbgMcx2dc5Qds44Yam8WHzEnSfD7eXOO4QUPjAKnj408Di3j8NPiw6peYPDGI/2iR2iU
SlYd0X9TGhqpc+oflWzVypsmxsZBZjRFz9UTYKSNBEmMCs96EntpyOg/dnF8rVXdXgQFhXYIV+Ro
PRfEt7hvqMlsN9p2zZiFvsmETR3Fjn4QLRCUgQWQbyYIX3jZBrztfomYMRzFzd7s1s0rPea6/fik
pzrN3DIk4CesYItouxlbo6JgEl1qUj/XmmoS1bgiNGiM8vyIL8tCbAQIuNpbBUUlyvJwesea32Z5
EM96H3V8AYu2CZlB2kyudTNZinegWmBreGX8a4UViU6xoMCEpicmFNDm9IXI6IeuQEs7c9Sep7jp
qLn+pL0JYwrojcE1NzvTkCZoHzM+GLAFtpkSLs3wzOObdhh5jnInyvfZbIhJJZp9MdxQxOg2d8e3
mMY+X7Kgy5IQVn8B7sj4f3IxM37WDXxxpqOkG1c+pURPPPwKSFaQeT7DBONft4fgZwV/rs4ubWXu
AsHnKBF79JClTCEOdo7Y2S26km0ScI6ygA0zZfeFfXTcNZMnACFMlLmd5u4hA5ocXVxAmAa2g3qq
R/6wKE4f2DmSUsbqgEvwkIKb5QJbFdg1oE+DLSEYNZkpBuU6v8PWLqnY76pjE19N2hg502DtHSgH
LReRYvZPfG6TDy5K0sj06GYJLYj1XXneICubOnuwnzRVE2oeZWsYi0Et/Q2j6DBZELw4DRfs43cT
Z+24j81adLYcmiJoIUB8ijtRc/oiZuIgBW0B/yuI4HJoNxaotdhwjy5wPwIkbdJNkdFLt6O8qvmw
slzSM3E2qtQcr2531Bvz9GcYctEgOqznzg7HOXPnw1H1pX/cfIPk6ioitZKMHx4O2R4b1P8J2N6k
Y9JhfJrIemUr0rXLwa2H4lJgGp+ZVHFCd6PtzTQYumrmuba9p9CvRGPkVO/zyGXW3d0z/8151DIV
8nO62rDdLZ/cQEnYSgg463VuQJhlwduh1GHhHy/28YzRdYlKRhIEs85cgAMq9tYOy0AfMyvnrx7j
77C4/FEo6hkT+A5l2/z9E0JB2/VfD1XLdPeatRQS5FXs45ILRK9Tvd6l9uvrX1Jorr+88S3nLz2B
lp1Gii7V+Y5pdoVQDfSH+7z6QC4jq8K35CnceYU9o4a6lVRlfetFHtC7kuSBK7Y3Kx9Vd5InpjLA
v1LpI0WTvH47LPemNsUv740aC83jPLmU4Hcc6huSSRfxUTYFOElmPm3Ex2NJWNN4ZUdlVBO/oiN7
Z9zcm53v1dCqbr5ypeaVAmusGj0pnZg7uAof51mTuBbtScLSPKugkIpzpN8F6RhsdT2PHjeKiM/y
7uTfVIRg599EFD63N9lqg4Sm3CMkwyf9oMPikeVfa/TNhc1CdhzK9SX0xpnB0ZTyzjjNV3XPBcD0
EOZnXx4YEEWn6Qhs1Os1x6TYD+uLMYuMCEZhXQqK16UBONxgJtp3J2kqlaJCu2lNx2xhXkWvzfy2
jw3iRLK2mB98kV36WWL1PTGOBsXDL0koumJJgkdRxzX5Is6jiTtobbb1RAgB6wc3UuiWbEwSvnIY
slhfyG4dTsRrqdnIsyrFJ4+3CkxWx+/tLXSWD1uI5Lgi73pDhvRqJq2uBTUjvUPifNbIzyAmp1tv
Wl6XmulqY+wuVEDVCIGxpaYYUOXA6qWm4mWGebFx6xWUWSTQ+kfrPBo5jM57p9ARBeRc87oz22tK
NXCBOrJYEYgzaL1WsUyt6VCSNmv3pEkHxgrZ+Qmg+FancA588b5Semg3Gr1czrvE3hJALaovj9So
INZ22JaFYPfruxH4DVj0WuEH+EuHEY9qZrVlkSrBGFOecEtFdEAdSyoSkbXxMXb0pH33Qrr3ykYa
Qt5kP19UBe+U+7CTqczoZ+VJPJoiZj8rnKX9tg3AzkimeaBVtVS+FXtaxPP2JJA3MGqFDTm21ZUv
m3Qe2doUCzo/HAzg8UbFpAhfMdrx3aN+YMBXUAvRx7Kyeuf/Rp4S35SSGubuex+DQs9GLK+UWA+t
RAQ7RxCtndQeRmzULPg2HH2nxCZb7hPhqeOS1tX/TOXww2MEEYN0b7dX+d9Bpk9XlNPKmwnwuKup
vJWeF144qbav/OcSsMKDQtlvItq8oassFjtVV3VHUAzVdFhol4aB7V7Zepda8jp340pTFFkGOFd+
9b+JT73ZoaH/l2FjkgXANfmhUkIt1/6nqJmCQX5coVfZl89b7D2+CRKbDGq8V9PxgloBTGtZHruz
9t9+J2u/W5keJhbaeCioD8TCpXeoXPqHU9XaoXczqP92OZnItCQNHqSVxdtYDFjDveIzzbcSo/IQ
OEOIqS5CBFvVRld/F2YTRA1+efaZGcMNJ4W9yi9GIxw3lCikxTjepoFH4fr+xosUCurJnmvlb8Q3
YFu3Fmpw72NUscYYDhDRPKDY9tskg0zaGhJquW+1j+/udAZiEWyI78OQg35whyyBfLdTndHOdAAA
iBPOYPpNSBa2mL8mO0mmY5W+rzSMkDXv5qwQBVxm7+Nt6oUN5L/TKPThCG+QA3j/95KOaS5gnr8M
VIKh834Xopn6aCLBWWv3eAx4qeFQfP2mMS69Q4Fim4nAudT98FdtYFeM/nj0GgexD0ev57U5KKgZ
XS6TQbk/O8Z6079SPzJUEYcsB+z0bU6TL2YhKGWs+YFpXIwuXO0JZ0W1DZ7b6p027ktGS1tVCbM4
ECHGuCc1TaGW/6pFQZ6nPMOxUg9IlPFS6Q0UFjR8JCscTY8A4YMtKS3swP2vpoUD3H9mc+IX+k1Y
SvXIsobKSJwNuRyeQIpe76NpuPZuwq/Gy9rFcIeldGImxV3UJUwwKmAYG3wCUzXRhQZ5Q+vTP16d
BhlYVY3omckbUZLUNHVAZXDX0R92sIB3vjcLpwYS9TgPsapG5tfYIwcUzK4yPBNctIiIfgUpjCnq
Wj0UnxjQWKbH/C9BXUdxqg57b6YY840sJftOBfrm2XCMqlSWZLwpeq0hk2+0TG1AlEoziL6eVb8x
qp81/l4xLZq4XZT+5JccAz6Cmlh7HinZkQg3Jg48gvNtMDzDOU6BGyezb0VEi+IT81nO+HTZSHAD
k+6VynTSPEra98r0EdCB9+hE50QUQoThe+BLDh7or8Zaw9KdbWDwvFw77MPiSYFXDorbin96z4NS
eZaUyBvPiD261J8iK5dabjhf/zkjjnxOPyxQV0keHOYwV1pr+pfHzJX9Bbhu3ZpP+RwiB5XqixN6
WKsKdiPWs3o1o/zngD4t9WqQuaieC4bsNm0CvuzlPyt8rfWHkGoTKSd2Yq9Zl6+wqfzxVzOMKhWC
n++us7zPh90TdSnTm7zc+JEnQUae9GJ+nd9haSgzKOIqS0n6L2gwbn6Rr+QdSf36xtHVLkNaFYsc
EdwJMeI3xsKex2WfQ3GmGF25uTuX/UTBZyyoV1Tr5X+Mmg3KhGihS59vgreK6JPZxPVbdAj2xnLH
uIQpVs3OhIv2jdFrBXCjXiI5naJc7W74QeIgaywAdwvZmRjWrhPkMHMHnWZHqS60R7k23mOECMXv
xiVJtmotzxe834XqNn/BBK4yUuTemXIyPk4p5e2Kt7oKJ9IRsDlrIaFfC7XttQNmqGu/vc6TSeo3
O1iCnUxLHSf9Bff2pC2Xr9RA+TL3F3GNo3cThrqw7ZyXbtBPz6cooByJJOGwxd+YPyZrORMWCdaD
jKN5KYQBQ+W/tXo4DUD8NrVp4CpepT5HZBGzyY2cRdmSxlugdTyMzQcX+4CxI+Vhqu7zVgviuMpE
XhO2ny+us6m2CBUzlovZjF6qqo8rsCD9ATD5nyQAlmyjBCgKWMS6yExbosPYEpK7xcYfFjhDPUDy
GC5HlBmXYa2YSE4dvU9uQgAcDqSvy1eGLUFB1bhBrQBhrBUmY13p0KLI0S5eWdvINjfc9kqdfY3Z
IcCRys3/udr4uG1RkCYs6vN/JrKHNhDLdxUdi6mTJtFxDDsDsdsMimTzqPBN6N+Eqo9An+uNV/mn
K6GCRmTZUDlaoQBkGE4Ti9pbeyGI9WaIASL2AR3KDxmofIbguHZuUmv/Qf2eQWdzk/x5V8b2POO2
COlIcKN1NGfktdozZUvG/sh/PnjkjlMao7qctNHZ0u18Z/Wb2Kq0NelFukM2JzN586Z95qLrfj3W
Zw9QQUQz8NrIH2yiHV8ybpYyYrIQRwIPJhP4Xx0pYwZJfy1+0ob9oQqDaAlEi9Be62VrEMbpl806
6ljiZzJdARFOF+2qOsqdhosQO+x+VD2iaizqfdr04+Se6rnhZvkze0iKC3JcoNVUNyVfy7ZueF3a
8ApbzO+n2wI7Abao446vgW5W2YbKg54/kOnpiHEhGpZGqM6ZXgOJHPyWEfDy6iqrhDnT4bze9iDN
roHcaYjA55nkK4PgYYU/kxw8FojDjjpHndAniMPp62OKwayNDk611uFWYUDXy7jiAyIvZqtNG+5d
MDCXaBeDoz62RDT9m/reQT7jTXfRopcSzXs8j1trKIyv/355AxXeAGLSTMYnQtudxNrmXUDZhpzn
QWq0tQeQd1CpeHhX1fRGr+9Ps5UiJua57vQIad1TRKkQjJgL/LtZJFlwGAj4wtLtK1rTrv8Yw8HD
6x+3VIihxVPYy3PklL5xOcq41Z2it7OWmuLm9GoTtV4WgckZ6EWAe7aa7s6fzgPpli7UFbJ5KKnK
ibIxSA04M75R5uk606M/MwYP7dt5s00PLFaZKPMj2uEhsFAlIvLspDshgSGs5j8kK77I7/W3JehG
LpkOspSfn9CNEq92DCGVgIgRGY2gHaax8WipE1GfDYfOd4qUUfMcuXQN0Q3pn9GgMYER3GRbE3E+
AWf2TysrZ7x2xNIx79gEGt6M3bFJUCu0IoSwZ5hbI2TCT8URcmrhXoRiBqaI8c2+J21tEjDWiCZx
2/kg573Ws5YtEk8RZeTrFhwjhzlfztVilbjaap4y1gAYb3fd7EsyqAsKyyy0G/wPXoglgd6vp8kP
8/9sxlSucwLlk/vywZqymU4VfBw4VeiopZofGRjebBQ95Q/Z1SqjapEpZA6cRGRfGZbDULJ1SY+m
Usv8UFgatMGCeWbd7+h/QlMOsVAtY1aOC9BqyLUvT+VRHToRm1IbKRFZs5JU5tmRwOKSfBCw2Tka
ByO4XZRS1PYaZztgSGRGc3N2yUwUjRICLUYoC1iNSo4inEehHBXb1BnrzIU7+Q6b/imk/KCmtebV
6sh3pz56Ayw+zht38v/+4JAoIRrbigKx3OiAJg4TU+cSS7zKUACQjlcqs/aH4IYoo+uRYL5/y9lU
or6eaHo9JgaE2H/0RaqxiG+RlxOLVvbT/6qcNe2iZqj+n9klkaMUKYKvz3K3SNdDMLkL6MXmSX/M
vMyZKwAJtHDvaEA2aUkHVwOom0cIR5W2KMbWlJtpHPmnKgJihOLnoVBbf+8n6icNytpPdfZefMTT
fWho1Kc112ai7nYW6UfaakpDiQ/Q7OnkVuZ8q3JDO5LJSNmZV5hMH43REWcHNVRnJeM6kIr8fYHK
xbfIFgN2T8KVcM/aZcl6hUjvcxe+fkeqBxoakI3fDY5EMJUDBEcqV2AjO3K014WicrTxshJ41SBx
IzFC/Q27VIeEnGs+ZrGjrCysiIDhy8MxTtF0kfWSMZSFBEX9mXetjKXUu8K6wUPbcqPWHB6oHUPV
E3Iab/U+kLNQg/SPkbC3ddOICBUcXcfPed7CTivM7PsmcLMnAM2rkHosTq7sXMJXZXJx2PsXKwMC
S4sy1nFdONeQz1IIRNWRgTU8+igaqA8LFQvdhn1MjAVZJRxmDzol1sS7i4h75EXJBI3NsfJ17T/r
QDyLJw91XKHd4U1cQozmA0azVeXp4YB6HNPfAXIyUhUnTXjwdUygoGJFnrMw/3e6jRzgLqC+BzG2
Hc1MdKPSVgH/htwUR7pIkO6AMVDDt3dl8hr0J5kCaNSBTB7XCf57VgitX4eGRyQLsNkd9kCoN1eG
AkeHxkl8QkamZdrjHc/H+eB05d4nn0DTp0tJroqZDa1RGBrZGH8uLZ16JBISpnrpbrKFzSQjW8z+
Yjd5kdKEiZJD8ApbuYQIer8rsaSYaeoJFwnWFGSp45tYCH/1teI024/7Ioyj0p/xG24TsM9F8Qp4
oDgcwqsf5bftQ6shTTU3Tl74RaOu4wY1FCCA6RfxPY0dPRXke0UxWoNYfBjspIeeMAZ+BqqN4X+b
nYW06hv2c3k2WZ+zQBOP7ldnYT4BgEmNt6JjP+Crx3gienqOqb6uRLIckrjJuqRLPvcZtBpcQKTu
Y2Q5Ep7V/wTpL7o47AqiwNw3lJARNj9X7WwiR7AAMRZm3ddFuSSNFVbCQW21kMtxTyCUWtdBkCH6
K9g9YQX7vgAmeaLcvphYvgCOI4E3Uxy3Ag2r1hj7Zws86JpjKubkkY63fExNfapLq8YUStOJNptp
LckZBtFSUO0CZGWPS1iu1KPZ4PMmr0hYYQkjO8mlx+RALgcJ35J659D1WlmjJ50vj+5l9uPFBBWp
vb2kciSY2z+F7aVXhj3ftjSyGz14ASeIZ1+MXF9gtJ7eEI6HzFZihvTL9WxWxbQaD9Ztj0mWKbZw
eEusrUYAG+fOsRxBLHKp7Z7+W/EEKlp55i80VOlEUvSNqfZeoAGY22HXsudjplfpiPnhL7WFGKjT
0PV9YYdfrLSVwabnT6o2EELmaBgmp8aRIPSClKyPVRncw6yOkqey8rcXJ3rtSJbJmx11lCzh5oys
pyZsL1TeTsSu74GyFgc3aNtdpfLw1fD6x8lTBWx0+ld78ePmrWaiZdutBivdo//i6my77cl0Bhmw
FKktFeYJPcrchde5iKVEjjFOnjV58LDa/NAF4fWkMPzLvtPkoA2O453Hqx3vNIRK8OpJ+cS07nGQ
tnAzj29wWrqkxDGWy9povcM/rnzLvPu33YJDr0GVRjCVDlmpJgplQ8mfgxj0RyWTygUo+BVugwSw
hR9ZYuCbaD+YfwxQaZd95fEj05S7A+aQIMEvy923TSUSeipd0bhSzza3siikcQ7p/h3Pd1LEZqim
Y4LfgegoIKXvLok/A/yUWvzkD/vRmncFqhchnQVwNlq0f313ZFrNY/6kEa6FpCZAwVGp83brrbru
Nqze/dh41IiQR5UEz1SkUGD5sHlqQYPT6PNhPasPWIkJVPQ8BXMrNOhLKUIEyI+J1CirvDLkJNXi
eVt0deA8CCmG9wFyzsUhcnH7XWL1dTqeZwh0L4V9JPHHEryoUkMQV4+7aYHXqWj1pDlK9otS4Y7Q
1fIUDw3ktOk9/2rVvZ/jY0gS/co42Y870myqlgy2790nuq6LcTaPqtgzSAm8cBccn2sZGlS6239U
+0ZDCJQMC01lW3CrKbZqCDjj4vrwLw7g8rGUyyJjX9+9GyrXpU5zVyzAhlskVgL67JWAnKRaxIBq
qiMwJRN2hmsDPGwzEGSDbPjNRfjODLb6lRO+n/vrdruqB2sqNrTALHbrfSLlipASSoKy8e/TGsmt
8r7tgkBw+ldrJhtyQdDC8bzYVqgzcpjhnogrZOxg/oo9gd2gFdXJnpjNgM6KicSoW+C8WIqgNyef
LgX2IlKGQG/eDh+ABrQ0p9O2eLmoHw8CxIe/IY6p4LWO43wkGdlcoUYC2f23+E2sQpJbTXqlJLDD
Z6AZIm036Gq7ag18oOC6xgk2omfxKfsZ9f+TcovdUCvHfux0TEIPEBbkh7paJN9Pkioqel/i21OA
PBJxfeGDrNurwWM1oTYvqnJfWW5tNwzRkHpSCwdqpQxjIUATR3BxzTgVhGZ1DJFESxREEAIS7rTQ
OqQWgvzl1SXudLVa77EYTlYFQuw/8VK0915VkioVtsxxRtACPld6joMMDHx8woGjHg1Q2q2UCN76
duFsQwwu8EJGLGmYRuIXQG+pbltM6z4s43m7mvo5wKP2R2ZHLEVVxh6JxlSTMQqTVYC0twCPJYCw
pB20IOIunT/U2JReQJ2Iofmd0V3xi3xtHMxAK42eDCBK+fZJ93CSqA0cqr6GpzRcpLNEv+nYDouz
6D4m8z8sLIPyHwEYLYSNtgOlfgXlTqdmGE9Cu6fOkEdMA/rJiONkgTdPj8Vm93KsX1UPCd418b8l
9qawg1u3neeDsbjziUKp+7Usap/dbjk579jM6KwvBr9vOG7wSq4VbO3seaKTg5g0rj7HJhjXAz9N
mrBwoGP7dIy/SplYns/KMlQpOvGv6dNzHfhQW2fIghI/HGCb41NH2eulCOqLBPkrR3DPaNKhGRrt
P4Z5v/DVTvs20T1JTymmSrvl16TNtPMOrNU6N47CIuDxkUSJPc9U0YO8mpUYnc4E4McvXe6fep/K
dYVEvAY+ZWTLf0bqotKAJ0zhiQr7gmQX+r5hN3NlekQDXS2RGM0/0r5V3kFENhy+fb3frVJghw5S
T2IPULMdHGfQEb/AcJWWs8RI6U09MNM2jrdew8bdTh306fJgVapoWEFCupRE0cDBERxg8uel0c6B
neEEQLeHDZmBbBdjcustmwPZc+MRqsWJ5plmFEd/o69KGLXYXEr9jxEd/+yR15YMIhg12oYJ6xe+
Bk8YUIdFgatPY9pwsDevakECeNoFyMmg3qCNpe9oGotF7n5EImAWuAKZ63NAkChN+XPuhuJolIfq
4MYIIP2VOrpwHADRtXF2KXwgFcQdEXvF3vYWV2aixEUmmYy6ayFqCxEKSApsJ/eTBKJbZ1Y4FEsL
WtqdRZlw6VcohroFQsG8bH8x7DTQBM4RzqCSMQwjbIx/GyEmNRM1/XDMTfiQGZK8ltkRAPyjKJk1
A893q2fGeJyoW73EFfeHkA6+Kae6W6acUHtRPyFYX8z/TCMvE3KCf1tE7LjfUYZQgyTNTBBwRIRF
KAxTIlkNcTFIR0OdLa26cjnSwjQ9soMEcv4RAa2fYm/RweTEGawJCtF5G0Clt5AGcdyXKdgAu4bf
iljssffILQfGS18G9dCYuY400QAiX1KVqi8iqnh9rrw3gUkZrM+h9R8hVRJTJWbHi8A2jn1d3DKL
IRBjEUh2cHBynNwnCqXvi6EaN6gJF3i3OQqivGE8B9MdugEJ3lTbWBChn6vHjfRNDobfZ2PUNUub
x7j1OPqJUcSwPhoqQJu0NJ5Z/YkKgDeFwzsIWHkHO/Fr0WLLR4DW2PWQLy4L8bNJ6qGiKnsQyTLL
3+CfweLhGvFLOttqjRicCiIjB4qNEH0HMnYOD+V+uFxIJYfEfL4nhrIkR6v3Xb439A6n8IepgrDK
p/eEaNtA/PhEK5vLAlxrLuEobE4/CEESryB0M4nFWtq31I7ffNRHnVIIW1Mb8qPRBIgM+pDTQU5a
gKleCLw3i5NwxTkAH6eITBdxTVKh1m7GNEsSdUKe8c8tZq72NdLm5dhslk172w7jGO+J6R5M7cto
TPgCfwIwuAlLHO+9+ZiNrGiaefgGvwAcNCHttplb/Mj9dnaC7gMj+hFiKGpOTuN1OH19+IXJtfqf
tWrHA2nnZ7lGoACN8z8E1LtR2coWoBcAhDR80baPhOkAPvq+dCwp4kpgyWub/v3ESdZ/ShVNU8P1
1Ipp2eLhg12i+AKrX0lmR3PbGYMgycDg19naFuVVPwNH5SO5fn5ZJVkEB8kivPmiTYpdT1d42X5V
0fPSRBecb71w+EK3YwqenahACwf0XMKWVFIzrHsRpIs2/krGFHrFQDp7RwCvAoyHKLQb9pKpNyau
jDci9+LlZpAwaacwXDKgpJA3kjM63OVtljZKve/0yzqwqQ27ACkbkA5/HgWfy/CXFsGky9C0Mfjc
vMXBFJfuKc68K8/Npuaih5ouOvqaDzhf27zSRCljB0KqASBz3nCwx6oP+SuzChY/iyT2YMWPnZup
e+BBhWDGGkmhxvXu0kE18IG/jn8OxnpVXHe/FHwIAq1y49ptoGL8cIfgfjJArCiAvFlZg9SEQTWh
ynZgluLesmgz16HFFInn+3bEZciDyGu0eoy11/HsJjtJ7ZqW9aEiEEpe2pWgkJ6ot/BteVNyOzpL
RkaD48pvSSWJ8dg/d55amz21FEL0yR5Ylqg+k0EuPvD5GYfG7xbWNct8fX+Ts+gmmCuFbuZaOfVm
4L5L4xsougtl6usepW9uCG2skuqh3aVMySjndKIPF8s0DsJyWdWDEyiOcO7syDOsDrmSqt/KwT++
xp2J9VskxZ0mx+35LUnXWZyVWSjMO0zeaYfB8BNQN0uand1gHORxN6LE0DATJQtSdQXEkmI5zrMP
O1nTZ4V1aP+3THDzHwWII4dmH0F1WBXTcKgan48tDer+Kv80U4zWSmVPr51N7pX53LHz7lYL/W0A
lvJMnSlqB25ou3jGtgpROAYNyb5MlYe2IPlz10wu41HWl383LhAWqf52Q7qQ6dNdc7vjbHzLp+Yk
yQiWU8CoV5h9PAF37YTsgi6I1U/S/o2O1/+SAevpqXzWAlVsFOovS4Vnb/h9NgS+XJ2NP1KvSqIx
gDtX15Tan6YwbEaj1OdhOgdXFKlR+y4nUNrdCvpxaHJjq9I5sVpf/wEM6D+DYh7hLi4x0E+yoSmk
4e/ZQ/XM7IS/ul12RbxBNbALhD7E7sbHSxAaBbLNACdbJ2jeMA78/lWZVJ+lNjboPFmBR9uaUnu5
qlqBxuge/YdPTgo0i8HNfvh2CcJnQIhza6AqF7aGn5aQAFAqIBo3gaivFVTEAJ7beBZVafXCF6LJ
DlUZK46OMiymj8xOpSs7vkyGa7xyRtXbZ7pysTzCAdXE2hWp123Ej7+EfyFV45n8ESViJnpY9DGq
dUKxKkL7vLqp1UuetS+jZNfyp2bzvJZiHf2oDNVnawzMhmjItnhwsZL1LEO4j8l14+Z/SQHHogpn
/BMUfA5IailrwHDDrC2zBp/X9IQNC8g7TNUwsmnR2Ia5S+iEYxh9FGP1jcqwAfE1sIHC0Aw1R0n1
RhDMv/P4jlf13ynfMxxdMrA1z14Uh/aZgaL0VXoWAPWWEaFKynTMWOQOG4PWM04yVWHk0828To0e
7xhUPtchQwkKVj/VYZIB3YHve7Nfho/miPMOzzmRcyPrhUr0RNzJRHYXAkupx3IsTXsGJW0ztlqL
gXkAzAACckDwZRds0teui+hJXZT0cfWROGnuIyoagUyCgYRMoyUF/JslX7cwppk9cjcIzOvyQo+N
q9dh7gNIoWzwwbCtGwyvm6SPYGF4pculnNeUfaa01dRDMlHIafNG7plqXvqKnpfeG+K9Z4/+a/Md
xc5aO6JQ3pZDngtagXGhwIzkdVTS4BrhQ/1Dzq+YOSvuT3z8O5v8Hy36zDZ7SHDIXIaJlLreZNzU
JibAiE7Qh/b8ftqi0d0LjpBsQtPgPDqPDWQQ44atjIFxbOLGUvKIY+Uj98Dvq5lGm0quEXf/txyN
sD+ju6UaN2gQ5KsArqPgVreU8DX+Lwb1+VLTJzHY5CGbyfKBydhUvCktYb30LOd6/SRX+hP5QtLh
Ko8rOpgYJhx81NvuQlI5pEGL+yoJeVSg5mr9UoLs7kIVWnp/WSaHg70yt6mHWzSuUe1BW/NkHXQ5
0GGMEHWr9cYZdIpXptgRMmvSM7/Jy6zNQcmA5UsnjP3MZpV/NYuw4ydkaLydPfu6z0F2DA9modZb
8Gs3y19mHlJYG0jFWc6QHrVqqqQAo5PtfxtIEKYx0q9yjFE8/jAT5IvSQH9SRbDBsw6Ul1kVZGpT
Dvpl9NoCj4u/xNp79q5lMZQhmgXkQolDepKBUMA6MTRaKq+mgKSPf3i70Gsbkzby/HiGKfKuYZlK
zZb9iYEpdtGic5iw3abqOI1/tq6lM+ehs7Ya3agG84+AivVoUNij4rDNNnldCzEvG3Bg3xnBW6bG
h55w8m8v7tlwPm+AkPuEknBs9vURPi9GlqFWxvJAzKc7jqYGgO+WZbag3n2ZOoPqVRDTReZHI+fm
QS7rMPDKaiN1d9C0f0oC5yNTUMUq7dBd82By7ZIQsRCgbV3p8FauqGYg0KdERAuQR9uELSJHvdUC
K9TfxSyZI4cJaOPlVSm8cA4Tn7Jzrk0d5EsU/AsuPCBxde5FxDnpQBrV2Bn0QBznbxXH6FbItL/7
LrFU8L0CPcVFt7CYVjaSdWTvPs6OQOSWk+uUB8jCt+DXb72c+EhOTLokr4U4LxSdOnainYOSg3/X
/Il/47+1+rVnR6UWfUlF3Vky2FJorl1qpLGLKGEfgEoVkWIDq7+T5iJL60WoazKa7GARVsHQzX1D
x3Sre2aV8WG1ZuxeHCGk05lV6BjLYvcW8PJ8DZFJqN2rVWh801AZCWYZbeMDpg95VnQgRF/C3S+m
1ZZopr+KpxpnSIpMzNtIeHq9rAekOdi56NlN1YC/rPfC6KnOtU6Q/hUl296s9RvG/LDzzxfooPyY
TY6aMOPSfJJVxDJUKZlG2cLHel32sPTu7J1j1UdgWQ1Q+O2yOxQzEHFAqyAJN1/k9ZFAE+Bh3LDy
BVc3FGAQk2xWa0zf4cyuAgDmZ9zvRbg/mRygMtQBZOZiR4UKB56HDedqJdNOookow7eegSuykrT5
/hvRaXRN56PnPNKjCtF5gawDJhi+N1ogUaVVP2AH8wBF9RnTxa3pC8mZrsNFLtTgIOL0YbRksmLo
g6yyzuFrdLM5RHA46Vk9YNK8NjKH81owStLsWqYkWSoY0VQrDxpWsSGyVRIe1v1I+8Sl55jkptSt
dQFEk4s7wTOqpH6dN6xhPmXKbNERh65aC7wKMEivsrT8z1cM/nYQ3PgKxqRxNdiAhOG15h+2K1Fb
gICLAC/HgSQFBi+PrIozikvM3kKcY7AyxVx5OveAwimDWBabOBUsBKLDNpfxMpxgkMftH6o/SIrA
y895hGofQGxPqSRWZaki17kJJmEqVL2kbjJaEW4Rrm20U3eD1qT3ozkZWZOQxfGM3+5jnjqWuM2r
CUheW+Oau+CRgnBZpZxTRHnbNnhrOWoZNPKxV6qxnq0ZnhlVFU6DruJzP7nXCD7Lo0k8K68xDpVP
HvIpLiLnTqB+/5ZmMRV/tJQnBrH/LL8DYXnFCTMU5l1+ZPfRw60mRnQFdIMWrAIiMPTASaYekxao
Q4cIJAB1siGRsTqJdnFJN3Ik/FJGUI3bC7M/GgFEeTCMqBCc+KYHjXpV++6lvZEV8P+ELD54oEha
IV0/SG+9kInh7sTT0ebUKki0TetLbqUv71ToFzk0U0xKu/577lZHXEGA/9cf42hZiKKJx8kg0V3V
dhWyxPLkb0ZzIFqZ4OvDHjpAkDl9j3GEueAqWYjCkknfVDw5QHczjOft43/8OQ3a2LZxyhZVQ1HL
GnWTyx/F94B7eHfp6y8/Tnqp31rklCaM7sgxzAWX90hnUIaEdZJmI3W8EgjdH3gmneT7mwFzD6zD
9DcDAlRSJJS3vIeS5O8ravHYdRzqfXG2VjUfEAAGgJTomdi85KQWydu464SgyWLMAE4XNhgGfsA4
Gt99R0OkaJzIwgdDDzdo1dgf+rWafQrVkJjvZ/Se708HTHN28AZv8kxhNV1WRxKImD65B79wkZI0
I7rs218n7ThqQuJXZVR67DZX7MsIEAisJ5BaHShuJBNeIz6RrlUM9PSWdUjnKHe0fy2po+Ozvinh
1c3Tod77oFMEbAhURZw2Vqtfo+MpFnmajcoqvVYopBSgUe7BgC4qC/BvZ9M4s10JRK8WMwEuiDqu
+A+5MLgUfLg75xhPAKnjpya7HkBTjPoaKJB5o9sQJXAC0Eu0JMT4unw3dYJeWNxS6iKl2//gAABN
6WaXny715gUUY8PlVz3phI5MSgmr3iegM0t9U1x3rjaZXCssYZ/xe9lGQLTPYY/CAeueUWE6TXSu
ZAmi5xSr7CXPAZmRi/WaM9oQiFRplMSlui6DqIOHfYOjizgZMQbQn7itJqP8yLd6RVwn8N8RW0Df
9VmZAIFCYASeqbgERYYXAkSUGibS9hyyboKtAenWoydP4jHYREpDZ1qH9ijKKGlsvAHyycud5kyF
F2glObEkQ/cpaC8LY/lxBQot7s6cCQWJjj+MnI+qvzUNv85EGOC4Eup+A1aOhAFnmdo4O9f4eugo
JS+iqJgSnIvvlDKD3dPuAXaq6FpSN1Iip18sVJCpS5e6LTeaSlxyOd7QHJzD8RCBrXJ9kub1+tQm
FDZN28xQ4ILd8Neuyff2Bml+lEpR4ZZotQbouaoXgZR3qoWDlcElbBTu22m2/S7jYxdvX6ManS+e
raDPrnrkXaQbOTdquDOzcQc+waYjwCAgnev8YUBkpsS7CdoKVkgbz2V41mj7sYeHmULp3cJhK2vL
bhN/+9/Skk9uJBe1/7aaZtHQy55+SO4J9vbWVFBChcPehGDWqUW/9vJOTnozLhS+NVw4n+vdpbmr
ytPzfuptkhcX3Toe0bpcejdPXRksZpzFV6DO6ke1+x7bMWV0rreUXRRwnjK6A6rc6pXM9dhktL9N
xQ2m9AOoA0/l8owT8eezTCCVy1uLsgcudlVYExBgNVFXyBTnb9ZXy2GBGwrGH5YtIcOSjSP+6FE5
XPCm9LZzMhqyYlvPbA+0/O5Gs/5+DHTmDXkfehCYSIL2GWtfi1hJ70OB/cpnROgMwq81YFR1M2ne
gKMlXsKWcKvRTuqLN4urN9+3QTpX7lhaCj8dr63jL9BR+TAlldGxoC2Yc9vHLPYSNyML7/USvmkI
D5hnJhHCNlR6rUd2vq+Vt5b57Pm+3sKRZbyo1w6bagvLWYGAC9Lm85hOwuC+tf/t7AY3Q4J9j4c1
nLlUiTb1PsF+KWUcp1uTctWTgzzohEHw+YRzuCbLhXjU2ZT9mVf42Y2cxxolQjkn63RANv7TK5I9
LMtlVrPmIIgzKyplkE9HdZA+Dr/O+FMSvIRQINAnm9QFzD/treQgBOloQ6xsgGblwgCTYhTnpJCE
yrLcDqW34tYYlijkSq2HOtFaMZKnIKBus1suMaIueGolfrGdfKocZjDPPh8nYdsCXYd1YxyzZniD
gJJPSFP2vfhK/hlkuDN9SuJYxQX4gDVyRFv+w3Dcuk+WtmE+nqjtC5PIXh6Ke2qC0JTxGj8dWbb2
+zuPG693eG7Wj30nOh1+r/xC4IbCB21y0TcMeUQdPnxi3oG0T9oi5G4IZJ9ruA6LZ35tOG0Mt50U
XluLKFayev/qLAjqasCUqOzP+YssLPML6zJV7Wzi29Z0LbIZvMebj45YHqH5w+TI5Lbn86moAywb
9LEopGac1lwbHMHmHWd59kwmwOG8BepuSdnjgW17PPPHVzhkdUCKE4be6cd10eDyxzrUhRLegrMF
xbvCM6u5Wf2MkioAfb4/k+vwp6zeQ2kLeSVRkB+adLM96Nlu74nA/5pXGDxmmSJLTE08ujUzNCw5
U/2A/GRTwVDC9ZBkuE13qqR/wmtKWLyHlFLnd7vvVILAkgeEPNKKcWWIeAQjht2HSoiRStIyqGF+
YyAazfduO6no/Dj15JF1swNKLkDErKcr0VMr2S/dbC5zM1BUNyQW+aVHn5Tn0pE/EBpnbDMRBxi2
0en4cIrMLzv3/wGaWQjv+ggRbXma+je/eFHfBepB84k3AzpfQmky2YA555a6PQDwCcyNchktyeIV
4fLMSz8q6KErN5ajLk5lTcHzt94RyDNs8pBs/HQebNINyHzxYQF4tVOb2cAFkpHzlhFAputBgc+n
aFOUXhbIYo7CVWTRlkTa3yqzlRexmvhctX/79BBA/UYGCzhCa0Gi9r9CZZDE9tUNkUXqLYA32Xsv
KDhdk0ObQNMmPjxYX3Xi1eNSMxbOMJVD1/F69T5Qvb2uDtqh9990lAfs42sfkyUlF1RrxEZxibA2
n7yPUULTLpl65Dqfr3hGcGF8q+CPtGEW6bnpXOj9tNsvECuug13LhyFuwHNANq5IkNGFYtrQSrLL
50WsbY7Rk2LgkGLXnYvQMDpgJJjqCFt+YxXLumNURCXhiLmnlEi5LSTRomy0nDSVbL5RMTjD5oxx
YfbxdQrm4TG/CoekzILlJvSfJkYNumXEwasusyMpyEpX1t3pwxiQENfmyYIQ4rTVpik2rmxIEyIg
JNE2ZHKfFIvqQPSH82O9V9aqt7kKwdBmsxX9X//DUYC22kllfMZAbMeagYa/5KUW21ot3X4T5824
XeiQ3SeTu22d+nJ/+QqErGaGfb24MIZN9B3eMO1/CQt21I6Ds1S+Udqq8lG/5lJXhfwbGNA45iia
xYqa4HlyIcPpExKjUwP71EqPyCTFQXrW/e0B0AI5T8QclYjzUaLyKIPzxmHWM7rMzUqyBdt7bqHF
lPZM/NtGaet1envZjWGyDPnN0mce37Ahf6epFZgXLWcP6GviK+WSjbo/OGEO3peQNxQbYfZJRKC5
lD1wVMdGt3LN431i9XM+//qqep8M0S5O7Er3heYlVD97Y0dhmNvZXUpuGJ5gp+OqcpD0CSbuHdPv
WQDCoNKpBbWR+GENnzpJjKJqTP+tRC17j8kvaWur0JuR+bzNLwmgG0NPH7BnW2qO0G5CivP5CXhf
ALonYLWlFPK2hEVZfpjDYwmW45qDjigxtjE08TYwKODsaFGcNeejpvcJoTT3q93AygV3U09SQR2H
0Xnnr7gfnPhk3lxx5SQA4PNq0PU8Yl4tyKAqL5XAR6L1YDHxwmnVyOOnG+2YL8dyqkHByiNNfk5N
FwpN2RYAGtnSexGM16qDOch0rv4mTw7ojozhHrSU5lkORP1uIfNO6kC0c0V4Nx0bWBoJmJ1p+FWw
G97VtcKcpHZ53MeZE4xiJ8a1JXS701gOQ85YL3pA0+TBqJWu7ofZH5u7XgiiS5T4ZG+QdSYVKTCb
W/IUZuK3YVPWSWp7jC0r7MT8heBK7UKeQjQ074Cl+VqJO4Vofhj0wQRyWI+Ar+MysAHuntEQZO8E
e8Br8jZ7TjbEqJy2ClEQFjwoQApNyrRf0UEbGvYpgvNFWv1KPgg30Kq0S9IAqiFNOfNCb8MEcyZh
grMC343k/VQpmxfFWbYt6s1Rqr4GmV8UkXk0c0ZHNmFSDmXJpr+GG6/Ecql/gKxfZhi0O/RrogeN
1gb2d+U881M32QjNnAC4hmlPrIP1nFxZcn8TEJetyBMqOCpKBk0HDihBoSUqRAmiV0ro9p0QL3eh
aK/rU5vBVaIuNXViBnyFoggg0hIgZ+lLwT0QZwaFy6tXabmNZPXRFfX7bTpo9VxRGdla+oOnUSZq
CoDzdnc59rz88l5vrR1USR9Ke4iaqj6MpgU1tIuZIArzMHohfndmKiwKlTKTLTh1Rvx5BQ2DW0zw
ancUyziJvda5Xm2Wgl/5VxSN0kvAZEFMcZifUSSxKQKAykfJZ4ks4FHCIGdHE1QNIGSuWR6j7BCw
fnhxP5jb9Xk6NcI1qMTynWxnl2c7IivykJto2hsLpWm64u4MuxJSgyvZQ/lw2f7wgKH9WKneySXQ
QpvMZc3TrpXuDfl4Rxn4cH3P3Y1A/wrfj65LVVJIKQtwA+uow1TEosb+KEI2uR3OVNCWjLCh8dex
LHqC++IgHTXxDpPwcRUElvXiQolYmyTVcYhCp0WXRteGekCBRzyEA/akXKpnp494a8tmw8qWBFYd
kT7xdXFFgjNuoIm9R73PDXsqawy3bgTU3vO79NnRf1QGPkWnIiXkZU7nh3m3MzdVbKFknxQBb3uE
RevkBJhzAXRtcQrriKI+mWPM1kA9ACWkeqXXrpmZYGsK5G9s7P81cEKfMDhDXHZN7VeWgYLfP7dU
oTbaiJvSqG0WtgWlemLQYKTxoXgHI7goAfsdmwb47Q0/jpDoGr4siMcsSP8f6N2TXxBBsYYUGhVy
y+v1eyvTO5Pb+jKWtaBM2tqjIzMpjl0Rfp5bzjAogeVOajZ8j7zHTWkO3UdHtNHrFcYV3coq0Cqd
mrSihTDszch5AOgrskb2hF/unaSoqFjEvhtqZKTSC1JRUzSQrtelkOafkkqYSdOj4Tq1kkE9GEa8
lqHufE260RsTXa05Tu9C4K3cFVrx540QWEvPYEdbKBqiMj3TGjzCTqT+mdSCiHSEc+KmYcRsEmIZ
8rGbPGg/MbS1y9ChSpUgoB4xNthAzm8vtbfj73ZL2i9hY7sox0ZOraTcM2WfFf2VKg+WhoQ4zwTq
9622X3P7lvqmvwaZDSwe1iV5/FlyNXTSIMphfrWQbAp/4tCz0YVec3niiZO33Qi4yGizYVwOH1xS
JCI+HGUfZa5/LSfmle55XTMNOlRVuU5fcwh7FKQuR1xAgaciPrYjG0VnyHOysQlVrFU06RONykXt
t62mmi6kdu1wVAZ9hBt76UMXHk9xk1tgUaM/7paMK1g08noCE69/sdnxypnn1wFm3hbyMki9jQBD
8yDV98kFvNHQqHuC3MiuDgTU0zQP830yhQfcuC2nN3z8WF9WmUHu0IfYOzMg+ErNuFhw1kE1TfTA
09keAmrmXiUulSP8FiZf2qOAg7SGQDE8pacUvA9lCvqCnmoKbad+KoR7eJFHEEfi/vpyeFO0DapN
rHP8Cloarruea4D4Eg2zU7zul2M8qoHgJ7IApUwgQIm3bMZ4vi3NFfLIzpj1evKP6VL3+ATSVlQ6
9gkGNzZ4+8/Fl3zntjHSKXnmArXDD3b3QkQL4C+TH6nwfXMEHE1sMT2y2YMkS/QqkdU+RaHa3acO
k/dAVARsGk7LgTLKt372rmLI7YeiMoKD6xLz+0oLi8RYZO4JmuUmQAUzaQqQP9Z8/RfrhIZr64b7
WVnwVSlU98OJo4Dv7nty7oXAzx8OyY2uenr29aj+osBst5ARWvzhvYHmUIN2HWKO+w6IuSK6t8D+
pEfXM62pZUyKptuShz75pI5cq5vCgfOpba0drM5uDOUreK253E2qOt0lMUXA0ihFufG+shQi2ShO
2hJXLXn5iJB1RPWQG6HGfp+pah13y+VI8i3NCEzUko37Nrn5LtIfQo8hwpaFphKyE2HTLEf7SnpU
/1POzNnCRD3zuhI8FYhtBeSB0hI6ADmAjHYSy4vuOEwxsFiNTBnEVOM4giCUm4FPpw7vGJBK3bCU
jAXigYNn/GUWx4BUvePDmgBH1KMQKeGtwTUKmBtutXu8pN2d4k5vHM+CdMRKcr/y3J7Uke/cHPYw
0SjjJ0isC4HFgpdNqJKekPryY+Bvnp5VwXWajTW01a4LuGZGnE1As7TpzP0/NM/TF5jfV8pvc0fj
G3784oWC38aXyIWS427k6ddspHz0lfE1RDAcXJzzsC7OPiSHlzq0Yu1cUxoi1OtZy4HisQk0Ks4B
WFWLpDT0KuX5V2c9Nlv3hhkGXnnJMNBwjme7iUUjQpMbx1TdTJnE4HTVQRm4tMdI55gkWJFBn1y5
5+ywE+JooLm5YMuQmWr0m6Y21YzdVhOQeOasJeKRA3yp5eNun8GoAII2KaL6JfMZ02i1RLscQvSo
Nbnt1KL4nUESTYIx3QmcOfUEQGzIS5ibE6TPNw4QjTrlE0cX0s2UGyE1+NENtWAdqLwI2eHV6Z9m
ijOesTuiv7nPBGUg5IRULcWDqeTJLeZ+LSDrLpeMo6KsQguaINbQGb+HSYh/KASVNoicZ0svZXGj
QZRToaVZ21cgctRf7jg2H9Mv312jWvhD0v2aaE3+K3ui2MG1JfWwNqkMSWaHLFL1sgu4+NuMuPQ3
Vt44T6uhnLa5bnanDP3BKQR+2Svp85jOLB7E3sx61JXQl1Qu6R6+J0KVyt1vT605jW5yHdJfvvIr
RLDtMDR5hC+URMtxhJt+tV/NwQqWdHJYYJWR/4IVxAF4DuK4nnGlaI0IO4oGSqVrJ5hXZZAPcj16
+2fUOSW2Jj8m579xogKJOTW4kGNHQUuz8MJTbQbp/cs4qWKL6+5kxjrLbuRJsnCfzFfuioHX3BcQ
lQC2h42z2zGy0uRV8+S3/LkUymSePFL9cJbvgBcqAlor/VK1FaZbfC3Z0akzH+M94PNF1OODR5Co
DVYSN/wLP3NK5l21FDD8W1zPhTv4WDHK/apKmto6GRW6A27yOlElJUELx3RDcEWyKcp7PsM5J2la
oBD7ymcosGri0iCaC5K3Ip8AjAbzx+//WJBtrx6oOJBWn3GlzIUjUXHtopT6lumGtCgw8WbZQM20
uiiWRA/a2h+FeSm/DF9ErQgcj+sMpEvNsxEyda8tqGi8hUTkY5CeQXSyh5HXsJyABafSHAI6vCTd
RO5OCm2b/DCPdnP1OpBaYmThxvjXhkknk6NbvV0NEo0XAAfCnJujBe+x20Z0H83zGTUDux21f6Az
ItXUg6GZIpijQ7S21FRP2b8HLfSR9jAuWkCaaLMCh3FEVhQsNveTriKiLK54WNwOYcybzrJ7J9k+
GMbzbQZd0b54hBXsCISfCvrq4M6pgtnoB+2UOg9M2kzpV4xXnDhlV2ToTiARWUOT2q2aaNCc7hIn
7j4wvPWYdIdZDKty3PfJF0Sm45j/nTkR/f2ZnS/K98XLuHGUlViuYlverJwTQPsDCct9MPo6tCwg
nRAhUdT+l77s/rAPZlsibZxtZYDUjpdYJptQ5pK27Jda+VQlhcIiUrCEiIcTyN0rtcXa9Zv2lQhb
KL2rosCYzVaqK/aPf2S4zuHSMsm6hQguwGrIvoOUI3E9mueZMPsRsSjZAuZXgO+xJCsUW12RKsyY
u7nK32C9LfKgMUpX+uvtvk8Tsd1aBHHyi2m9Zr+WmGpG3SGSDdl4RDaazimeq+Seo+HQV/vOBo4q
uk30nktF733gjfWLyKx8OsPCg6oeqzCyrE8wVD9sEpLJFMHZSch37xyQgGUASxhtpSFMDNrMwQV5
6fpo8rWWWNuaE6eN6dDwXm9jERBYL7AQy+OmK5KjP5/Fnr5u8o+9yFgqoWA6oi3ev8ASB2ir/AZx
uYhMLQlnMPtZPORt2VDV54U+wJrt1LfpMILZMos+VJvrKrwPayi11zerOpRROkZCMUvYYnsZC0vx
zD+bPjHk81DCmkkDvmUNERj/gC09RorONW23M5XTdASCk6453/pNW3xxeresjSe0czdiY8vpPKj0
qmX5bC9Ei5Ka2zNY5ljK++CjMqN6PCcrf4bj1S5Kk832kPPGIRzYeuABVlUYnelkpqU9jb9f6Znl
rAZs5Ro8L/CXaQXfTUNjoEPjCf6fulC1ZIF/U+Ku9Nb31t4aPdofxNIlzI3N24htNkxtCWN4FZnE
FwX/zQH0rP6SjOUw6L+GL93eQeOdBdRFaVONNU92/FxVz0pdwSH08cU0LmRdVh6Liwlub9TloAll
F1KM/Tl2EHc5/6BvtuD8py8vzJ7/1a3tFrmcGtMQlmcfg1oT9JEB0qc2oFlEC2HG8az2ZipsgOcL
9nh3OG9ss70P9n9aOqM8n4p2Danf0NfZlZ4oD4iJr/8ZbAc7eHb3FIe/cXfFaNZ6AFFtynPnQlhB
Y3HvUvlVJ4ckNT56cLNh6FW41Ott/6EfGRZtIOLuKJvkvf88WxAZ3Eg1X78LN0C3wXN/dmR0XuKD
9dOW3ot50GQlmlrC6wP7Ues5P1zFYB8bL2oYRtPgAHRwbhpkepkccO2rl3eDku7tMoYpZlYGWNbP
WY1ANc0uhbJ4fNi2jZkPXTX6Dr52aPSzDZLeVMi59V9vx4y0uCgr6n6XL3AMDNPg3/VTsDeFBjr3
JYe55soqG1xdADPmMWUigzhms25PQPDNXTJo1UxViR4WpDXi0TpL3XriGazn3RJzSG9niGH8SxTR
/jmfgUR8c5pxnFMUn3Xcb5t/TKBbJesaL4pzVvEiINaEjD+RV9rli1x+KmY4LEutxY1SYNLOaQ40
z+87/Uc0JnAK6P+MAHCKLhOEbaxxZyE5Nj/CummTNz+uldO+yhjpeJ89HYE+fn3DDT46QeP/9pEu
CY3LpOucrIJtpga88XRJgnwkDPdtu8AL4kM5UWKzX6YDWcdGebzMhhASvEyYN2wvGztq/CrKSncV
Kzg3a0Xqq6xkH6Z/xUgVRJA63iC0CmcRi27fHerOlLc4TGYOKQjHVMyeSIwp4k6n33LLkMmGGYB7
h55Y+XqYEGmoNaslMQ6z2zoSjV1YMcfgUzZ6Dz3YKG4DWIpzIXJ+aSxdBJMxSe4mdJfVjZSlAaF7
JVGHwgs5tkjJJsN34B10pu7E4hGzpvfzdMHc2F+Pqy74e0i/HApCckjQfVonMho5vXlkJgXCzOHD
EfmXqjvaWWILzfsLKwZqULo1AtRyiNgl7CUN26UIMtydLy+inm9vKRKFzHWD1uZcpgS3NyadOSiI
6x+cwFAdwCXaFLc5sA4iaZgiZ5r9mwECXoXPsYKq8+g+hHEEKjmjeiaXJ8Oc12HQTBl14iXnaFzt
zD8Ipu3APeet+93Q1O3Irwk7vgWpxDSBJ4EwJI7TE3ISBu/X90/q0DOOa3HDIyFwgU7lsP4NVHVo
UWrnp0ifAd2grxKbcfw0rgik3goTERE1BHx9oCaVPUDK0X8Ff4HpclpMgczxLPzlQNWE1bLEwGNy
SHwE6xRU2Mq7U2iIGHluG+H4aLRHNi/B0pF84Umx1Jtr73ZJ3EEBPPGAepgMtU7gtTM2N6zQDt61
Emh720jbt2Lknyss8BnCblQJ4BfGP2kGoa1MVhPhDTfLQHNKS+p+fFFA3hsnhtr0nfdR3Q057AdX
O4I0Jud46hbkUXQbn8uN5lAORB+wucfaJUEnp5OOGyIVPOXGr/uC5SuANu3zRAd4OrvVd3G840Dc
CSFYeG4TcIixKhRM6/Z8FsCmYdcm65x1hPt8ot6FCcxy7iknQbCwRYeTR2bBLby/T2HqYLPZH362
HT6C3wEjTk9nhF5KeCwzCFq7AG3v5SqFRfFzW1IC0w4CtyKcQy79qQAq8aNPf9+T5QNZ9m2coAaQ
yodNNpm36lIdGYqrmWXS1ZYI3glZLrOqEOzAhs13ZGSP7bW08TX6lgd4GG2w9A6ml0r9q9dTD4xZ
s6g4w9Rtq+tpmjM3KEKdVrZbzHF6CoQMkDsd0muO0oaHVfqh9mnedwxCPubX31s+DVzsOxoKS2EZ
psQ7dodVTD+OEs0r0VrE/t82u/g914eBmPd5s3juYv6ktESSqO2lTN4oVJB90YLjPQqUWJoHMQ6D
AjbnNfmnBWzho2SDfrp/AIJnfBjxA44RdgaoGzBoXByK9wlsTVhSbhpOHZQIOpoVyenhCYKbFRU9
s01KVFDabezE6jZcmtgAfTkO0a0kuj+RrrFZf/Y0Sal61KFy3iIqSoh4+gS3MId+UGGWY+GVDn3P
WAheEvyxj83r92G3mOY0Xgpp82mY0ZOCCz4ILxucqqh+CbGAOQdur2iVTHS0MbFd8rFMzkTi6V+g
Y303M69+lCix8uc5oEJ8dspRTFOiizNE63M2XJvoV3OMD4wo2YNDOCvBumEQUWgSZ2l3LXJ/1NDx
HqBcNSzE+1sX7B7KbQaOcjSQDubw8gd0PT0W1B40YMlpi0C33QPyk5ZfvjDmbyubTTsBp+b62SHt
pMY0EXYcHMygFTLXxvn0mhsnl64p59M7+aB6rbjqVJqHJwiaQir49tRl77W11NHQjKusL6DzFYiv
HvKG8wPQWHs7qE6A4hqThZ0jezcQgQtv3olptz4kV6oSpaSShtTA765f626s3UpXQLz76tUd/idI
JBpMxA9Nt/66QSRpX7p+n/BTFDXGpyfBrIgf/k3++5ysyFpw2RQT+lHZesSisX+46as1sE8K7iWf
XUdXDozEH+ZyaZ4dTolOp+axUNqbIJoXuYwKPm8rAp2FdGxYgPQVLgbIHv2zLCbINCjIvXzjCMu+
ArmYT2i3Xh3MZ5ro2fHdSzMzsfVPuJUSzOYIbCvxAkc8af83s0lJH77SI1dSD5SJC7+vWBruhA94
QGbbtPEVawJ9E+cplvA5/JijrHOVZcZ0G3wDk2MEySVG8andPAGedGRmWXhREc603cQeZBbUTK1r
1cft/XWkY8WEPxc1NFQFdMPfSINS3FTzrzsmNgWoDM97QCU75C4lnVmJeMMJFaDuA6Tzac10qNm3
5vgJh1Gat9wzwYcxqCqsC/U2h0KLNMtlDZPoVcT5F0oe+Yy26T4YLGamrQlhqajjIE5VoGuZv0ha
NwyobUDsAcokrSU0+W+PZYD/1PeSXSHFQVO3xAfwqBf091V18pteGVGwrFnRWPWJRfM6PGN2DyBK
eVkYoLiEsi/cB1ZCDPVnWaAsKjHcjpdqVTH2x+wRgWOh2JgFjVgShq1oCHW+roeKyzATRu84l9+K
mNFHwoCDaT8Nx8GBO5Ua7KXk3KEnU3WQgakm3eMO8wgi1XBhn6bveFGmFdiv9wt+wN3E8R63M9XW
Mm56ZkQNwAbJ5X8+stDlsKgosZdgpXI0VSHzFddeEARpRtvk4pntJI6ILk8f9cfN44OeBXrS9TCt
bh4MfyS0zmlOXyaE/LgM1kosqJuLxUbkTqGnY5m05iQZCGHDIEvW5WFRSYd4pYbIWqFXErGN+ArT
IRhMpn9eGZlI7dJoQZZMxgE/1r+D8tUsBW1Vw2EE03mLGPVt177yyU2ZKw213FIrCgF4gPrujfsN
2ouRgVxv85kZS+mQkacnnEAgK6TbW/5T0OCA13YiN7XfO1vrA72kVXtldsrtaDAgHZ2gXf7VFNNh
+F47mCLukMdjA3V5JnBbYDLIwOpfjtPTDEVl/mI3XZIcUT46LjxplOG34T99kzmqa0Ek9YwbULel
q7bZKXkdAapPaTG3Qhs4E8klvfVpRYNXMvgLPpLjiHuHzvq4ysmuHCn3GNhk1P71ZYTGFsBc2qf5
aANvfKtmxaQCZ4AhuNzkDrYs9IsXEOqoya4pozh90e9PS0SIarVWX7RPVcOmenYy1zof6ybusgGS
w+gC+jlnSTVOU0HWHzMUjJEUzUYZ4AYKOm01u6aHVsO6X66nujQRHWIKzlLH9euRWKnmtqvB5q1Y
Kb0oaiQCzgtSgPjltqp7U6rxE4b4yKQJyq00bYFao7NvAgjS/uX5bUED2p6w2+8T8mFp+lbzS+MI
r834oPN2M/AcojjasG+VcSSDY0dMUhCu2cAAx4wRruQPvczSJ0Ub4dJCcqr3IsO9kurFg5gkJbZU
IzcosX+ic7wuDPvwCt8eorRVS8cgAHn/A1zNZCxD8l14X7+Iz8mS9+v4JmCdyCgglLw7GB9D7A2B
8h0YPGZL5dHRi8GUOToF6rUlVSF9btDzVhkYP+MS3OwewgtEO69M3SswcExRie9qH9t3kM/vvX9I
QdkTQy2Vhh2hehed/6rVZD1/8e1TtJvx/kEuk3csimUDA6hfyj5jc9gxDYKpxXc/1AJyzp/Wfvnd
KEfO8mKp+qk8rb3U3Vpp2Ho4fHizGZ2FmIJoXKt3/LIEIasmyQ0h3JT5wXQfbqXgHk8u4bGZXTjz
iq6QMolEzeLY65/whzFgDSal2luiogWyAB/vmJKww5c7O7NQm68ErDKGe48Ly/97dAdSs/dM30zM
PDgqCVIfEsIL72SrKFPp9XqVOD8XzBwB6FCK7pLTr55x409LOTn26L7Z8dJ4Rkm0t+1IhP6vXgU/
YSo0jfxSIYcv/EZdM9ebDoBXaCbIW8t2rzk4XvmpjYwTCXjqqpg9IRiRdrM2YZ9ZXjEbwPzi7Dgi
43eMp2lXcDhLAlAmiGKFpT8s8D3g0ihWSqXsuxSnhsx74vDH6LTHSTH5KebaO21hDYR4GaBeqvbW
nk1sLqsf5S2ivyzQsK1i6WOSkbzcRI81zKkexiuWZ0KmaLMV4n9S8aF5l+P31yExZ0BX64zVX/63
+OAtT3sADLaRi8SJSYFObSmqdJ1wjJCqKjxI5MKTcK3oQZmxtJ/6innTWGyM230IJgu0q5E4Bfmb
xHlRDQCZFozpVHnqA4juqbzTD7IGAyT+yUBAvxxIYu/pXE12UA5AuKD9UTZbulg1WhJztWQiGThe
X2geAWBJ1roukK3LstUMTAajsWTKGRyufIXjtVkTZC5OTceLPg5PzqCGsXriz/pPmiE0TOJmtqfh
YwefmqzN6jF8CdJ9wOv0PUDpU3z8D6OiHNTlUZZHAMdh5rFy6t6CDB6wRz6PrbyD2mCkLd6cmMK+
+868INdvPC991Lpi9oS29U5PfPCYFyUl9b2ySieQWGuu2t4P8QRqYpf/xO4aNNVUd9OxBKaRZvif
GBcNut163wrxiRxmwmRnQd83AoKiPc5TvOEwWNvowo67EjgblOA1kELZgFERIJI+N7f8hZrcX+KL
a5OEEbH91PPFgN12KBCZJaPDuWrZXh6QC2tM1vb+JX8YH+wMAva+hyJvpEi2+F/S7WOYzrFoBreS
StqhewQfBpAwFho0YNrNhL8ipxEpfnYDPh7ykw7+Knl0ktxDdhy2CjHb5M6+OC26uFc/DqiFoa/5
gegjBC2Yg6/4ji9iZrNr9EkgZTHRK2MKnuLw06NERBE0opu4FGi02HFl2+mW3DKhOnBmejmydHi4
bqeXHd/+hB5LcO/lRtkqhsCHJTJpk0vf+lpUQtRB6YN9rmGG/MTV93Kf36PGP0XXb6OgtZDhrBYf
Up+7BnlT4bUTi+UtcgX/BnaEgysaL4xtB9RF+QmlrjkWAnvhOSOW6qtTp/+pJ7rOpF0vUfvF1ukb
PkONR+mC3jBWy2yeroRH0VSOBPEHLZIhTKImdZVuZzEpG8iEDtN2fw504bP5m94vIOH2Tl75nUVv
WFuFy2kuEy8kAyVPDi55DsWsZE8ZyCjYju+zMJR6BXNAkO57iDBj6OkOtQjgyzbaQbxvim2IgPTW
YlSYgJLNmMvuSwPMvkpprkW+hZ2jJT4x9ZR/rm+PysUz/bpHA5bD9X5nWBRCZMapfuOi1m+m9KHB
k4atqyyXEvJhe1tCt3s3oRQajFNHZ/pVSmjF9JXTGC8pC0GNwXeQAU6exKJjR2SXrD3cbc3HhwAA
95TtqCw2iuEka5v/QWIT3EV3IsOLVq1cQr1rNv3MDALQ2XNAJqNEg40kjhZNcj3/tiHm80iLPy66
Lm2TP3tZUD3zRtt5lByF/kyAis5zv9hean7ABCUNwKVu3PPWqXa7qLK1o0xC8QFN4Qxh5UKghpeG
M0FxcKfN28bKKPPdNel2QkBnbEPovSV6Y/lFL70/2Kb7kSMKnluZr5UOvTYOyi/wQgaylEcUeqve
PAApuD54wgNRIc3f4zdGxvd49b4+EUy6jy/3zazysf+Ab7iXEzfTx40iwTUmo3/nVmn5IjUoV2kN
1bx/7SpOPuDaEQHW/5YXLTdH8UkEzWTDrvlquJ+jTQRMn5SysvYZC8pZ+dBHu3BZMKbcSfQpdd7Z
CX04dtT4fIQvIUkque+uXdc1hG1ihzbGDSBpZxtocyt/QLcHpPuBNRjhLe07UO5zNET+qEnNjEvo
IiCcEmXag6QKvsSQhfJAyf3JYhINF/aUG8Svik0zjpXhwdJ7qG6f8u/3t/BQuOhzGnizFm8UdLI3
152he/EJW2vViojGU1MAypsRZHNQUdbbsJdf8nmZxBlHQOqvyZScZ6GKd+nG1knFqdr0HP9BEldp
Ux1m5kIw0+Y/r1lBZI4ES+2AiCraVbSGH3DjAFKcJj48xs2EWdmm7nRvtiyBKDFRJelWORc8njfj
sMjc3Yb8cnD1w8Wq1XhAxxg/j4V72taFxuTX+ITiGKxGDRaCi6a3lZ6eL2zW7DmZ2IICPNxajcmb
HtBSvjoRDetgetDOAWJLx2P/upe1Nu3X5b0M1xYi6ZrvYqYJycB5VXFUaPRidSWVmvxVVPBQ4r78
vtcMHpr0CADKqIbhF4FteHIM9Ez7wPPwGQL585gjgLPwISvsB7vSixG2GOtvXtA5DIVOfJ8Ls2JP
f5vrVlaj6m2usBL4SPJWZiYxNYL/TSGZKYQQBA9KpweeFCzGmetCwGY9SasRkfQkKYYuFMRpZsXE
Xc6mv0PdzU7mmfNCTbnqNxP59IU6ByAlEkEOUMDabu2G7k72TVWGso8QaQFaN0ZR012IhzEUVohw
IJNKlTyABVB1OYbD7xZvovkhfkc193DhsNpnDnm1FIKVn5Mj6ErQUjm9yL+KUgUFAv4XnsghruvK
ksuBt1txtlQhzOe1zHEmvnKSR3G5iChdKKXd85InVtmcud6C4Wo88YeCc1Qhkk0ljeiHDTPDipmr
2q0gKtgZ3BojD6o9n55NHgtleo2BMy+p/DnLFJwcw9rC1kPAkR9NE5FETkTLy/IlkQrwnysxmXn7
FRXzqd5T9PJdFKtdrTf98HZ0haPwq4YANWlWZAEHISez422IppsVFFX4un0nGTNt2GOtTJ4lQcmP
IwQ+r491U29cn2g4/mBDNcvIZO4jypbTDei6ja62WWa2gvpNpNgNkcYFhuVBmLH4EqBzSia9rzYR
pAN/fhEvP09usht6jIUZKR8DOujkdfOcFeAmuNFcDbM1nQq43sASNOAd8J7mXnfrHEMso2s244T9
GinXycgpM+h5YmL37XII7nCBVax1V8iyA3wrXBL5ABNNJUBg5xlCvgpQTXuGugdSIDJR0UQQnYyj
pCcXXUVWEt9sxsCp+CfD/54EQzvAKr/RokySMF2J/W1rqypjHe7Fg1+ZioZplzxbeGxlYQnZZrHy
Y4E+b+AQbWM/cleUoCiLr/r7qW9xaX77tEktvh1Ls80VoIQw/wiyIH/AUU3aoE0Y4AM5yuKqVymF
dphlOc47g1AibI6v+AY4HQ0nGehqxm1qkAXWRIblr5RUnme6kNGccRAt8D2n7sh7TrGwTzi7/Y1z
LdVJx03SnkjDtyMJWIACGBwvvatm3LbKqdl6fZOaCFLm+c4zSXUCc8nH5TAnrgMFovTnacxJYfZg
N80uI3hU13mR6qhI4MkJJB2ghrJIv1Q4FW+DpxVO+5qyq/VvzUBooSQHy17H+IjH82YFAEqnEwln
rcQfIv4slp4vf3B19d2HwAbzzs05KuXtRHzL3FQ/XbUFDwEp72h3zi/Kv60Bsl6svxeBQbkD/Q3c
nBJvt6Q7AXe0VQP3QsZTN/2n661+ozhQICCtSbzgYYNfqGhaoJ8avhriVVD7yVP0pJ9KT2zfll9o
vDU4Z0VxD1XZg1w/mRnvCwihOtYQ9Lsz14u4A+l6dSx6E7JjPIBxuG5DUBuDMPMpoM5fZBtIwP0f
iFf2Zw9fZEhwhDd0Zqe9iiPCkhKR3DdSt8ScyAD0MvNQdOWxEqwYtqPtvEdpY4IxxY9rQeYNdwuB
mU6ZcocmDqeA/j5sPammr0oM3mTxzLkHoowJdfkY2MFL8eAXYrz5pNFgHwicbfbGzHyRdNPLzuh8
Qmd87QH245xP1cJcmD599Cd1sjrVhWL3GG309Lkeb3gjXGKPbF6kepV6xJY/iJNbipGKcc5uHfM2
NFNZcQJ4npU9PbXhY+SDzwPfRrOcI6NstUqSmtXm0+C5Iblb9BVoRSqDOdbBLoDdvHSxHtlTr8j2
5tuFn5uKv8/C2TO4pAqgpP+TMPdYVVrCIrqwV1RBzxwh2sPLxPnRs78WqYexVB9/r1SSvHnmzeH9
1rceP5u/45OkHCoMfCx1XPofFimv4L5PM7mJXJpsrH8gCZ7qIqU/1Dz5ODs9Tu0oRYAk6JRvpXyX
AwLcEOrdu1GLi6OxAHl6ImgJRpuY524xe8MtrR8wCHNfDEc4fTQIdrlRIl24teoQBP5N7kEHFgqm
/wqeLFhm6PShpHs5h1/V6unlcbh8wuEaWWqtc4lWoRpzG/h/dbtA4ue8Zy6/dZiyh4C2JHKLzxDn
XzV53gxQH/P90L87JHGHL9VXB4it9vty9VpIi/r5VyM4HP6MNNugTvTOzA3DEj1e2pu1bJ5vo6Fw
zxWoH1exzoTJnad9TL8V5CBYAyZcpVTZz/A64U+7sc0bjzSLf1WXi2P+7LhOo1MeRK9VGFxv+PsP
hs3WPa0tuTr31meBghyHKDObevoe9FtNyN42vk39v1HgY32IAnby20Dr2gsR/5smlmj0FtV0TakI
p4w4/yqJkstPCKrP0p+sTk1Fhve4bzdxE3N/jXYfChbxwSErGcVoJssck0YLuZa2RiZbt8Dtm+Nu
gXDtmDhHQ9z8bHcqeGji7xHREfLLHnpQXEzZPP8Z2sPd+H0CLEU8W2474dJ/yKMuNFtnR+yZlKJB
A0wU9H23pP+B8nvyoBSVaB/mrHbdWAKzLdTRNq0qqsmz/dO61NtNZnn9GLf+y1WWKulvvUrxD4bW
qC1aKlVr4JlN7UzfV53s4//N/GarBiptyL6BHZHq6talLvcVnxvi1bEiHxK8Kyyz76mKiCjCp0q1
/Ouqj7F79RzdFoMSNnz/uOHdH31p5Ae/NbtmE6NBdfVTdt47VWcqzFGQ/IvtgmfFprBb/r860Z/G
9mwYRu2D9vV++ea9HBntgIHaw9g+PzqfwWylp1BtYbOO5WZQyTOWtvMtWWVBX3QMftiCoeQ/hGxP
qtwi6Eiw+JFOwsOROHU+WJA2BaBeVpF8RFlcmF7uVYuVaAU/SSHHW6E2oFhlH5K5I9wRnsgEE26X
dw4rvEk+b5/Bk7KakAsK6d9vL91DZJkWbSEqdbhJn9Uk8ltGTq+yEvqSOdZPeaBXi/nw0vxfpkg9
a/p22yH1vGvxSeXE0gSPVw5wuqQSws0T7fu2etkVy6Bs1soG9OOMCVNDbB3zIMDq+j//LfLd1EYx
w45wEJVoe6LBO4/OvujlModU4MhMdfUfldIODgFWVI4xZ5QKlE1P96iwspvYf9k4TkZSj6Sq7mKt
BpRAIfB5Y3EPNcZuWlp0wFJ6qz9kulKKtREUaCItY1YyIazYq/hk/2zjZyZGrCDQR30ROrfi8rWu
FVACHQNRUwJyS8HNSlTgK7wSmfPf+I81pYTEaLLCDQjFrJTiTF/6x89ReG34nC2pKoqOKc8iz7Xr
O55xFBZYHs0A10xrIIUY1ovZ5skDF3ytRjbo4GpTwxZyI5n5Z2kaJsYs3mB7huVcQcDlI2ZVypxW
AUktjqSTNFdCeyvL5v2gkH9wFHCPdnkpnjdURWiJMcKm59YuOf/28SVP85Rj58VJYvI0Z4YHcODB
6On5/GnB9GUZySY/fCj4XnB9T6bATOSpjBdwrlNtM2swZyk1VBknbqBEFuqB4CmA1mgZp8O82Zeo
Su1JFbQeyXQik4DEZFyZuzaCoDRtQyS/+53uVFZGK5GWpu49w66dC35DIxivS7xVsyjrtsPnToug
GrcGoVOwWSKFtKosk3icBBzkcZpOnpyEBM6qVHzwFO8oqads7wpWXkFk6hyFnyAJK2y/yPK0UE1d
3r1MvRfqCCpRya+KAQSpuOSlE8oSFqCF4oPYWmBl6ps2VxqgsY0142VGsJXqbrTGgTEmcxaQE/Di
eNdqV3uDRWD/+l7JDlIM/gDd1CWxhMnIZ/LCyfGT8Rg2BKf2aqI9q7reoZI9Rz9L1GChiGdQTtwO
GYecz8WICmQVTeQM6wh1N5ALMH8hfpMbPp3NKZJXjgnqUXjNVaKkzxyr4C1LxiPjI4sEwx8aKfG1
+BbfBvuhz9tb+jjvbjExvklVq3kW/ZKQ/JsccOrInOWUmFR9DbUvUTqxG0GN9cGVVBN+EdMmvXtc
xXbiJqZqVs5eYeF15+M9cfTq0NLEQot21JgTP7mJmVbj33Y2n9hylOi4uBwzcF1JveHLA5WRVSQC
p5tuZwXsG7iY9/yS2MbhHMXy1ZlOzhap7howzQEUkwVq17SiX9X5mmOTJ3OBV3ySkbIpR/l7ndlP
Kyis16pYGuqtNj4JRlAQntKmVJvVvCKXMwi4ofqjWkv1Zu0s86XqjlUG1fVYFX3VwDPpO1nKzTgm
0ACfelMdMzT0Ry02G3xNjJ1UD2n7rqg5Au3lo47It1qRjPO7Jh0r5df9WRUg2me+RLmATlWbzpIq
bACuVMEUDjw2S2E/W+vxMyJKoqdRPEX+O9KAuWaEnoMKTclMGY6jATMS7nuCleWXshUkXeBcF5np
hUp/ps76VhuZ66z+xBhG+eWkjqcvd1RVUBQ9jEn6l5fpAr2dsOHk+dZQ6cOvwy5UR+UrVkFJ6Uz7
WZPXtBCz1w9mcMA5hiiuWkesG5uMF5myf4vhfvoYK0SERWKt+JgTbIVhaXIhEfhHjO4GjwIFuqhR
HihB75xmqat0iq4iX5CYEr1bpZq3HrZuMLmz5BoFdS5A3SSpOINVLxBJViQ4e0XrOP5O8sIB2RKV
uHjcc16Q0SVTbD2LQTFdwjGtj8r74rZxYD5XKg984kAIQ786HC89dgo2zprvnQDNLWxFXcOsJZV/
FveoxJQRKM7MrhyCd110keQLBy8RJUO5StxnSfC7xVbqn0wgeAmcSRnaM7tjk1+KhBiftraZ8Nwm
3LddDhE6+RzS9AK38BEztYw/KT88eQBpC/9lrwJ7uzVBvqq6aAFLBwonrIBAWNtBnlhZly9cyD4g
3eebeNWrAyHxyODRhi/L40EZJnzl6awrH3NE8kxOULpsM8dZCy5vto3A93tNjdTIlSVLRuzZcRzV
EjGiu70saXjYocKFQq6N0nsfcZWUzUjZYnS0RMgUsbVujEbfBqDe3Jzku6PqAOMuIBVqTFHcADli
ltP16TjjauPtZ0WfvSSq6lydHl6yxmmeKsI1UGFOPLVAOdmhdo2L7B8xsYPRfQCY/boChpSq6jOW
9aBMEJK41TlBCB803l/imhLq2xmaLOrHyms0PrbzUnCWC4cdkeg0x3WBBhshams9PT4TYx0nO/ze
6HiPONeKJVXEZYqDyIfhdzhhsgTlkrpnTVCpPxUetTHm4pOmyaCXvrRZlgMMtWLbvrxWO8m5HsD8
y5VrrEOXRT2447Ph6Ot2FzLAjqxG8kAj/K2+imM6/oLmbHvnsv3nn1ZNoFmlfdb15RsZZqjun8Pv
QAqzugyqPLHAW0EMedNmYXAm+Rp7duuuo02rFF7mIZ3q69f3Vn8TILlUr23Mfro9Eq3QbkhI0Zx/
OyU+TaCXgHsqY/Nv5vr0ZhSFMToGi4hBKMQ2je9rx/EyZwAtwLHVixx0N6a4s6ZnD/+KiXOXUBTt
YM2AMnchL8g6nXmbWwOZ4GKyGZY/AiaRYguZeGq8yLFY0NIbiwvRrMJKpWv95aPnTcQbAWOpEVfy
jNijtZfDyBdqFzKpFhxf+yAWucQIA+cIHiw/Bc3h7zMl36zdLFp1vwdc5Q3zkHtXtm1zniXHVriT
rJhp1pC0u6ahgaSSl1LxnGm2DVeKbULxu1QCYsu01rKHSDGpULKXD/J7a0kduNzwLs6YlQkbyncu
MlGMP9J0HX2SkbFCK5dvO0tplGRcAqAoqlCm0pxqjAvjfxqC4NSnusrKqV5QV+JU8CH7sllOCqub
qq/yE3fH7YMxE7gM57FFGmc5d135PipRGuh2KyTEZrhpxzRdyn++N3bwa+ED3XrAjzvYEIbB+bm8
UEsjdkgZS6f72H8e917n+V9DLsOC2UctPIuSPQIcaGL9uZkYwEg3EDsmintUGe+f5zSBiCCK1SH+
qAgfyOH4GM2otaFYO8zdwAkTmYHIjfMdTTFkXEPYBa+S4kAer6PKrBJWmI8lln8VW405vS5CbMwW
Q/n/DWe1kY1F1GaGam4KTpQkztUoPWqwvoG6ee9JL9XLRpNCdABe11YSn3eQnBMnOhSvJmBU0K4T
iKYJ4kKMlJoho7rH/cBli7OZyhxGf/SMAz5UB/71AQEjiXv2NS5meOk9gztVqipQPP7guVa3AeOp
b7nj4eITdbBJmY4xUg//fZlIHWm82hVCzf95iHNpvUCH0THUuqewK+LTPqbfDTEf2RkArHnimxuZ
pE7MZkROm5BcMfmRO/1o3R2sy3j/1Vdlew0VIhsbJnt8QgbWc5383oKWCdzktdWQ/4ayoe9ce7+g
MZIZzFv+i9AOcCv+GsqLpYy9g6jyBZpSJeZIYKbEOpm7bIi5m6N9f6gu198hgSodFSlGgz2nO2ur
P6Nqe0mDXLJmAGaxjiJ3qbUvzK2cOYkz0KtI1b4cH8Hyz4FqbuvYFZ/la/d1uWhxSjxXgIaOtkXZ
9EpltHWtgP2qHielu3aMEVCMlztsQORzOglyKI4sU0/eyuj14OguKt5DEHD5U+M7uQYAFDo1PbpP
TdWm5ALD8/dd1dHJ4PAU/o2ygPVgqZrllzYfztAx25ZnCHT+nVkEk/DG879lO58PRCPMHoSq5LIz
HW6KKkavEl8ov5coiyazF2BW31iakD0WlaBTkBbqRw4EpimCziZe5qtIhqPNJqR4LoCxWi8fh2E6
1BDlHYZd2O0TT1nvmFosMQb48nyddwSNI3dpLLw2kdHi1oaWTxxdMUjBRCVIGarN8RaFTXtPWLh+
zw6x3eCE8hSJQCdj9rdE+3E6Kw/pPsPPQasYGqGF6F6i2p5Pxe6HD3OJMOS2dS8r3ehTRqcdT+1/
OTKtmnRyks3WURs7GTcZBO6CZZK1ocMMcob213ecPi8XgrdJE2Qzn246rXooh8svTVEu9a5qTt0O
WCJ4KuW7KWa9qCEucoMQEDqQY1l54EbKBxIbImsWEXbryEadMNIkOGFvKtrtgq5LJgEpRGr44U5a
5i7Hil2u2NrysddilaL3oLf6NSu5Z6425bK3dAVK6fssQ/VmFtYo39pkms2sOZGck+SpetRARPBj
gOu7DiTW5731WYlWOc+3vCjgkSFaAbvaCeoSmCTXKzYPPH9yT8aKoDEuAPiUFu2SCvy+nRTmGeR9
gBOcMr075pPLukCOX+QA+wGH39bUZLXIOxzQy5NVf4tz69NFLyDK3PtaaiQ6PC8HvxyNguYmO5qi
t8OIdUyQIwtq0f7+lHs11rE9dUY0IpSF2pNNpDyXlcxNqMgDrICWmRmqHOSeMy1b6WTwEApoOI0r
2+l6aaS+Avr3Jmo7GRcbdEkH1qv8sGsjUIdmnJWCxcRZJ9CpHhmjz95PpW0sKCvRVEWRmBJs/Hij
uKeRZGl4F2VebYRLAJGg5SJPQsGCAoiwr4/q9oeF08MMYNKJQ/hcNpPAD7LMrfTVTwIe03cl1B+C
QzAl3S36qh36VHaFPoab+2BuuvFraUpbq/AiLH0w+21zUluW5gKjZa69HVkqqOoT4W5LggS++UeS
s3x8FN98aPL9aSmHx/QpIL35vJCY2rW2uDsaEedmKzlmxuHTgJcHHs7CYstrH7QAn2gjDbwbCu6t
gk8UdaV3L0FPP2HHNOodBFXYxKKmVVZljIwlp9vO/6dnsKFJYByKiS8/WtBf77E4yUCu2lWtYc3E
qOD+qPuaJdoQiqduG1n3Lm/PRYI7bDBUU6aq8npB2HXsBwYEuQ6HBlRTVsQSoj/F5JHqolz5lfqG
mwi/BH7ZNCap20U+U323OGimLvBERs7EVds4YC0tybQIY3ETjmcq8keIyM+YtsYLPyLv6d7gFLPJ
59zNFWcuSaGWpobnVjfgsM3rBJmj2/EmrKTFD74e0DRHrDzh75bScfFrmwrnZwehRhk8lesUEqYw
GQ05hzP6fZ7pIiTPCKqw0EBP7pIs28fap4O1C8ORwoFndadReHkWv8KKm/Cqa0xVpHM/htLckpQG
p4EoslWD2FqnZF7aprH0koGJasgcawii/j71yulN1JwGIUsZiltDSzxF3ijpqJWiwkQx0nE+h5AV
y88MkJhGsVXCoIyagfIVl3aXZ+R+kL+kpONdzbJENDaDEn9XJsxul6zCKtGeF4Kn5bdE8Cz+Ib9b
+5jrK7GZLdOwvRAGlp60MqsIC3kI+D4uyHYDKUGMEpc/D5G2QB+pVPYO4g1X9sAtdmLdqQVeKihJ
NFwDvWqYaaNdDShgclakmJkqCoQVI0vP/a6/wNkbhc2c9IFwGYkpvOvswM+5ATkBt8V8zLJE5Rpm
dBzbJ4zruNspNbYpUYaHPrnDLLhxxvgTOGRR3M1Eoaa/p5TgVB81Ur2eMydgJ26WL5aAggGiRIHs
Twcn211J4EgLTNRF/sf3KJc76psnNNngBgTrQQxmD9NFJPy+0y90iEtHDHzOvkk8JC94Vx9KG1Qc
rAXEZseMtNW8mkfh+vovCvMxB0Cr9rDTdSYHED9p1c5kUUjTqH6USxuYjxOO0gKAeHfJ5oS09PUt
jf8sGQqM73BZY84OVp8pJ7/VSAhn8XkWhqR+BbEK1qTsuB53LhaHvuntFDvXe+272ewiY0g2geXB
rmIvlcdNLhfmZwjDUQhegf8EE0bUrXPciKHz4Sux1AchH4XZInXPoW2W8mdW2zldPJ42I2D+SUsW
xtD2C5HPSezmji4DFX6yPb630FjF8YLaT8Gc0SuV61UtDQ87I4lbHUCe/LfnCQb1Dzx4lJ+Zbep9
XEwEnEsSAv3HpL9yQgRjG1hnk2zRTs9VMFz4DFr+4Q9a5hMORIXzbM8vfaOlCsqo5A9j8hbpgB+V
GlNsXUJ4iWbaTPrWKt8GrPg51XJ9mOUg2nDrxwAtWQED3vbWU1hgwq8IRSF3GnoRsezD0aYtaROL
m7PfvD4RIHs7njVFsqaktHyK/eC2s9IcwR4BCNy4ZGFgoHsjNIl2+Nrsfz2qZrDN+oz2QTWsVBfJ
KNZixp/ClDGnbmQe7aJ/EIzhks5GEM5HlRirItMvci+3Ft3SB70Tq/fNDD8TofNDhpbi50L99QeS
14atNNubcnUk3hlVwMG09jY6SCfD7OIXUenAO5TAg96sRti+bv+P8TRWc0aB2TVejVqfTlGGllCG
80Ax0Jqm0CLihfi0Knl6Xz/CRZy8UYbmSMTSEBsdyEgen5gZLo+y/uSFYmjq9Me+YtXXhkerd0eW
xR5066cMsXSv6MJPr3phUzGYKC+Ha05JOEs2pVoTnV+m3TrhWa6pOFbf/gX+qCDK89pyC03gTQUo
zaZLCyOF+A/KADMbljSGv4/FsSQ3dBxx4YOyAQA5vXduHYCgg+oUDzeia+Cbcbqfi8Wwxacz9WLG
Eb9I9R+xZ4EYHj+gcxjNOc9SS64W3lWafJ7rvETzg6D0RfAjmrEQMhgZpSVv4MtgwBA5eaXIJkvz
HVEKSrm11XstumvUuybeMlB6sZJDTYcf9oBtObF8gaRsDkOovyh8vBVCY/Q/JyR11KnzlAQFZ9b/
BabZFrbLlsFX2yWKH5Qi8xnGAXByDIav5Kq0/lhiJyL37hRGx9MiDfntkuQJ602cxuBasX1TyhYc
Swe4zJh3Ouv9bd4WPgwaPj48ZQeof8DDeb4kc46TuxTZ7YksAopds+HXJ0teeeuCbYceQNU+4Zk+
N40q6XhTzi3jwYrPgnErTaQZ+BXnCjYuQEMnhCx17d5SSIBY7scYurJfSgrs+etZAlru2et031X2
zpQ0x3NbjYPkxrIKj/VBYOFbx3UhmzUYyUzESJ5lNPFHir6AMy3gt6egsb58o+XlpL/izQrMAvyE
+16rcKuo3YhEAh0uwKmaCQooaVHNWa/ie5HfdrAn5A8FTgfViYM+3FLF+CaKZyF8anL7hamWWc/s
Ca4eF9apPQlHiqcEKHKl0mR6XCLi2f5TF72MJy0gvX8GmzVfDxl625QMdbCJjpd+ZJo3/CU1VnX1
PxgtRta/j6/1e2/b02m+qIv06pJZD6pGpLVZuiTxCD0+ZbnfydrxzskPVbFi2xQ8G773YGSfme5U
UuS4hWMn48MS2co09NiqYnUoJbGBy9k+uo2UuA5gNcS8kHG2ABaeFqQkXic/X03Al1uDnktDlD8H
x1FZhLBkywrwxi1J83wiCfzkWDiOB4DmcbgGosEUmcJWQh5qapkrcvP12lkCV9iS+4YBuCzgZ7uv
awHuLDhN8ydXZVkvIVgl0B3Y3KyjFmgXJBgzv6xDuZ8OBZt6lG5s2j/exf8PdbBUXgHA2t/3MPgz
wLzQsPVygTLPnbDgAkpU+KNTz5+WMH2v8uetgLcBgjETaoOEBzrRnnmOePwE4BIVVB5Z68en21dj
hqCXnSCbyFgDvvlBPdUdZIH8g7Ike1m8ZoXbFlVjFpgjtXw6JHaOv0hBzLmAL2Q3JrTun2/WAbcp
kyrC9gE0tVSL1cZslM6sSTbfSb4Q4pxM/dSeUK4f/fIoH4xo6mWcJtlpq8IItw0mYS6VAFxOFWgr
0BfRrN3har3tKwPjGhd3Lvv/tFBsphbkybdluZizHjGbhsQP0kZNsbEetTnQSnqprcsMVcLZOt98
5isf07d41e+dPCa7fjjevQhc+A+54B/HfBldVc6MDb6Ce9nV+FJj/Yv6yLkDvdxWwqkX0tH4nVHD
/dWjGkuxIPqH4SA2Q7n5+mC+VME/aIjk6k+IntoZulwvSiCBzF5dYhIdFHUiGCvjM0+Ln+Uk5Thx
jygoYFkaVkDJEVidXamkh2Jq1yqXklEkYoqJ57QscWq+eP728KbHA0ZUL3HvdPAVB64nZsdprnaS
333vj5mM5r34AGnOIDCCGosiPIzlC5wAe7wpPn/ony3fFeOSF7JmiOrCQRHwh4hoJHkqsxqzxgit
QAnWFtjYI/zLQbssvkmxgbuvxgOs0MiRHDw2TnBCAIHyy6SmmWNkkrCk+Oyd5xqkJ898d9n45RL8
WkFgw+CGvoeE8Jl12noqITsWFYtPK1nECu1/xsauaiMSwzijdvBGvcz9aBHlYYY/TbaoQoK4cj82
D4/iSi4zRJypAat4uC3U/ZYe+BylPyeW366K1NkAgNaoNrP0koD2FTBROmREhi883j2muR+BaxOf
BTkapKXi9mMlFMX2OiKhgkbnI2rR/4625MsUKMQX1igm4jS+XJsIptJxvzn/FjtIrBovn0Q1K3Be
GpF1MvSOhBhVVMT5AFP7FqsH9HunEpT6KEdSfLuK1OJIq9d8jrNZuvaluqJJ2MBkajjOYdSxZQsk
n4k78hXYAWlIZkp9/pONo1j111dddLZ2ZScHSM235iIic3CtWLIYOwh/JG2rQQTzzD1AGDTpaPl2
pbuRGBwiw3wm78+rTwUxW5Mt+ircM70BYLg6uuO8I/wpxGME1r/OyJHARFRLJBfHgfsU0SxBzfHr
x7Eej9sqG9Mfs0H34DN1fXTkpTatptA5gcPTs5KIH+TDFnakbm17mkwKeI/rHUM77DV0o4jwgfab
6XtJOYMlah0vDeZlJwiyBm5g/VnKO6x8ZDXyFIhuivOgJkbn3VZMyOHcx3ZSEZLLlftXeYiXCYg/
FWDL3YL7iVvrDVkF3SN7hVu1tarJikKZWRDgbIm6THaXd+ZP00BirhVR0f6LWsM1sXFXg4X+9giD
uXESL3V2+BqSd4kEevOnRUuEESH5PwVeGUvKsXke/DFPuTRY6mrXqg7QjGWZ1OCXh4efKEiJke8Z
3VPNJvztXn0yoQv9blfYaEGHtHkr0Kx6KKkWf01rGwj3qzRKWgfPKQoQ1Uk0UAh8zXFKGmL2ZX5T
q7A1CtrKL2yTFaZNGKHL6IAGCzBqolkHp3gehzMStmm2TEE/f2sYP8MOmadfIR5wUWkM7G9FFQ3L
qBfshi9xhuhR1DTyRWODlpZmDnQgP+l6SehfatmtZdU1wfsc8MmmgAFq4JlQqN4hIJOt8J1HZBCn
+4m2Y5CloW7X5yjYJyuyGhws7RUAsq3GbCILX8OV6cGi+Q+zKtKoZIADEL1r2f69pgZfN4U6twI6
J0bfFgswDkQvjPouPDfDYDWZXUwalHTQOkVM1jt0+LgUj3aTF05V0arIynYqC25u8qhmpy0n80Rq
e7zcG9eQWPZGHqL8JJGporUfKU8rf/kIbL/zmSCeiQjIGci2BPrzTap5P9vnGdd7VhBJ0ICg6tKv
VlJboMQERFPXVF3Enl5fDe7zyZSuRSvAFJe19enQFu6BicBIR0vd7hiHscys/e2VBIwIfEm0NnIv
wQIywDym/SpqFt0LpETygbnJCFhhOoePpp0KYHujozX0Ku2c1f77UZd9DHuKKRu0M7doHs3mjkCV
rg3aPKuV/1U4EQJfpjOrie3hctoJdZ4XlVzA53f0LI7NvDwEOUqw03/GgSr2QadMyV+kUg7aGN2E
4bFU0D9C0TTCw80R/FziX1LcoqjsMeJQf0AL7aRwGEGln1geEZgsjgU9djHoKHIUDFW2UR3tH9po
emCkHqbaWMERl7/b6+E2RPXbDNq+x0CDphNXbsg+IgJLSjK8148gUO8Z6jHJ9Da0JEMwGDuEMK4T
m7htpmcBeXYR6dWva1q+rgt/r3EafHcDQQVoVVcyk9Zw/5D7fHzpyMOwqJFekWEw/UoVz+91VIoC
cU8CHvNya0NtTfmPYeiU6Vb5ugHLc9eGufhCp+yk+9uwCOedV7XHfXN1oA8Bv1l3aUPqeHIH3DTX
ZPc5XWvs1j3B28rtUKJiTgCdXdEjj18D9CtZatFjbCpSLwiQNZ7UfdhOj1kFY5HDWe8rz6wXgmzu
fGooezMA/J6GTLLgo1FSilnR1xFgt0TY5K4hNU3RE8s9KIRoSPpM99FjgLvogVhMfAeeYYEnKiJX
XkA++EZ5Buiw4Y4H2gqjIWf2Af5m/z20G2S25J+yiTDYWLFMOHrYeGsZ8HOBxmyKIQykcNeYAgKj
TjPkiYGikL/P4W5MQlOwjKvihXexqmB6HcCNgoqRUvMKYd5E4A1q5qFPz0LKswh+LbHSlqPd1OFk
OIXaejZfAMbyskMQNQclzBg105OmYGuIQgM5FKRJOTPRmctBSmPkWC/TL9zc8m8dwB4MiZLtenfS
Og8dMDVZj4PJ/OwFG8FL2fG3WfpLjnqfWJJisEOJgyY8telYV6UX+cwt0UIPpHFKjwkKukPHquwy
1X/T1beV+tmU6LtYVsESk8R92O8kOoqnkiOg+p3H4pOPOJDNNZyjUpwOb9mEFTENKOWlbtIME2AH
Y0/rxZDW0zlxNu6q7rLSixOigMmsaVXYpYmXb5iEokQghYJ4p9/28QBMd4QOV1+94otn/mEvzr89
HWwyygSz4Ve+V71AeN8wE4fb7wOC4rid5SIR0SVilTkCVmE85BismkJVZ5vfMYs5FfhCehpinFll
N625XQraqLsZBdUfsoahTEA+F9XBA7D8sE+daRnMwaPZyoWQxhtro/eVcIJT0NuGMOiQbnquJaMH
AwDGfApUDp19EcFpDzLSCvqaXdC2T0dty5OYb97ZrLB4BXRBD8WPJ2shWsym+3oHU2xMSsZ28gtD
mDRApsM9ytFKjeJimzU0UvmC8cqA+nnzHjzfdI3LJQo4AfvGEd1QIMZ9j5sBix+TAGgah8aRzbiB
+b4x6zTq6dRBQ2p5UaYpTZSBxwoJrVuM278JRCHtaFUpipY888JqOKkCzRIT82B5cBvDWqiiRdV1
CJlzd0dFeoGAbdi+FadSUOAo0eLqw9VI/z7NZDZEIw6UyvRG2YJL/iwiprpN079ZzoDsE2Yh7gsc
qt+gkDnvW7h77y4wMcnPxFIScRA19sk4wQWhrNTN/AruG5rrHrvnVJtWHiN4aTHkD7VILDuXjKCm
1ApIvGoluboKkcJmzkUV1TCEBl3n0nhuD3zd5Ft1kx5O0ijMS2nHGcz8r2AJk/eNN7N/7dbtT1Kv
a9S3PLMphrk080wPljFgiYtpzH1ZtIj1jkNAUv4IQ/nwsscGL6vKJ3p9AJ4phPSfZnGBW6X9GFo7
NEEwVLNppxPJvU1/3phr7v+C7aaO5wZWM7+Lk+tFdFFycSIaWlTT5mgHyPxR9R6rnj6816b+eQG2
/krAQ03OyZH7yyeWvKCNcnutLeKgylwXt6KOEF9JO41/hBvwSsnuWc+kZI21uLLfsdv23dj6iH0q
d72QVDn297jJ9Z9FpxCx/wFG0vR5UKvI+w9d3CM3gvadSVnwwNv1Ff2QLiAztPUsCo1vOEazusLI
W3ykWMz0L4QmGMGd/oqrbM02JOaqP+EZeIDwPBc5BUUr9gk8O1LATKSAzAZVK1/lAnzCsH7MeVgu
InfbK+a0FIiAIicIKmritt3AAX6yMp67BMMWmCP+UjukFm7cfFYfKpV6yNjdJzi1zhyMQtbmuQTm
TTGfcp8vf+EI53BCtTUBmWSwgrNavG3IcuMYA803JYyogb8IXtrxDbZR9E9LBdWzTHhtrYpGO+gW
g01oJWkHgZIT40E0cv5VuGWrIc0pc0SrB5M6ZoRsn1RmDvw2jeuXAirXH0eCB8rTGRli5xrAS5Bu
NmAvXDoxZvcMG8uRe0Ya8a+kv6a5j71wNAOsQXVN/EE5UyJyvYpuPgqEha/l4c61zSYB2zgJFn1X
XzpWmJjkedsFVJG+JkjWwYZeUleIgWTO0AHkNerPSri/ZqETDqD26CMnld3XRuHPoPRdoBDtYbeX
MB+gYVWUfYlqeDh5mPKfjhDUmr3NVO+0lpZcXej0dIrTGU2pNCKPrkEo85ge2aemSkH0fwHDf6pk
o+ShWxPi1YC6E015ZH1soUHeJbIdxHSr6IjBx5NCVsZVVG8tRVeD1UfhyxLBzU2wTyrMzwdx4y5U
c8jpDseX/4pEjv30XfdrErWaxJwq9r0Q5mcmb31CppZejX3m89uZUU/lQPVXX7qn2NcVlERIXp96
vvvSEXzj8uLkMc3Doyo15lTlVC6JlfeQSJp5cbCasZezcl61fdgKTze7DBC0HeZ6GT2HD5xw7snc
p6Ds9paOFsjKRQi2OdV9LLZzLBZ1h6zrmb+EJzRu734SzgeOiNmRaqKyWUNndfAxfZ42BXlegzyY
KzK5f/96LGwVhoqlPowbw3X8fm4DFsAaYcTiNMTKBujc3GgUFOnyzSI4CRVmlLxMgC/1VQpioV60
k1qtVUe05fgYVddQI0kvjrfoU+PeI5tStksF2C4FlsGArkN8S4QQZfxIXGlt3n8yWHU1bSXXku5V
9LFNKJwaqns1OzA4ZgiBqBGwVmU/EOye+KEhp/RyQEMDhptcpgExkZgy4A0e1tKf1L31Y9tukkr5
GJlIsX76qTetkcVWCSry3fzco3/r/1OmpfqeKe/2Lmwk4CiiJbEYrMpNs4rrNPFVO1ADI0FKPXyN
AHXSjKrybG5EedXO2H9edIrhOn7bk4urkGnXcZdjvzdwC7q1cG3pd6RIjpeEk4WSXywGR72VYu+3
r2g0K/kwd+OIeLtljLiTI/wZDUz1TyT8KbFGcEgXsnUhnRH+UWwtOWZJe0RgHwv5i0j3m/cWRK9K
CnkoDOfb1yIYfqx5gyCPX1Ic1NQ6EPgvlSaaeI4ennsyrPDVGmplIV0OPUgYmhmAwLi4r/8+TmI2
MJMKDlNvLuMY7zd9iFg+UtF+7dTRcn//x3MNGFHrFdAPokNsJn5c4bPhxU3+buWHITkSXUbxc96H
5y1YN7bbvTH4GseFd7dXyMDmfsKKXHsp9LpUloV5ZOJY8Ae/DmWpygKqIub0ujDSJWyfLSAjBthC
NyxjcwcVT1bvlZ/yDmx8Zv4M1jpaWh/kuw+iP2KpOi84W0D+yF5KwU4w35QIvEMGHFAUFAFqjiNW
yOKXvMlK4jviG3yBumF7E6EBFSAJ3Bbppf7gNi8L6/Inp8B0d6u9lrdKbKThRwdfSenkbKy5Slt7
VPZ6Xqtds4boV5IpVXwnbtNndvGhQLgeX3+7960ECQg4safy32qT2bSK2enDjNK04qCQYdOeKboW
+rHlSIoQkdm+tF2IQAQHhXNA+RspiCwLzVcXwb64jwcjHDcljuXCLCPP/FzDU714NctbhS97dd/X
YdlWgL0tuHsXGeY2tuaMgCIIwcry56t8g9gooYfkvD0L22Z8QVQcrRJvSqIZ2AJqtiYz8PrijiHu
etX5mKRVk6Mbfn5g7W2MwePeL7ZV5R4TMYvpGK2N4D2E9z0yRB+HS4a7k9ShmtvSRn+68J1YGgBB
bdiKo8vDn7LmQaqNOUMCmfQ+sRBSXhCvPwBR566n46+krE74V7rmW2AmCWcj4ovZxDc8sIda0Rj5
6N07j8/ekhPCopAPZ6zcGBZ21AxK6jdlsVctPIXFzh5CDsl8z59hwJ1QSvfr43CWMFkmf7cTIHVp
eI4afmHszv/cMhv45+KMrO+ACRAorns19w1St9UX5KibOKdyMCc/auP/sqW5AMow4J58i8UbVkVb
32R+BXwAs5EthJS4G9Yu9rrs7m3ZpsDkt4z/5rMJ7yJeU9dFpGeSNVG3t+Lw6pnJBVavRqtZidYc
2L8DehFSvr+vmTpGoeVIMD1YSI+M2CDltASSq1ipM3+AP++9w4OH6XXnmUTKxqSDKQN1KXVD8hlG
ke14mlxUg++/evVLk37kbV4V2D2P36Z/rxfh0NsaEWsI+7Y8CyegbymxoMIafF3DsPoFss9+g2xy
HfDCBJ052LyuERWLndvVmGkitXkIcZHOzxGMpyz6blf5mrQK2K/bCwH0wvbiqCzMcidnDKNiISEP
fhi3lXLiJQ7o7rJbD68gYGnCoQGD0ZzAAO4+mrZkU/wZTvp5wA+5GKeNuQQtmJ4GY+RyaYkaPiEA
t7yNaf0XA2r0s117jT6CZDaG42IOhuTS74v/DEWEdLsemFMw/qUjVSgTnRoLoRN7PjfdIxpKpEXk
XVpDNzarId/szYuVhOtCoj1FUwlil+RFB3aIpamIia3stWkeALVNv2IQmPZXPEmnLZLtJEI0SY3B
tY0usT/tOBQSvXork/PVrF+JXcHDXfDjsjDnrBbt+J5vnyDiTR3AY6y6gpCJopf6NA8vKsea5ki3
3dze9ozev3rZcd5kVE4yQ3xctXuNm7aF1U7WrUrAXhy1/oV5vtIilK7VoOyTomAvi7o55JEpwOnb
NEQm2yoQDdwsvj//voes9wpEbxeNi5KCfZ7NU+luZphj5A3oc7N3Eg8+KvUvzUGx21OmlGY5CP0i
/XhEkJNy8m031ZSbNhxEZLf+ZQRAPvzSQCI0AzN6QwbshTG1+SJJ7BLlebBvM/4J3OyYds4iUFVs
fXlgJG5/8svgRz7zg8WIiNSydWNQFM2VysvsKQn28KYGs+chOq6iAQQGkg8g5mySpp81GqWaIR8W
Vvj7DjdPATpEnYJLbWSDv4ZpHQatrkUbXU6DSSxqJTtpuSwU5jxRCUVNL2IuFOTLwlKsqBKuMDHh
3Au/Slj9qTn+s8iB9LckGh22MTAKrA9jXSRd6zg3nWr22ZkYQ6SJCWm+txHOKL9tSY4WMAoD6T2p
sSONVcnY53qe5BI320wbk0sHnYAqLSa82XJ++Ac/oHVkKB/AcK6FCy2rGOajCGPTiT73nfyhxrGO
+aEZ8TrfWrNjxg1q+5qzcgbT3vDqk+OCKsfZiegSXtf8wY55dAgRue0tDg0lbZ4HvDnulov+LevA
Gon4xPYGIMoflEQR9FUa2FTy8p30RsNMEXcV/AHvO0UntwfAvePYB9qdmbkp895SIN0lNlXMndJ/
bdZJSmaYcN5NID/sHebwc/vO4Za8TJwv3TxK2i0q09tLYSqSX6tLAHcso3AW4e/N+H/u6Ewhg5c8
3y1WmHjmdxSNpBqkEotWTVRsAg95OrCpeFX5agD7j81b/jxMJHlD4ma4Z6kvVZBbPJr+b07lASTP
ru0nuGU0PsCOKWV6iKj1jZpUaHG5/d48obTn5LGI1XbSJrwtaoaEnjoou8L3abP4GKCrw7uD1eiX
FUXGHuj2WP6J7jKzT43udmfiSEA/l4L1sE/ReZ0eMyKryqBRXb4UMlUWtoNqQbzbdgeqNwrasOSO
pFgD9qIjndE87B/+KO8LjVKfs4gjLhXqf6TF3t2gOQ+M3lXn7gc8gHwWnUnQmuUSc+WGJXkwEehQ
MZALEjtnAIfuKkcSVQ312XIwXOl2Wj9/GMidfuGpLVfQJ2k1y3V26b+CmdZqA3+Z/793jl+xfCts
GkPMzOmPIW+9qnLJdCdxUE9BMWgEwQSwbYJxECjAi2naLgb4YRfg6xWSIitB4jLH6bn/6W4T7scO
JlgV7q5gyctQdxIto+v3X14Iq+CQDweZqTQr7HaHVbqVQKKWk8lsF6u9itAgjWhozrVUUYZ6IoLB
edchQ6I6yswcfqAr59S47vnBjDM47OK8+FowBR/8A+JvPrSB39BuvmBDqD3BcLSUtnWUZ6Am4stj
s4+sSB6UJ42mY42BXjO+QbOu6Co4VCzLlwcHiHwIBnvwf765d1fEVOcw6i0EHL1dy6R1RV/jXMwG
p8hULYX9MOV53nLp27RQzJCkD3Djxcvv5kt2/3kfDy1EvMyA9voRcnqkyMDaitRy9M6OrZx0ZTOh
f8WfnXjQnrVdNgeLY+QQMSJKTkxBr6NQCPZsjwMrf9LnlWkcM2WGOqbbiXGoCHC2mLaGR+NJ5Rj8
hIm85ZdVe5Oxce8SqtqD9wqaJONbzwhVmWNuDtS9Jl41vE5JKgt48WW0Pj/XoVuZqopduqM/k/lI
I5c2vO2V3HqWLbxl0fOjVz4xW16zhnRU2Qd+9p+sqR1VgveP02a0s3fMt3+tIR9jPDfFS9sAAVlK
Kn0Hde/M0B5KIX6F/SrDzpj6OxSPZX9Af3U2fQRizCaucD1NNpad1Fr//gh4JdGN2KvAquVcNwir
FjATYIEC25zh6VbYgYaSgxi/F1Ul/HWxquW9ppyZ5CWcaS5AuOGQhZ4eoyxgmUzfWIFndd9WW74J
cCy5xRC0GHIvVDHX/hrnWWCfO2K5BRvYCQItFKhQgmb7Yi1/AS1WSRL/0c3ru0hlJdwccJYJ1ZQi
u6dZQi1Hd/0zHEVI5/iSf+wg7lw2/h5WILDTxYUw20eFu9UyrbB6nsqaI4NHzHU5IZOGNKP1z9ym
surb/TYBKpJBh0qjKXd1OdDCbfCfsLdMgt/XSZC+HkddnqkinzhtrTe7saONrR5fS79zsZAa0QlZ
SSeaXohriKpZevkMPaXxB9UGm4q7XhmiI7OnWPYR/q2o2GBbxb+Gt2c8oM4SyINTOTqVHmsTTzaK
v9h8o06HK8eOKfJ/8wBwWUV8L2Lq+Q0v4BPxeNlWolz1Ib3/1ykB4Xn0OM1CS9QieoxzA3XK+hRL
eqR9ej4K7E1PKW4is5+Ffj0tynTaZDCs6h+isLb1oisrnzR/CsFfTzqgcqpPi2K+0O+PrrgDg/yb
JD5xvLaaYrINt6xCJL//00PW2/ek6A398CIBqflXal4z+I8kXMd6tfrsCeBgW4UIo4qkxXy4X4ix
Vm6s6XZdb+zojIj8wiL4mo8FPRfoewiyWpDX4/NDlg2n79s5YbWqu7j0oa2qMWFMtWPFUYo0OKlI
fYurZ096QQn/3IjTWmks2UukqaQYCFiZ/wWg3yU2gCaKsoe1w+we9Kb2lNigSGmrWf8lfb4kQV/8
SHxt1zNeWDguwc1QzAYXHO2TBQBmF7xyDjv+1egP0ZnicsBvgQ5D3NxLaceDPlN1zqxs+3zyggKM
mB6zkHfU7x0oEagpoKu0DR8X5UL1FC1OMlKO3fliTMwIY1ETRTtKkNN9MuqOYpE2GdUKBww4mKB1
MNSIJHlTPzJfQ0VInnoB5ROsm7zLozBQf8NPuty0EOHeN04/EVruTiLb9Fow1yw8rtHv9P5AuPje
btpWGpjC/LoScavkyEOYfanbB/2l1bR1h0eg0O/twAwFxEWOBFgPdQwxO1mjs9Gdm5tXug0bnTLs
rYHGe5bFVGfX6o3RsDvmLpStgbWP0qmCgT6/boFXW7wjid1444L5bV1HMN/uACVvo8wjjByYDbFq
J5mZvbooTiEmPfWKarauUC8zVeha4UDfei3hklB7KQOIRrW2DjCbNkPeTzGQ1YqPRS3jXLE9WHVR
eOyelvP7tWdxNInHOpFeVbbfxqvLDAFc7r0oksRzffSA0c1ne9pKEDkNIbs1JTId8lEtYdBx3o8e
X/51SVnrsAs5GprHcy1uOEl3oQDuh9k2qNBh/saAdD+C5M/ZqQTpBQX4x3idHGG+1ZANEJNMgCvh
ra2RxnxSI9gkKPQ9SlZH+qIv4d1jT7jsPi0i9LR0/EQVimEBu0UE37IKlThyGWL/i2nt88mQH8nx
DvkgqavGV8WedVs7eBBr8zSN23e//5aafVx42l6sZ+NfM29WiIVTlkroZJZ3SGkUmOate2SvvfMP
STj+mkvbSGhLhGKq3x0gxrvqGIyOIencc2sI9xQJjsReE3/Qndp0HfIqpvAbdSCRtJuHMeH1KTYS
t1UmR+1nXsUPDnP2YFcX920ZR68hTQoWDLN8qxw4xwM3fuxn8LQUxlLLF6jYSxlXGvHkfIudyTI9
LfLhYUeHVprhu/JV/m5IVMXrEFZ+0oKDhXgBuqKirARgfzy+Rdmu4BnKz423GrlA7MObi/Pf8QmV
3s+gT4gaCOaK+ZZm4VWhJlbu9f4CQKd6Hf2leN3AFByobxtvwbuOXRCT7gLikF8357DqxGSATZZQ
7eYZFCdbPjCdE9SlG07m5f8ktg8+2G6yhRNftVS+AFq0vkxLRlgtOHjhz6vTPeGar7AR4NoKMUx2
AOVmxFKZdjMaTGBzJVNe4wdaImzGHWK/k9gb1qiLMeUMW+TFRFW1j2A+XyQ9buBKHnYnZHthX9oJ
Jm29NdKMRN+24C0d5Adr/T+Lx33U62cbSTOS/yFclTHzU2+aNg97IfRmJ1ty05Q+ge8YggYnwELA
yommI1RHewp5vCky+MLwGrrqeAMMzr/6+SdEFtxEG16q37Wkyr4J23sDmz1U+Alzl4yAvOD5NqSz
6ZJUGihbGT71MrRS2/Wb+3MMe8q2A21EdBmsGMsnjhKRlgDNSr3efOXXAdJL7kEKPu0u9bOD8res
BTcjNNeSOTMPI7B3Kl9oR+rSnlG89gXwb1DszspBV9IJArqJEcJhYruUiotkJX7XjTExZ/iN7SOR
uoqDG5e56xuofr8K60xjx4gO4bAneuNAEvcw4ochw8vywddPSdBTL9nEEsFWo6JUO/U8LeytRF2t
78pIc08dtVopDYtPXeWk3cNCjcTh8u92YadduRI1XFw7E/dN0jZCU090AZHrIcSY6UJiY/Qu85ck
tMPWE8chHVcMmaCuYxwXdTr0Qy66d42f16+gKoLViepxoyX8wiVVcUqTXV+dgBS08h5Gv8Q9/KOc
YDJzSA9oyNvMl2hBWGqyYA4ZfgJwXmat/hJ5DwjgHGKZTJKQbn8bcMOIWH+mqKEhkYTSfTzOymY0
XJMrOak2Mo2Fm+rqxwsqc+LfikCv8CyP7l0WgpJo0QSy/HFkfqqXPoFo25RAqytMnYFdYLAYxDA0
8hCJHtOFj3gD0KxVXwnbPMKyt2BAnM2uMjs8mUm5yRqTKeUEjBdFmThiLBGJP0NBW2Zjtk5qXk89
Mo89SJbo6Grl5IhMur6S1JJIGCdT4KPAKsesZcAdEGC9HtiMhUr0AQnS6O5mN3xgQqaK/ntb59OI
buPUo3LJI0NBjQH4LBp07EjqmhYgnjIHuLcXgod+FhRZcfA9PaRuKVkbx2l4nshQqgYovEddiBgK
YyuHhXjnDXunrROky7f5eWy49RJnjcsm+lI3Ji8V61LWzQxzh2wsjzh67pmh1Ry3cZSvAK4RZp8B
6CKipfkDluL8GOa3PPT/qsxxPM2ShcvZJh+AaRX67PfME2RRGufq38nEXBbyg2YV8cht7aGsNPQb
TuVV2AshdB/UgR8S4loduWgAfJY1AisUPeO89hqcH3/Nwe+o8mGjUmNGQ3wXSLsP6XzrEautOd3E
+l1+UXQovmxiK5DfnPFdfERNZyT+djWwFwv9SayEz9q5xPYj625TzXsxyQD+jeecWcSuQ+voZNcH
951kdvxWEUkBRGRXo5pj/lwME1lPDgwfUaYSu44AhU8eyEXEKNnGC8U6GNUR1IVR9rZ5uN67MxQ3
U16tP1NsNEPDYZhpnwPdkhvENQKwQ/t1rDEOrdkZwmXPLcIkX0sYz7pF0Ph/7Xc6py81WF7Bt13L
itiYAdX6U/QS8YIsX1Tl8eKUE98ystbt2GBSX69iaSNuIAuwQw9uAP/tXBwiijFJLQwIWg98Zs11
/f5/181h0SjUfJNRjkY4wLad20QtyY5mj5+j8OPIiFD1J+aWOkyJH1nKjhcOI6aV4p7kr3Eax1KZ
LNy0LWeGVSEGHyDzLimk+EiMN5a+ODJRciEQLTxlQCLRopQ5I6hD15A/ifObLhZswTnVbg0jamGi
BzQlWuD2lCdS4u4qj4p8ctQ2X5yOQ/zCMH3vXJuq50rzHNPoRraV4/xb6umJPzcuJoDyGnwepG3y
HqtL263HmLvSV3RMmndDIHDGCXCJEUqnP2H8SziwCnzSvaB7hVqlNV9ZuTCmL3hLSo384QxdFiFW
Cw7BUgArdumBNgZqEqrDYWT0x8rrlLeFe6FHbgwGKVrgy5bhnBUVqTuAJ1Qlf4hO3illk+LwTtSc
W/JbvwyxKqsQkjHt6a9+mdwE5OTaP9+A7GYyn8JvITIP8mFgx9GyZBBJuxbXda4QkxfrNwRBKyYk
/a4a9SCQXU+7zTd3PRnsw7lZo8ipFroo3vEzV2EJUZoUfjY9q6iwdesA6i0j5i5hHoiVJv2/d+F3
HdQgP+hAR7UFq2S6DG76RCgZ1q3R9IKf/JSuHCmfjN0HicZf9ydBFjzQESk4UDt1weaM4lJHu2iY
TDygR/u0hJJhqvymwNis6lVGCzxKCproZCnqV4k6qtGV/dAYpfTTMIIFlCb7AbaaWak/3yiOJ0ln
pMjBlXo5Rc3v7wrbHZ73zhMOMeL97mBBve8y4OdIWn+jK1M9u2yi8zTpOQImMrjAd0a0CYEc6Bis
mN8kRRQrSYgmvp+/WNVxokYjNyGH/+fWZCgX3IOlnNxxvrxOQhTEW0R8ULLX+PnAGEkF73fswtIp
4uoO2+2+v2mbLw8ZV0dwrcpkL8jmhKsvnFPXWvjJc5ppq7Fxkv1r9t3oIa3PG8sl/L44qw3+5/Ns
UZ/UtZmOQgxiDoozGEMiLsFEGDYNyevX6X7uaCb+ES7zeC3UXITTIQB4HUPhUa8kIdPNQoErkgkU
MLN1Awj1M7jGnF+rwJomLlcY9RJczQMWkF3TNGGx2zqGqOfOd0hdjBrLyiD85pkYSd6JZMJujJkB
PWiuRwK2QZJBiI4SSYdQFCVqqQP1fqoQ/sTl+9/o0oaNGBbfQlRosq6ADrMHkSpufm0E+7UNEggm
oVZsLg5yJsJ2EBwkJG3bytCTVHJjqC6r2/sigi6IVyR/qi/Xxl85iZI0Aa9oLkFY/l/nkSbOYkvm
IT+6YjhIAjWFshLMEEfjwEPDjZ++CZeiU65JoWLrFMAwby4IFFRbr3LnPsbE3UXF8cgUP8Zl37Wd
htQCZcd/uvOHCQ1rgQlvSyMH0bDiyeNZYCqQvcRW4U4B/lrIeu3J1q9AAi5KBBLCgsCB/p2JuFXs
aNow9EQ4BkFhRGh1ilwSO6hvjfz4L4PBY+n/XcFOLI729bDBNAztq6C3KcqFVJFnOoKnJX3P09q0
N0X6ejPgzetKfzfqB5gXLi9LlivkII8L4AGSZzR6KncUUVZXs3yS1KFYDXGrYSq+KXpALAXd97BE
OxpjcqW2ITtNGx9iyYYjQFTsAZqFKu6dIauBTJHWkAFw1V0PfbRHulvhl71qn9AdGRrxW7ufIlfN
JXC/gh7IyXuJ0ErHObhww/Fs+Zhd6ubqSNRGeC63+LJ9Fq72ITafB0xwfN19qyuLuBM78bGk9AaL
fQvEac5nQH3z50ymy1+HxbxXG6TtdbvBHduFqX7ubkrP7iVIClfA/ExMnAfFJhfLtCoEVqa/FThG
wicBIsq4kLgIFSvy6wGaKLs0fdtZlkP7gnyikUoQymMGNa+mx7EiUeV+O036DmXzgXLBI76ntAkE
lGIwHu0xPmfl24b2gG3AI0KeY0eifrWA7rDAmMrdtF6ca6ATP3dV+M4rWeQQkYpemvHXh7dsauS+
VqGvq30ekcxCv8ppcF0GmXm7CJJBquulhZcv5Tu4iNU95mobqomldMMBXCMYlKLyc3VZyWSH0BQY
Npdnlo9t/ouyMa6wKxX6A6UHeFitWIOhhr8CgXrm5PRZtFIhWzBL1G0pPLNhqHcOvqQ6g2jfTyfP
RaOPgqByGvaxHQDIoCGAqU4ecbiWW2jWcPidab/4gVyLvSXuePte138ZIFjtwUQyp3Y5Shze0iZk
s88d5hbx7iGZA+rf6gRRMPCqwRJxYG/314lPvsTcUnfaaDM26zK4C9Qk2JYh7KMBNWoYFWVGejYL
6NGwdZn5I5fAcVIpNeRfYPVL1Kh24zkUqvswB0Ucv0She+nfGZmqELu4MNPtgJrdon+UuilyuVhr
VWegXyRyWy2WkbLhj4ufyZixTWPciKCuLaX3CGeV+mIAwqs/4uu5/qJJ86klb6PCjtjJ5URbY7zm
gGgASOutnosFVdxoRIBaww5TeSErK7HxXnsTWUY4bQZLkChdO9lc2Nqws+tr/uSShbSxalAFumhU
ea/HfWVt2RwoKB983fGhGhGQchrQAXzml8XygeI+/CrdhazWSqB6WcBIY8KltXP1/v2xzY4oBL9i
ybcF4/jpRx71bcYqx5QPBBk6FhUOqQbLIvet38WLr/HQTQRWgbASuP9ki2tRMjr7ppw1K3cynzub
yv1cfiUuBLaHYOMUxVqBtZ0qF0WAzV6Ri9VeIC82YBVbknyq1IYXMQI/ifGV5OIZOPFmG51sP+jQ
cZFgBcAnaHWqqlky06qAX7JgNZfZ40+z+xP4XfKgFZBJ1eRUnSbT5bgQErk4kdt//dSkSvoHZag/
4biTuL6WJ8IZ+TrCbr4HOkryLDooOITOd1AFXMdoP6gkz9etPzV+OvLniodrV8kEqY3s7I8HQfUc
ikSfxOL3qHa8dm3mqGHGDU05XBhF+dy3NWmCAoHTqKGbXvlRXGVu5AVTIJDV+SboAP5XIXXcJirz
w5b/8sGvWUmnNX8kJeFQz2fqyMLoHqxoluSnZa59kB0j96SIbGPupRvReQGQZHfvOlCRnK6lVBVZ
MKrpcdYgRYgAKXgggG7NQYJvRwXzqehY/jKBgHCFvLX50hvTjgBg5HavhelVOCzbi2zIf7QYYscb
Mb7GECC9r9xwNdqLImcEVJOxbCAnu3+wqgBAYokYYOqOKXttDWyJLYfrS70tj58Utq4IggQfjMu4
ZAdO0p4ny7nOTr10gccJ7r9GDFOjhbO/tEBvB3Ja8pvGk7+tEA4WRWYldJO2C9YxKgysQtdS3cW4
/YGWvrsOqYtoBI/fBCaVnCx+b2FNxJM/M1vkKwY0o0n4Okb7EPLv32cj8zQvpzVsgAMxiYO1Xany
SBID8L7oTK4lqwj6luTbbcwieLDvdPoGbb+NemOULb2UIiAFwZjuh5FPt7TGF8jxsL0ZMaPk0BQD
RPBgHfl2oyTUm6f+mRUfxnhUWapLWeocXPetV4p4CVFPHXgnxQxXHdAG3HO4J7VcAGPoR9k+j2H8
FgYC6k+YJHFWJVGH2mrnk4iQ4q9L3IoPjL5J1pZojiXfy0j3tD0dh1akh0AbOsF+/1FqBbCM5X0W
kT/tyzMg8RzVFS4FdRkNHPi5lOF2mgACAkDEDgZe9xZXG3uouuqClyxV4HZn7qN0LIym7L5Tv0Yr
IzGoKfk57p6mxhzMCXrhjqSmpoIaGScc+ON6D8fW2vD4ibf3fCO17ZvFIL/U5HRHJp6VM0gxxOxV
d9UAY6gUKk8L9cJ7E2d1XPs1izlbPD7YftmB7tSuja/4YynsY30rLQ/zQeDHo+QUcMJoo/WoPSuC
ExqwEWZkD/s0krDiinMkBKWPWM0xpmvWpbosC2yiad7Y1p4WGGsZork4klAHlKgaMDTgKfTuFPt/
Ol7RO77ZQYr04FJ1zcfHYGTP1FAC+u+gN6TdVQPhj/k3envFhtbAgdhm/H/shCbjptBwy0UV4lig
J9Uonk0hiFHqCK02NWYaCKa1s0/RYmoq6C9XblrhI0TAOFsRtj1bXUhX9lKtiTPLws8TtOJNmhCa
eI+FRvKoOfhyaLEuM1VIaK1XLcBBF2iTR51P/xxaTugmFtM9yYGYChchrWaTO4JfUoddzXwIwIME
P7KtdLkGaKqufzH2dHSUfewLohPCC/gsM04F/IK6V5sg44FQ1Kec0BvA7wYi255m1Vm/L/y85iWe
7y5J7SYFjbWWiUgec62JGEXZmw2MD4Qwc++S+wvnjTliTPWG99KruO3/T72JJJ4u+ZYShUXuy5v3
vR0sxmazrAFD65Vy5R13t+ouo3+wNyEwI87w2S0DDTRfBj8Kue7tH/J1jX9/hquZ+FpFeTU/Wwzw
y6YtoWKtNQKfgHBhc8zwkgFQiJu2dP3yb84nh79oUpiQSn2nt0uCfO6voB3tQ2Yhs2ZN+OpGiPuK
j3jNK9QE9+sqNAL7JKJZg5XUka6kLJ+XmLpvNDXJ8YAAFPb83Y02GILsrVqSZXWnm9UjgKerWqfu
t4RBaUeq9x1bqKJ2uf+j3vlrtZD763K/Sg6dRMg3xCdIEN227iHh/A8RzXC3+RM4gb8a5Qt1OaWf
hcDIoO4cjpfGrhfsECJwlbNav3EgjLlWuY92w1dU64gcv29HBXKq8bYL1BvFPmqpju1RYbr0A0t3
N0B1Hj1wSIQ4/4EUf/VkNemz8mjq/At0qk8otqva0Quhfgcw4HgSyf8/NR9zzGFVvpBQ2bXXSYkN
dJ6fJq5xmPwznQ90yuwm8+nAFJAZeua+0kgPHm8j5xH5GBC+5otXIHEz8RsXtrwh5zm2KZXqgbS3
vjj1pSbq2vkTh9v9EzpzGVBWX/QmdrWicnZP1hwmLz2R2baBvP66jmIfI0uqvEbpkcLDOL+3kVsZ
A4sJnPhToB1AalD/JZdfxV5/8UMsMPE52mKfZEL6iRB0ISaCFUSKeGGx0voB8sOn2PRfGQwCEjAY
BDUUx8BbdmuaWnhTj3icK76PPGnokQHG2gZLkyjxrU19Pr070GpPEXQ9nwE0y0WPNtyrCRfx2vc4
4tAA+vo+vdZ3h3gyUMLpqhAfsP7aO4xWxEnZ/TM3wRQO3pomIFjB/0CmmcDZLxA9xxc8brMMjOeK
AhrEvnU1Tab/yqpTH5h5+Tbk3Jdv3A6jT6s+l/UG/QDgnN4/Uh9utSx6uOuD2r3yVq1ThGOAgt1Y
f9WQDIcc/M3gK8iMmJsC7dU/uTBN2qZEV3Glya89uV484ztgeBPZbmn/d0qFByApsydtNFN7k2ij
cGMaN9QzKpTDDg4ZVE4yHPcrsmgedUwCekHwaOUrPRh7pfiZPrkV5hKBzg5udq2vUlTv+QApXNbe
82nBnNDniEW60w7n57hPGRBpDHcjHAl5my7iH6DooJCGZwsFGREIwHKC7bkqlxFmnXpLLinm+X6L
7vFQbMvjfUl8hKzI3cZNcyjvxvwbLx3iDvvED1fqWIshpYOceVHmWpkYu3152W2ROw6QriNBaiTR
oddaWw5YTGSVqfukBnJ420nwWUwnomuSWP10b/DxhUxeGQIWIHZDSH5vueIiZUZzldU4p8/GOPrq
u8VzzYqABJHcNp4YSVstpv3X7EgxTYeZleymSvjx8Hn2bmPPgQdinSEucphLdO1oTmFVtR2pr1hP
0rQ3z1uESZ4PRIJKnBFpOywzAVzOwKFR3aL0dtRNUYaZ/T0B4zronp40EBz94h7FOcfMl1nI98pv
LoQddfYYOwy5PgWo/VXLMH4ODf/5/9BY2KYScbDiQzySCrtSrs0C9NBSg/QDyTAPVySWJiUmNQzX
ffD0oFdZYO++WDlNQZx1P+QMjcrYAS3MnYBxeWI6xlw9IEeO9X2vyOzj9c9vtG0+Nto+oK1emCZ6
nVNSRpCPNCrsfD/UiqGdLEOyvZ5NIEwGo9zbbVKMIBRnBgIh+Md2hoDUMqfAwB7hY14ILYHFesas
ntfixk+TNR7xrWR/ak50r3mYxF2M5uLPfxhj17EQOkd4NPNdGojgEZ/WVeW0oM96VnKyWj0JGbCH
8nq/O5rxMFW56zJ8ECoWvG+CjKFVNdsL9oVTo1/imyyCjXuNhCDJmKxubpfw8FfVsQJheGyyiGAc
YzI8vTcIV9WbTF4P413DHpLjdEhhDaQKTnKSD9pvj/BY4/j9M1kj/yRuiXpVe6BWVAA7Z7uiMdRL
vNSemzotgRaGG8W7b4yi8yFEwh03UjBYbCJP7rBhKDA7WQLy8M+/RJR3E1JtBLZi6UZnXPUeu1Ef
1BsuyeCHtV1iLFowgO7Sb1Nhn3kEVVDQ0Y/H3fPgawlFfycsbIk8IVc8ecXmSNh+LKkHRum7kpdM
2I6E7M1Cdz8NFhgT7bwqczcuWx2D1oz3B6exO4M+nC63fatHBeXCXuB/rYzdNSHIzBlj/VT9+08C
Qi9+GwjlvZ2aA0d/St51PsbQFMK5ofAQwRvClbPOQmfC2YMK/+A7bVu3tuIL8fH3/L5OY35ZClUv
LKlm9m4USo7gQNvzFmC7d7UqSHpPfADUK0uCxKO45E7FsshvBrVxly7eEl3ZG89wbHhCzi/mLMtg
edoJ/aTwC/FnjqMzviBVRNG1D+Hp+UliaMgnXUOtrNhwJ+NcvZp/fSlwUFVL0u1vcggj+ivqAuq1
fpPRGVwJ4bKm9uSO3QYsSsD+7jAOQ10TdIo1brc4POFAqftppDPgfEeQdacWe8YCS7roMbiv8mgn
S93pxwEhEw28en5e0HNGmLEWDDtoYgee3RJJlr614yZRQ7BBlbO9vlZ9BwlQfWgrcLIoC/oKN74V
nQMAT79wl8FQx2u6PgOOOw6q48eKY6YCJEzWOutTTWY2vVmGwV1yeSAkoB4nr5IkKmUlrqZ5OGaC
bpQdV3p2THYA1dcf/rYwaJp6iWgnur9sgYejs3Ktbu7QoM6MzmZASdvyAAo4zitMv7zWu91JIn28
ZGtcCS5B3SoGVHPbpHUEku0zmUXJaJYsTN80m9DmwGR+ggwXkYmC/e5VpTXzqP/9T+NbU7gQlPFV
nwGiOYkd7s/dO8Tl3bNU0hIr+cScHC9Hrlc+i2/YXXBL7NmYOQ08Xcf9296T8J6aMvT6/P+TEYXU
fKv92mEbh56sadZP79gjPtBQMUGBdpt5sPZxLlyV7h+3eMO08+Ws+Wb8O5w1gYEK6d0EYToIbQ10
0uPWzi4RRXusW89hyddZuwDuwCDU0vAWgB7oU4MUImIzdxF+fg7RbJ/sGctIXHloFj5VxAfpggNE
r7opRjGnUbNxZXV5HytyFKfyVa2UbGJ8AWynx6TdauJAHvliovDQacdQk+oEifF2zqtXofRKhn3E
NOGPhSXXZm9i34/5lx8p0i8l+7DQRU8kntjDyB2YTS4hK/N7kuxZYHYPEoRiJz+VZV3aUFU47qnQ
hBriLcAAWGoc0wGNWH2wFdj4dYkrDWOry7DmV9EulAFYI5xGJBdivT3xi/2weic5fDaco6VAn2zF
m4O5j5Y0kt9xrCv6uAcKkuCc94wduUe5zFACSgVqWHdCZ/iyNi69LGmaaeKK2/9IEtjII+hybjI8
6R6pBu3+oaJWRylN9tseex3IuTNIvgBxTpPVjrQdPTxitlyizpRVd+PLl1CJQ1ZH0TamUT0o+bAN
Vcyo57ChRvKXmxWggsGyEqA+539H/icEmIzwHY+Dk2fsVLpDdZqZTGhCEXg2Rhp0QnvxiNXD5y6R
tVxKtjDxsbBWof/Z0bKByFEq5qq8jDfMjVLgUEI0TEf8tKzWBz4Rq2LICUFZKQiBuvI/TSP3Zc+W
oCwnQpyYCBjipvl5XXuhY961Tlx87958ynwWCBnJkdwbDkDxGuMFjLaBGkn8vgVuUZstsB/yg/ko
vgxeePfih2gwXfIGodb11mPwIQQt/gqbk6aq8MnKlAOTeEsZ6S/Kj3OcboVcJm1muSsVOifMuTa2
6VgPexcPuq22JbkCd+fqV4SIuiSEHr2uCrWzdYaav4nQTHXaJeIfsuVUo9TUnqJtkrblG6b/iE48
nMl4Hr1IUuXH3F7skePdS67TBb9jDsk0rR82ZR8Xu4+i0J+hyCzNr2tFsrda5SfZhJEpbNDyiVZR
JBMgOvo5kucNpIF+azWqIJK/f+D5K0yG5Gtpw+MfOcjc7Yz2mlL9Kk9hLqzCHNke3ICf1p/RfwDD
ki3lSzhCC4pjs7gSJ0OtsVwxMYdM73yuQyuIXAEfhiTZNRmrr3OJQmajUJ518PkiwPzTtLRuyMwi
LttsCRRijm5giIPSZmVLJEG15txy5AdT9VE53WUt0zBLh9Nxo804v3+hRj5Ls41UtzndNSw+K7O1
wpd02jruUdOTizUkZyxGZdTuCMPzu9R0Q65dPXmC7v2wdGQ3EPJjcgFnf5lDU/F3/qVbIN4nOyI8
Hzw77hC4cC7e7hBHTaVe5jAQawJsHftwkcz3T8rfDPfsmt3g2nwpJY/+FZZr3XjT7yZg//xf6VDd
oF0WXxb8osELzbI3fDMNbu9wZSb2N3IlN1HFsQqIzDib2UyjozYt8sPqSm6ZXMHqG5KrQ60U4AmB
i312mueSaH3rt3ygSzMHRyS1E5VAl/vO0W6kLWC0pLtQmd2quZbxmKuGM9cn3j+EMpgeHWRLBp4h
D4x8jdHn/AUSXV5CLLH3Fq3Lg9rdIN4k3Yn+4iOUwZuOxGUoUq9Phede+/kTbrEv+f52TNIuadsw
uDs9/lQBJCJBsolX10z4PyF4gm2SxW/kzuLel2NYTw3wYH6Ie8Poz677VHDulZjlO6Ex9pS5W+Mq
lwbhTC2DQgo6foX0FvSsaRjFY9sh116EqhIPM5PHhn0DqEudYwv0xz2Uvzhb1Xt5PS7PmSr2JhRG
LqslFf3FPiCMZxfuViK5jgok+8LTvCzApnCXie1z1oVahNUmfxXeNSByzMlP0qI0Or7V/9vtvS6S
slVfPiRS+dKkWIF9oy0DIvjLZecAfYhbC9zA3RTZZ8/SJGNZuAIi1XuhXLfims5Y6bn//6wx7hES
yygNtmid526GeXmexISm3AtMHIlPlDjXdjZHkxmB/uHEyEmRVGv2neygB2CLe5P4AXTJLD2SD4eI
plZV1zb8javD/INqYd3vd9kzEuttHlYoIhn5oyLxKlFqJUXFjNKiX5J1x6deeagZc6uONJhfSLbx
G4PH+RHiLIWNhEevD9Q9o18RuZmfDa2Xh7eaCmOO6wZcF77IjokAgHuWNh2MFEmJtbvx51MUUlFK
d2d6QJf5RQRrgVW+DxYJ4ppPndhwj2W0dp9FtbLPSD2HWUAnwGUny7mwSwjP2MCZsxTQqu+aYWVx
TlxXavah3j4TMhMVt7ZwhxGjpB7i+QEzynya33U7Al+XuikfOy1OWTGgiMZCz4qjuMwSDsRrqZ6b
M4LKYpBZLGFMoCE1aL9APdYrX/R9wpUxtxOAX2hQchwZeAfvrZ6EUiMdEyYOhRe6qfrFT20pzcFU
A+cCtWaThGmzSLq+scsv7YE4HTsXxX/FaLI6F4n+hoIvgcr44EW5pKGDrsctrWdix/9K0NqoZkjM
niDOuQ0J0TjIz3mG5X22G5ruoCpu3miR+1IF/+IpVDaFzTHYSE7z2oMAceMbwdksnvdb8wn8uI1n
gr9uBH/WXj+XKdsCPgkx10Q7WDY03v7WOh7I8iYbqWFSiLg5/FLgl+KeVljgnDp7g2LtcTkTF0f5
L+ZjDSQSiWeEiyxtJxr50pBWvEpWKfN8dGHmdm/AZn4a9XDjnz6CLgeuKXdf99ZqBV2QuYkuJQf+
/rnN4Pzn7gSDHxP9oTtHDidDaQcpCVZIEyUM4+T7oKEGTZJLQQRoRy6Swtj1uJnlZYcmBDOGWM5g
E8T8xIma47EBEUeBkG/2g0MhHb76KausSRMwqZnUff8t5kigq/MZrxV03uc62gl+MqVunrkk1EAx
d63NDscYxMZ176ETlC9e6Hyxz1GGzZKHg61uNr7qoQJ1J4o7xQ1QZNMQaoezZk9cx8P3H8+xiFcn
H5hV3xBN9kVlffBVAYKecB1ZNVW1CVyAgAt+SSr8N8Bge9pGKjlzBfQ9AsqD3FZF2qVNtelfBcIX
tCJF/29Dy/tCKyfQNr+Gh7Qwlp7pL4RJG6E/q9Eai7NloTfB2i+nSAQ1jIwVjsLwz3NbpkGXcvKf
P+REpALE7aOJcXU57jGe8oWfdFt03UC9RYZEYQPNMQAFto70ELGSJjQ74xw8mpqN6CiP8Ek0d3b7
NrQTkshFCH2NWiEW4EVOkVbT3XgaYGtzsmggaZKY58pJJPnpY/JpLHX/l7b7IwM2pji/D0BY7RD4
Y1Ne/oQzL40FGvfY24vSMjIjvnoDABAkISZGNppI15zsJoMLrKPoLA+z5OHgYS+RPRbI4wyh4gEA
O5tyH9vCyxB4hQZetTByFgdTLR+UU5HwUw1MMKQMkfGV7uTTkx9wq6RwWkXKxoDmmWMp80oP6yDS
jjNJ5QEyeBW7+L06c78+DBDe6opMGpZz5N/WMg8UPKvXotE5AM4y7VDW2JtZFw4xlhARy3Urg1GA
BrHkSc/4dSownfIMBAHlEoi7OqZI86g2+YbROaG07pbg+g/Zs/rAbEz/1A1qdpZOxTzVyLCVAQsQ
Ld1vtaXk1RyLNvQqrMfaXaacC6ZzdK3H30g0fd+F/dmk/viBNVI+Jc4VY7Ft5NVhr3Fyp9OIo3nA
Ijjq27MXjwDroKs/XZZ+Fg17NWL4AoBgO8u0NPi0ETR1aQNA8uVqCCkZpIkuxlzq2g8hpwB8QRGH
F165B3tAnEd3Jr4LmYrhD+vSodt3NDYwoN70it9p3Ifav6oNcwGliZCJ8K3ukUShin8IgjawfDVj
f8Nhf9yvrk6FgMQGH3VUlqKjM2UTSssXLmm6k2ztSy+W0fibmwq80WZghOSzXMt9x6QhR+JzZuYy
n4FUFLvIkRXfS3u1Skl/XVTBiZJ63YW+S7gpwD4nP7xs8vHA4+qwpz6k9JrMyl6IKQGhpv9zLZiG
bd283YOmQc2qguVPZyBUjcbnvba3wpmVNQIFlRxiqPuCYO/+vvPtDFwoZdVTQqIzTgwLsh/2F692
pvnbH15QtEV0ZXrZxt6ESt+/DglTWrNQ45kIphDA2sk8LX2SpXRmuDP0f4qqDgaXgQkudBM14QjF
5s+LRub/7VjI4nrrGTbiSDzpXOPJEs0+gR91WGoxtuYcaMXYyEv90dg9AdjxzqxSuHAz5P8Y09q7
fs8KJyqrfi0X33mlLoi/FZrW2KoPL6HqWE5Qa+iwQ+Yk/mXD7ViTmdtGr6OnAsFxVspDnUEMekUu
UfWO3LrjQ2f36A5ahSjfEI8ep4YKHr4HmaBUzfyDsnPnbbPyLJzsqlWTH/xslwzEMVQslAUxcNz9
3CD3XdVFdnNHl5MBclh4qlUHEUomS0k2+0i+OcAkjsr28r9G2z4+xsdYGhQnjJTt7FLp5zzOMEIP
W0eJ6/PnJIWd1Yn4HQNfFKVL+nLz0FTwhilXqtsfQ5N1TOMElXcBEu60Su1Id6Z1zXHnLo0pT5v4
V7Cg6NF4BH0+DAe40AGsz99T6VzRb5pw3Nmcx+iSfw7VlZT8rfmVvgbGmrUEQZ+WlPoVssw/bNRe
Pchy6oC+sk6dW1KGOoV+E87WtnF/31bvuhy/0z/kLhqz1T/7FJoHzYO3lqdOem8DVY1E9tpY4KaS
Lcox1OF74ouFUutqW8AvwVifyi98DAaiaxhl4FKcJsflfkvvFv2pcB0uqeLac3ZaRLwQ48BKO/KV
f0VMGgqIth8loG7tRk+W3lGv5ruYeeJ8L9xxql5u93iTBhNMpIVut0jP8nF4ouGfibbu5cOZwKEU
H1UHQiP2ygb2yk0YUjUfR5u2XQN93dQnMqx+Qz7riIafkzhvE5xPQXX+TnVyr1O1Eg/6kJaQRcwt
PQd8QyQDNo8U+Vzd2WN6a5tfRnFEpzHERJ7QHw4B4qQpw6J5AAZQhCemu4reACOiceJCSSaNcqaX
8BT+5u52lAhE9WgvVUtcbHR3SeiON+R3Hir9CNBV7W1chnOWYbgz20tXRrWLOTdWqYX+vmM0Zj/G
0d2nvi13Qp23XMadheNJl7YN6Wk3N3x6cfkCVppEGznE6JG24TZoNUw2chXImEWeKOAtw8G4N/sI
cVozEsdhnASqWT4NpuuMP7BnD5oSAjkEsVci40S2I7rgagKn6R77i0qIvVcftaPXosoWZ+2STrJE
swT5/h9kK6dPnKOnomHOF4g3g/A7ov1fJ3n4ngSX6LtDgF3c5LHZ6Fn4+6Ga5V7dR3rD4EeLhVUT
XE194nw56oqrytGK8GD4N/oY0/f34DXcjVIo0bhSF1EE/kjZ7qT3Km0Eo+8jw1v2TyHzOGUdmqa7
EAvdlw2tHCQNUY8KJX96L8PKSQgEPPE0CmuqGKiICtxdSti7zyaJnv3t97PI2RIyd1CQjINiJ0m7
NHbmy7JKQQHRweUT78jvUl0EsnQ0+Slu0FmEmoIf6rupnK5YlkBYWGTSwJLHyyT0p8IuWOtJxepW
0+jpskFutI6CpvKzi7RjfIsZlJ6zK7NDc4dJnz1CJj05jsa5xwad9a4jR+uVk3BeMBH3cxKAEFmq
fa07yC+culf9ng89PlEusmC5P80z5HdBHAm63zmYkMY1R/VTidfqmPUHtO6zn1U678SPj+ff1Bgt
c4GZpnilOD8Cf681rqG4UdBYWpCC2rzQBGrQmsvjqRnZrrBCi+bUBdN5lPV6WbUGZpLg7KXCn9Vj
jS8DMfL9XrxI7MFcfao0KT5TXGw5Ncfb352grrV/e2mEvWdOEFFFMSAhGl+r1Pe7zSz+phPyrXeX
niui6nOVhmRSMaj6gzJatWuV5AI9x4sdhaCk6JQc8r21BtXw/UrRE2OuUVqjZB+Pr8fbpSGi8dd1
1Kc6lzfw7V9DrKScXF8+QSaZ5NTBg5jW1rT244kZ9hRxvMWSBngbIB0YEv0P6lFfDeJHbLf6pBCw
olXH3/SiUxgKVXj14bx+HtOjxDqJbud7Q+ITz2ckLMz4kSi1gZto9z/0s8FVmgrYkcgIcNJNTLD8
ahxptUNpBfeNHrFP7xSUsIuTyhS19dTNbzEdjC+p5RDIOKpsOL5eJLq1JqRop2Aw4NhVS+drqQ7l
nkN1rDTyol3LCZPxWCzYEplTnhFOjxC8kels6NHCrneQWAZ5su95GBjOfJFqntgno5PhiBlkSkmt
wba/e+HENz7zxo599+/EQfqBfJC7BUDNE5lnXrbRNLKHCObkZaVim6Nvs4+WFbGrE+Cams4byDBe
o3N1+ZdgfKzxOkExtP1roCdmjOSzvykcY6VSQOrb1b4aBSo28jcWvHw7Q7SJzTtCY4B/TKFI5y8v
4WJ6azWLU/3AC45v3VmYb8810lSunLIUMW8ZEZiCC6AoOxxberI7ljNU6cg+lvZRYz0FVlRbAz5o
ZNePSDU7DwY8vu7k6QRv5antJf2Mzu3TsmElO5OL24IsdeCqoRS+rCsaomGCFNdKH4kXOvaaBzQj
rzTgyJTfs0WNezH9mif1N85qXf2IyHgGgsSu9QYoRc3+XCKbVuMdHFfV8isyR3KvmiwqR1OBnCZn
ZGOTkLfsom7rAif9XBrkM266l3Ytt5cuKJdZnqja2BW/WnWdSda1BwGS96SlNLX3JGIv+PRX4omZ
j8p9vrB9/kVTCEBfDWOniz8ryMMb7B8mHJ4ShANyufdR00pgGFwCmYbQYXe9hH2eugRuyYxWcPii
dkb0a1TQJ/bA5iyS5ctnSyc1YhI0OFnv2xF5NqjXBQAJbIovx+oAVgPcpnibEQPhDQ3Z41BOX7hK
4FpgdlWm1zA/9v2NVYeHOEDfQYe7OJ9g57G4dsSjg1WhM6I7cNrjLPizaiMqiODUcDVXE2CXootn
naLQARE7jfF7LHXK8u3Qqcqd1XzMmuCqjSCda99MKBYxJwKvaMyMoZs5KCI/rNkK3WHLxoYgqldy
6vsd87h6uGwUffS+EbzdB3hhnTbVLx3tFq6rpvszK8auWJQ7XGm0RE+t/idoTy3rLcublxSt9WCd
MmQca4bm/huQM3WcMQz7dyUcBG1ceeZraa5psJqJVEf4NNZ5avEoLRVQYQISWNgGXdu+mRYiKyeX
gcZOoB2gYXH8wkrqzctcz3VDBEG95XLFcPdxolt7rQS8ZpOc8Egw6FJ91KIFuS7dA1z01WQzHDSw
Wo/pkEwBnupiXz8D/ywAr4S5XlOetmxUcZtC5xC0Fu618exZHphlXnjBDDLQGBgcN8C8oLLNVWrh
wqi20e8Aw4KURo5MAbb0iaKfMi9KVqm4LoPoLjr/E1z6MfrvdMjZbDWRq+eqegsnJyBMH/j0Ocpv
hnPNQVXj+MG6oULmwxwqNaK6F8ORPTHm7D0AfO4s2NPRpjlVEMXJr8tLrO3E4PV5F43S35WhhqgL
qQd/S1SXKdidhIFTORZNFMPk+0WVHlyVQXGZ1dMZyXzhaYEi7rqZ/VuH1svwBrvkWPh+QUy6EBYr
z9PoOwtuRCurimJmSGAjSTmMfJr8VYqOdH6fAn1/N1/3tmx2KsMx47OF4iEYb/ToAPftSaK5eXsr
Z7RPiXJSDBLrwS4zmcTxIs6IsdTcSCcCllg3k/5F2p9WlHC2voL0N7307NosLJHmSs3fS5vIrnyA
Hrgc8qNkjWu3rqD3H4GAbut3SVb0Xh9eZM9t4lQn5/2al9P2+k+ccINl00JBMzjMtQ3Lb1Yi3eSa
1DHx+pR7uK6zAhcOf0h2xvkXLYPQQhwy0Yhvr7pf43YyEvKZ0Jsf4hSIUimnifbLgdvcRzPE/nwH
2GXXUr82ETFt5DXYVjfzrn9TDvqNK30cALg1pERqF/08acB+krUjbuvcBGiqZ3Tp2/eAC6TdbpkZ
HF1WTRPPwhOtoYn+hJyjK8EXCeXvM5PzPDL505UXjnFisjM273oHzHGQvC42wKCWmMP+PE0ac1fM
LcRr7f+gxbDz82HreXusVo7wW4ac/SpyyrTqG+RhLx+lFmV/IWNHRgbogQBvux68PY3sm7yUo7Dm
ljPuIDqHbVzUwgfsMFTX+3KVqHUWyfTE5AlDJ15/ZjUai2sDnM1lRT58AVqwVAiaKQzPBFarlbc3
1lo7xr/Wac0sImy8oFtVqoLlGUtv+dglOGvsKr24cGK5aYUGPcatkjHV5/Px3UjoL7YQq2R3VnyV
7xfpam/y7+3BjTGOSZK9ftrH361KQ+bnjDlhrpguMAkSnvRGY1n5StE+ekOL1RSmhWikveUQqTYV
kKC/swKCQaY8ewkHHCOy9D7/t8lSAZjZotTXXZjBtkDyStUS54hieO8dEP2BGXwaYbbsb8tYmpHB
Oq/yH+G6rSS0AXUBQ160rnnSFAKV5F1+BEY6wQtvu0r7cwuRnySMiCAQtZYwPhjh5JO7HpZgWF19
TJCvmPQgrxaCcjiFdMszeBrJsT+xb2Egs/I3kqzCtxuWm18j+P0FxAm2MAyQtizMylMBX+vKuZIt
zgTi2U997RIKBi/BC2PggyTAcD/oR03W5S1EfomueaBoQ15cOJ0/fUokmy5OjUwm0VdkSOOt46dP
o9hY5dcObsH+4Wc37eWLoMehKTgwUaXeSsIKRURTmGP7At9z/QSqtPw4odYAqNo8bg26ZaN6dqtb
4ip2ENhg+jG75gdkIDW/rb1uzpJKeCNX2MyA7+gh9FbZzRKKu6aHCB4YsGPCPRsrAfCelUjQPCfJ
k46j8veHMV4Xa9DnkRBGiNJZc1dnXjKLDZaffNwTpNBz8mq4AR97fEv3+ejOd2s3/ZM/ZiFLTJLf
MyXQAF/TnILtdgEcoF+1K+eH18ANYY4Hnxv3q4TJkjcwwFUU6XzVa0VeXDmpCwsbP1nBdnVRlfE4
WErzXbrDzfjeo4jTQ7XynDOFBnNxv6yTKNaaRzJOCb7LXvx1OUzCMHJ22XyZ30ExGVzyk4QbNhbj
yGRUtwbVis7lKhq9VLD2idDno5PiUpamkvwXxrh+Gd+RI8/eEl9rPI22ytJ7hkWjKfulgjbSqQri
/pquid6hdOynDp6wq7n8un81tttMxDAo/P9KiyYn//D8Uu5nWPDcx8G+wZRf1okkLdFTrMa75Mm2
otauQcu1wb9GkyFStk+X73CHQdtz0BNzmYFMbt2hhLCkABVx1Joou71pT1OCjrogc39OfJW0CUY6
MNboFUNztplRWe3aiVTx2fNfz8dlpd5niDWRp1DDCg/RhxsmvEzx+9K0e7SXnJByzOZ0kCk3/9s7
YHFNrDsk1fmmeFhFKMR/QQzc2i9DhClr6PAz85Bf7sul1ORyzlrC/5qU6gTWIAOWkmO1yoYPH4fV
QS41mvorY6trdpvHTSArg6W08JaRBimms3G8OHa/DJs1JhknVdT0/YFwP0uJpF/LwYllGFLpyB2O
0ob1/JFhHfwJkbvvqzkefdICgUZXYF6uvEL1RgsBh6X8or7XOAjmj63U7atVgjf3jnXZZWLsSmSe
eolorf9iqJIsYeLWiop1WxDmWkDTmTI1VuZ6L0IzBNeBRxJZpsz80CPQDY4PX1XP0Zl+u8tqU/Xk
vZ13AeyO9/s4ErNyZWvbmf0cSYfcuK/3UKQ1ukz7++MrQjgJtXJLV5Dnu1vx1SPXnVl1sFg4sAzN
8rT5cKyXFK3jIDYbAjwsRQegXSTpY6tEq6FUP7d3B1QlR9/RNZyr+ysuwdb6+24eZObMgP9BiTYy
v8kSwj37O9QzKutsvAjcIavq4MpgVCGVI3yV/r4YZhX5vz9/UYd2Bh7ZhXN/tJBKJjW/R1yb+qY8
19Xan73VvsdHS7P2A+bcVJkayxF/cdypfDaqfPDyTC3rlfu0Q1NwUgsFZsXb1sm/XUR2aRUwuTAV
eZRBxB7NQj2MI8c1aShDk4V3A4Hm9CQfqHdjJT5sF4TjJQfqvTlLBUptNllWBjEp1DvRlqWjt6WD
+wfXteqhGWgF/Yg2QWekX7ICNYCTmEWZ8CyHZSBfMNyU9dFwvHtBqnp8RUqdHcK6dWB12ghkf6Ww
zUYe/jz4dltPJKoJd42zPhOvgsBPl9LWR2trPNq6APNkYCVQb55aCvpZkgOdBGqIdoepv5ZLTrUC
xfl2LZS38EQH3zNT2HTomOnkbCOfO7WSWbogNXnFsfnavv2knlK+6A98iqTE1SAIOrh6YnDlAtw3
9+l8RpfhV5jjKydkQKYgJL4YOUFaY0t0EVE9RtoygzSOZo7bVGgW36HW2WarWUKLOlnCBdG/uwjH
VIgMeqz8V1BjmYFqcQygjXmFaRZCA1vwIFGhN7B5FldC+qvxQg12sFDyKuJMOMn5054S9R6fvru4
v5ZlvvdrbOh1XRexBcORpYcBmrqr8HFhwntbJOidyuGuIGFcj8ulIOle4sXO8Ycelx7TJy2Wi0Dr
8w9KByyC03NIn/VMCFAElLD3CsXAvGnnKsbdrT8y6Z2ZuYzFaB/xi4AQjF+bndvo11fyHAQrGBo9
QgTvkSvsI9CGKyXSydJLJADJPKaV6hutqlHxZ5BsKfcnOLnAf7ahOISlS5ptYKCuhvfNIPvpYput
tVlnKFlTG6xRBnVQDcZ3/QhRxzp1UcNrAYE6ymSfP9VNnx7hvBkhUhtmVIt2hfY/zlZexUA0DjK9
ncXDwS3DA7EhyRFl3TZ83aEcngLrCi8o4LGrnw+1bNACXplaUWLmHsMhfIQGCK8p97Do+aBRKQ0q
XQcdyj8ibB3XRRPyeLIG8ibp2eeEBJFfk/XzZBuYI7hPUCoREw6lYcB/PfzJ2xcMHNqdr87FnJpH
5s8DhmAuKwAzZynEoQAB9+8QrSsUmakmuxrafOQoD1Nu+ski1SuqHA748oS1y9RbVDp3T+zardEc
tIp/NoTyS9QX1RdsZZydmZy/zhE1E2ujpfVpkcxO8IO4blwOjzbZMjEkGl+VbR6WAaxC4TYth6Vt
nEqel2votLwIdNKZGlsvZxvD4sZQxbe+Moo/o6St8tT3peEsUPDqzwcWp6j3vxbyqwfdGhEResL3
j74p07BcY2JWUlQmkppJK/AMtBOIbiFPNwoIkZK3TujxXpji5bJrKMzuWljqpQKXfPI0OHlQy7M5
+Jn4imeYOFu0p8YLxXYCh+8TtcPfcGDZocMlHWixrWfv78LsEiHJdfdCl3YQtQ3uebuKjALWyiIs
dbJvMLdA3YS8r90qkE6nVwTJ+PCqRVw4MV5OsIMOk00HqhZhyPXdvoIaofgmqIKnhcfdyKuxVXux
fqq9qVxME1F0rrZj3EDXmiYM7kuc+A8M3QpTB2KICMiBcqIAVDYTP+538Pmej0i91OTxPC8ktxMa
+r9F4iDTXXSc9kVTHGGVEDdwRfaEWysdhjw0HaLvKVFlzA7tx6UktShbbTamZim7C66CrbSU7mT/
mvM7T1ZOaeBLwa5TcmNORSGjAW6jQS6PT76Ya7FvcLzmMVaL5BF78RgMpZucVbTFL9XSmLGMEkPl
xloU0jo0WJjD9U6J4aQ9BmgLZs/oM90oHKgeEYCYmbn5RgxfXa1ZziyQMDlTLCoSlhhxwRkwDgGh
8Wsuc3aeTNRi96kOOdK6RuNCTJguxvWQTiLHrhtYM3vUat+b4jd2wDvvexhVSx6ubPhn5PpPU/2u
WR7GsXo7GD9JWAxGWPPmE7Vfzk4AwuoKZ+aXRmkZulg5J2cxWaCM5rZrQV/zAloCn4zvEmuGgtzz
za77PY7wzlxIFTJ0NVayuGw/Y264OXMdXVcifUmnwQKrgkvHf1UaHDSZo63Txrto//o9KAY+73lW
uYrbUKrAJeSMyNeQJ4WtbBSxkoJKhIKkCVJ2I4/zwNdgQn7ekGUZzhjoh9HNqKh4pICOP5EBXDUB
wvahGpJ9eHAoIfvRHne2NIov8JCVDS0mwXNHBEeID7t2HgBoglhTPGmwLI61mYmDsO9Y6IeOqAFg
SJcO6D6I/y7LEHa4bx6Z+SVPnB5Gyzapwu3tMB6JHq6ogbf1PmL/mE6RzGXJPN1J33+RChQLq3gQ
hyx8/wGlz8Usj6kSVDZHTICPqIqKKG3ZeXF3lJtM9gzVnklNFboTImriCXJmA2vq9Dhoy/lUgArP
Sq2S5xY7GFzIE1n9sbrYw2/w7ZbXzSr6KLlUZZFzA5dAHTT1sYAYw8jkY5BhRA8ascu0nOCh+Xc5
rG0EEGRMOLasfsHzUtPlVF1+LzPGdA8vNGtiz4ZcguV41FD9GSmDlJPaT5H/K3jzYQM0eBo3hMol
TqVYReJ/QFKrFXS3Ve17Sqw51pKiNqct17z3Z0lcKh+roViDzoXG/eVAgFMR6ABW8qI2eI2HrJYF
tevG67j/DxXjAa+AMrC/rPFwrK0cqAuwyclDqRr5DF8xGuBzht2tvE+BTqPlYqIF+gMNwAkfgd1h
1xQPYjE+oHSMeD0Dj8bABFlqpWJGKnb9/dvskEp/9TyrR2pWUnltikXED/QpJDTeyoPW+aFWbXmq
0ZLneBB496FwBRKTZIOP6JxSLbnn4BCD4AFI02ZyHFpRqOswjcJ2Uf5EyEf5gon1KZqRahepMGD7
DiXpqFg7/2rcBGN804V4MJdEYwe5IjrCWR8ngPu9DYQvvHgJVI0FNPBDtk2f9YZ2AJXrWxAho2wj
HP3SK024aJNZaIhIDQe7hDsUYHoZMXqO3L2h4Otja3IZP8tWwnEYvtjvQWcS44H4oRnGianxm/zj
gwmuu9vBkeuBIPdboY1Ni73o/Dq8jrOUuLPaljXoKwhJ77ESTNvTSLOfNRNwRghWbh3hdOP3b6ut
qz2mIaJvPMTS4pwlHjFdMiDUF6umgYwTrsN7s/nZ3E/Iobvg1k208VTTCCNjrcyvHvSyA1oYw+Dy
uJuLfUEhH0H8HUyzDEhcBrssddq4ugu3QCkzdXom9u0KO/kLjXvOvP8VE3jQmT8MMsUFX18veWzg
dqZOZXcuwuIN5NDh4pzs0bNY98zvGU+D6yj7GvGv0BuEjwzUPecXaCgAL+EwyNO21vQR5EmEJvmU
uym7eqDsX5lW4nE191GejiegcdYmyTOM4GhFPgyrPy+6SRiGDO7zSmQTwBYFYOtmo+mwrdkU9Ahy
CL8SZzFWXTEtP/Pyp5406yu5v0/OSa0+FbvYckT3v4sixeiCveAoXyhCNAlI+xmO97BxIR/9mRW9
i6o5GO/Eeh/40v5Ct77lWP00534p3ed6gcMlpWzRgXCWO/4WGLx0Usgv6EaaZUYrF4Zw4X2pmTK4
ZUnuBdz5Sxh74eOIywWxt7/eAgSuPVPYllVd0X5lUnVXQYhQVIP3oLUU1wQJ0msfQVZ5ANSBgBaq
5HjrmG43P3iqlN3qkjSVD0QjQanodcuM3+FBU8zd61EgkHaHYY0qSSmzBrKb7wX9nAkjg4Ua5RbI
Zgwg87hX6JP8VkBHtVZ1y2OHrl7cSCisysB2cCwXsV+oP81IY4A11MIhf8ToFmJWhD/LZ6tW4yVm
F+fs1fsAs9kx+Pt9GUOCi949nKElaYlrZQEVtFTq06z8oyxLUIVviaeuWX/3G3CfYIRathFLGR02
w+R9oymTrCb+E8+8HUfnCvv1A7cM6UxcWqAva6QMbNWJWbgLBDQVX/REQ5IDnnP18OwdBxyvoYoD
pwvq6Zsz2HRc47KmN5usoqwg6Ad9e88PKwccz255KSmCGaR7cIeSe70Y1ISrbXCtxdnJF7tMC284
YQknhTMOHT34ksUKradwI5m8RJFn/ziuZJfEaCBnv1MS3Pwry1yEy+WsmN0DRjOpDWAV8Uyj0wCJ
7ndMJ1O+q69Xs5oAHVK9+h/QNgbBvm7Xs5tv2YuxkHie1VcW/7jw2mMM87Cmf+VST02vjF6q7D3e
X/PhUGKJR9fXllSqDzYJoy4t1G7RG8VMEFG0P6g8kJF9pYylTPs1FrcGQsjIXFXDxLIhn/2lEIt4
mTE64/PTkQrWmoXJvJcYGfcTyyA6CSOO7CkL1s6NU/Xyy7uE4nPVNjN3D7iSzIEbs1Y8x0xzPu8V
Xst9UTnPwDlrdtqsHJ/E2CCUOtg7Rco19zcWnwKF03fsGQiB+HetkSVJep+Tl5NfEDkWai9/49FY
Xa3AGfiCqTufopLM4RdQc2KifjDw0QtnBnPhpUQSiEA3ElCVOhVbz9e57xRUfeNsgHGbDJWaLE/L
ss+aDBbiksNcJcDN0QbZI5Ke6bdOwyeczRtuZKW1S7JgMTrO4DoTK0nNwUEbqfhZXCvxxu1A8cR0
mHZoYaHDNrWvxrHuGemUjehIpDtJxbW2Uh4jvIh60btDJ4wl51rgaJNU5w+SNue4skE5THZjCMKf
aQmLCrIteW97b0JLqONH4SK3UL7vKrXOKydic+/tjjf7gyVKUkpZ4hlN2YxSup8uQAvitNo9UPkm
SY8AAHhQ2S67cbL3wKeCBY5dQPWvyzgo4qHraX49rbYBtKBNTaBwI4RH92NEcgtoVzPHxPr4Ue0G
08anvPbT3s5Y7KL9rwrWynuc3fEHPtCE1FvTxjdQ3qmN5F6jQvVziPUgZ+D4uMe4QjWwXjTvdm9k
vxLxo18/BNjxHYyazzMB29Kq4SRzmQke+Zvgke0gKSDKX2ZoG6y2AfEYnyvoTuLoqYFCt5d4T5/G
VzHeEm11Mn+Js+UQuESZgc44L+8hRaqtSUZ6or3vn9drKZ4lFxCxblCGmABKMBv+Id4nydqTWxj0
Jzf/HGw3JacTAZey6WOLfHldZFQk7jDYs0RPxVdt3ZPXMLYhQHgUknOg6S4jbEvMA2VZMS0fklis
mdLvysQRQGjL3xR90hYG9NoLBsELnRd7egCRVkmRrsMH0RYxadBd4R+INxq0VXBb24US6H5rqxvb
8G2kRiNRRGqS/BBn5DDMVYdQ2FBUMhwgbI2jo5T6P4JXzq5BgVc+ROdUgmDcKachYKwLeZeqObTc
AA9emA/UYv+P3JY/VcPq6vh/RSelsZOmvvQ33yBzr/CHv8jh7FXZHTN1xrtnCQU93IWnYgHcr8r/
ZbPanCihiDJSgppEJLC++y+deibawqnIHFauhdgJ79MbOYl3trNBht4UFglMo/r5A06awKnJO4Xf
aT2Dy4MRYxdGb3CChdrru5p8uTbxsx2+bvlV+ULbEqRd+HrubeZ3Od5T12Sjj2C++sxHKhXqRZgr
9u96yqjCLJb74Q4jOc5SwAIaivSC5ynRuK4uUIqzPQDzFaLc5Yxr6BOdpU8CN+qduAn68XI6Svyh
Lzlmwr74AKhlLmx7uwBzMeVgKfnEHhMsG+4sIbdoi8MgKtLXd4eU+8d6HFwSQwXLlAc3+gDa+2TA
Ds6RjbT2Lod/VIWkUefYSpfkmruy+S1FcWtPdrI3NEIC75mkJNOiaw/2JNYJbNdNkJtmGx9eXEyB
jpu0wwDCx3MKcUX3H1sSV8tzHyLJcJSkrOV/EdRP/znSalgrvy+zBEwvBeiySM/O+blg9+Patqn5
h4An9aKCfJNb+jmzc+RoRFtdxfY/ctsBXeraQ5oxx5vJIFobk5NsjGcGLKWKKcjuixP9G7k9ZvQ8
rms/ycLRXa0OmHfQTtz+gvf6YuxQu6zbb22dNFcPBdcIrbPVOYIk4ubPEYGgTl00tdqw6bv5YfiD
VqUn0jVcG/U9aM7u5tM5oUhk2wDkv+qzaibZ5FiKX3BZp7WXZ0+MegQDlnCqLyEA0BbYM4vcVtCP
hoZ4leGGd9foWw6LDEwpr5FYfqcCfQ5gdGbTl4FVEX9X72KwkZv+KulpQc/mgZXtB0LuUezSoU+D
qO1wT6T1rm2OJbMkmDxNFHg238kYKBtlTN8fvwFdnZm81ge0N4AQQNKkKrmDzSndpzCKHBpRaaRQ
e3xUsalY8HfO3vYpsjEPX2sjrp3k61sGmaQqAyJ9nSei47ArXqMViIfjsNZHRATuV+SSYezUG6Ah
N6Zp26FxYUDmaS2ggSkQH4igHcSM5j/7Y9jh/heQkE+FaibOt+yPDKpT6fE/SGdoi8TKmmkOZDh6
xkChFHqSoo0sTnuBE2teiN8mihB9P8bjPZYRWoR5wVnOmM6ajA3+TpbcrlC3qG9BZJYRr6pgNqza
P8t4IHfy1sbccVxYUVaRKxxw3ORWmRh6s6vdTAVd81DPo/76qgd9N641L3LiJ6TP8Do5hwmDadFZ
zY52s5rlAjgNBY02voiYPIcogdxxoFdsVcTzvv5XIlZ5fmEqboddvALYl7LGYJGBAG8HA44WR2Ug
M4R3SIhqUrlYZSHtIiQSJRLbJhs4xN1dBM7k3Pz1rSx0BzeNqEZfohcbGdyUvZucYSUlHmDl9VyS
fLvPInUPMlwhNycGAIAQZcuBF+Tg3JNH2BnnCoYgdG7j86J0R3EWoeItNQYfEwYWwXG65Urv8DhW
jaehhBzXkhhmQ4fmfNYR62EQWJChSfU+vlt4oZ9z+udw2Ncwl9nWFHwUFpTQlPxg2tvQm9HbVnZP
khpODKlKHe3V2khuKYOh9EQv2S1Rr4kQnSQxpp2t88hSDEPRCLUZSEyx3sTrQJcBm03V69XqmXXq
zwVkTGrogNY7viCTBo4StFD+wKh8Gchb0xAgle1+IvqoSqoZANJsHKGQ+fnp2chAsNRZmptrsjHg
r2kpA7iHN2aMsUpi1BYIWm0p6IYYhRnGIfBA8LuCSLOsZf66R7YXKNK/hdIzfUCi040G+bFJdTKp
aWmmQeA185sJy/9RIbKtiX2FtAUjUQMRACaijl5SgzhCIknA/7gqbAUz488DRiQu/elOmiiiz/BQ
hVv2q+Jc1UHxmCWVdrGgU63l4TeIZrgf/9o5RBwe7y8xLQe+XWrlwvb/QUZudF75TpRcq/bL6iUd
dOr5MgAcS6AsOdcOXSa0MSuCtBWzgadpFFO7Up+mi9zfLWQ6TkVpcSUOucEy4gOBGHoCelAoOdr6
sb9d0i7fiztt0/9MqJKA/l3Ht2iEZh5hQt7a2Bhb6O4tnkAUqAP+edPLKZSbymyv/gSvZDDSc1Aq
YEaX06VAtUKA7ARddb0H8q2QQbCX5pcTxKSkL6CiN9tgQUmIx3fvUBrIq3iIxVBU6TUWO1IbXt4+
czg+f0wfz4aiJEvWnZNkCFAGXMv0vI/7rZevfOMgiAdmxYum8UzqamCt5txJUtb6w/Ou62hyPr4j
/3o/4SK9iDqxmW/C0SJUcw6EWZuzUNqF7MyKW0Nf7vnwmHUZEhSKU1N5KPwLiNDM5D9Uu4vB3Llg
ZwfD5SeLbKKPulLIuCTrd5AQ7HtiOlYppE2GHqBE1eCDJ0fuLMNx6nnOJHo16C5qfxT7qaBMlEUL
YyKmlxrT8hv8ZQ1ENmWgogPpiSI+hJT2o66OrCyMQ/b2YBizDsbI6G5eXE+HEW8a8k52pS5WaXtM
X69+nalhTfNQ0VfnXqe2u4fFITSfphqzqY5NZsRmyEvLwjxPAWujtQsK5HKhBF7E3HGhxlendo+0
woYWz0SPODdUp/V6al9gGaNDdU5VTNfHw7NyscrlyDF5pY/9hkqLmUF8uA7HCuMF0wfqpotL2Fma
6kQDX7J83vdrhLV23FYIN7BqNYf8GQVQsSZKxQ5RvhovByYkfAUZO4CvG9SKw/eiu6YWSv/f4hBD
GNZNcfgI3ZSJyzREb3ItVsevnoTD8+G6KThA/r3eaVIYqc3TzxfnY+Uwc2hEQepAJqzb009Iqnsm
45iwWc011HRLxUdtfOyDcS5/AObmq1Uq2tbC0ZhjSjNR8ypmyRTjL4cDac2KkOCbFAY4YIicnLML
gZ2W8TvgF2thVMXzvDwFTFmJIl2Wu5/XY/7S1iqui8lVpeq1fSqHjteGF4WXY98l0aQ7QRgDNBGj
H1WaYHSZCu29Yck+r3VJ8epnrF/XkyhFg7uljg16ZpFHgyNuuyqkr+hoKz0jE5KwYi6H06ma+Hzn
tZsLYAxxj2KNjOtW1+FFEJVbPLG3xWKESj+0zo/HG39BsaibEO4t7w0CzfIHHKbvcFd/OFhObwuU
OeqAZ/cFs3VBmQVP++08rON+XU9CWAYAUPHcw630LFHIoQowioov1Ft0x2yv8Z20rYcNeeTXPf3m
gzMXHhkcF8p00HEq1mm96M+TzGnNbRTzUjhQPc7xOTHXGf+eys6MaM6GmsyU4CyBIrD1rBK5Sf5c
YMpV1DuPDIrt87w+gklWQcPo9L5qH6omL0s8jNKe1uP1Gsa3qtT88xJlHVucJnlv2Laz0cj1w/32
LZMnGn9yv48dfOMY9jmrj4OhUN0rvGAZ34rvWst4A117U0D6cUcpuTfmgP3gEo8FMYiH05YMmecD
KTqj33AKMhJXwPtP9WRgMEfviEq2huA0ysb7MAxolwP/QApyCCG4VSxNxagmy3m7hr0cbxqvuZr5
hBM7S5S+Hqc8OdVUiYsC2/8FOsIXym386Img0BvPZjtZLzRdD8mJyduUqzA6HFfQWJMzuWu4TrKN
/R2wNM8cqh8x0fJ1C2eBEN+0+skY1j9FrboTpz5OVKW1sJpENGpQQCdfAP1hPRIQ5cq60FubdEYs
RmaxSwgBfq3a/lDovEuJeNBJPBKoU5R0l1ZkxaeqeBnkwRDct15pTnIkaZQ6wTW5mwilkoCyDPIe
DVWiCofwJZSIDhTlBaWQsLHP6lfnB0aPClXQ8Sy+3gveoTJsNv4UyXRHllhnYV7QvI5pclnPnIbT
G8r0ING+Bfzq8vC7oMRlWruzMDZHuVQlspYc0wqXdw2oO5nWHTWmsAQzDUr02iXMeqf53qendBZO
PWyKu3Rj4m3IBEFktG3u5klR+m0GGf0CdPHLOX11G90OnNMhsQXzLzb1kn6kJAK5l1Avm3Hf/fZH
WIwP/Aev3uRtWEjboUNVDEqGPZ7VauPsbdyrwcKZk5tNesWWpDx2XUkSoneh+5D/Kym6BVGMfX5s
1oHJgpYTYDLsMOE9NUNu0T7sVTj9jL7v+WLbD5/tKdMpDB5DmO/9midVSlFRtfA33a9MEFQQSoJs
wJ3uN1K2BEav+anXujD6O5Gfuf0TElq8NsmADZZPQSWKm4O1UN0SBgOY0sFs8SnTkVuH2iOV7LfF
89Hm32j0bjBi1NoQM5VU5g9e3/fGPtm2CRB3mi/ayfhICbzuaH5rbzlSkpaI3aEBRV6Y22wJ4maA
H41+JHgPd5G8SDQB6vY/hQ3D8DfUpJu8w95Gp7yOh24spC+Hv7LZUofzBftSkk1XiAs31sshFwdY
xAlkw6QyO9HAukjdE5UMd0Hrq8K5/BOVVs4xLBXAk084Bw7imCyWHQFPovAS8yZP3jmcyaupowvC
8EMFBkUKwCKBz3DtbRHOFT5+AZwd0u97BcS6HH4l5/jQ4GLFqY6U9DnXro2Sxnoo3H1XC308j4Lu
0iQcJnmbivb26noQTi5E6Ny5d2GDktH2iD4dcwBAvWzfE4MawUnSvachR/RQx2gCKhczr4c39/lS
7DZuEOFbr3ich3VpT48HY9E8fhCJDXh95Gg2s/QQziBIbrWlgnftHTqZVbKsFX0UL0vIrH6oTa8E
jaUUp1wP9NYlR+rzeVwkBj2LNN7+J5oQeetbCQUx3dMocuZylNFVzn0E2FUDZhPWw5fiQhfLMG4l
W9i/7sQhTmu76ksQMJCriVEHYiVgbI/6ZehlApJvpnFOnvoIScapeIACZ8f/M9qmTeT+8CkmGILA
hrIQCmFRqhVhwR3MzR/9yDgtPg9PRRqKdzFbhcysVDIHMd6vsGHqZl2RuSdxnhNa5ycwJ7BqkR1i
NbF3exaqZehKXFX6ClICp8toPxKYR+sam8AzPVMNKm95FwH9aBu35wTTrztXMlXYjSS6lYpP3fqE
PtnuF8d5imR+s40o4BndefgAvU8FV1EjDY6iYhUbIGOZwKtFMXYfp72BvogbN7sXUpMmF7IU3j2t
s2moPlIHL9/Wvc+8TnjsEqbP+6xGKTWS6v7FoMbRtOhioWZicSBX7iRiDczKxJNvT/HpwOW/y66k
fvwyGMslCRpgvX2N4EZazMEI0EMrnC8FBqebYTFie2XanMGePniV9gB4dJw2NxGeXxemNxVYjo6X
7KMYvwaWgEUJLl4Pg7hhqqLgAbUlho0J9z7XE0un1nNpHx6cmXtJZAvwGHjB9Oy2K52StkkYCsDj
XX6EDowp9Q2onLnQDpFGidv8Y8QbEVsBIqezB9nh5BzOUHqe11Q6aU6nOSMEx0V06kqxrykNAqwg
bxNLztrTCdkjvZMrmLG6N/Ik+4/UMgOHxjpWjX3vzNN+xWc6Licmr7lXN3XBvOyb+20mY24EJ2uQ
Y6rSCXbc5mn4uaYYl6+ffHIWAM1XGiT6gjkixkCltgmBK3ksg9hiaKPxY/jdQH8muUTXtpAcCkzf
B93sf8sq57gKLRIKDW2Egjs6Eqdf04Utq5x93+YiyNaVTB7/vbKec0yp/TZJgwkXJqU/TBo0D83Y
l7nQNvhggqxtMp5qngUsJ5Ojm+7/aCpIO6kK5ZnJomxfKzJesMe79pGTeIwo2sTUYdH7KycEcSeP
vvh+sU1sfvkLvxTXwGA4VE79trCuW5pSZRIdo2Xi6q9mZ0dHyMhU9DVCras/seEqqiSw76QFSly+
PF5nphMpARsa/fVoU3HZHnW5GelDVk/U/PlC9NbhDItJGLZcaS4llBk8Fufur3qaGF9BC9u1/1M6
cbeRUVNxjWnUZXviyZQ571eWCQO90bGIMmbMw7qwccnxnpGNUvNmUSuZq1hd/ejSdc9ir8WYYGkG
IzD7VWStfR/tXyFjbIc+caD8VKgdix3NL+9RZQMqMCo2pks0CDaLJo9zqXA8TEqSCxxf9kqym0SQ
y3DSwxbB5kgauHA+3/IQpLoiB8E2oVKHZ1HYDPrnUnwQddzaiymk84YeJUIw7d9CIYJtBjuzWn4A
SFQR6MqYPZ4ZhhY8M9qCE9LldBir9mG29Ze0TfUtH9194DzMlRNCU372jYXMULNlH5knmahAe1z7
UBSb1czUkoBO8tlZGKNfCJc0rNEQ0l0o1zK8kP/aVZ3VB58Puj/tX/+SVuqcBh/W/q091rB1vfO8
Gu0ArjJv/JLuIKwf2SHpMVD6wlfBz6q7v4w+Qeh+tQw40h6tMLLhn+/j+8AKm2b748NMIhgyI2lJ
JIa8wEMZhAZkr3sgMDxEUKxcVJKPuHFSanc3G0SuoSn6inajxoOwmrzBqhp3GsdBKq2b5WiZkoU0
FmfAjWRPkRd6S2kR6fHpAUJoNr87IEWuFvbd6jMsJyOrvCKUX312+cVcwMO8a8VunkrIuDUf8hxS
ROac+zhvcBbZ3fQimkrLMgNJ1HyDjMteQKv14QGlkKL/gyc8KshJroniZPA8xMxSb6FCFwpQtMzj
TH/E6S7PLo4E8j/PPx169vvPswWVfJfO5wjSt83ZP17r1Ndj9cIhU7T5TrqjvbmqgLyktQiWBPQP
5nRu/ckfksyfY6D1qHVP7djrgOF3A7P/0HInZv42HBwREaPLDR7NXUWCTuuotw6yWVbgV0+2gd75
8mk0JIJHJQkSYkXYALYLPn0exVzotAKaHey69Yph5KyF8Aef0n0sm4jS+mVPV6LBg2zO7Fuv8fbb
y9uc6u9HD63yaaQen4kWSQ1oGNYyYkRJjhiGvHe4x/FhJoZM1wz84H8BXMWdw8GgyhLY29FVVnkz
LMuoM0lm2C1IShSfafyqiWPLWyqA6/oqJaVQ4HPTi8pJ3h0llJc3jelcJo4h8p7Acofx7uk2W3/w
WJn/cIxqX4wfzaEdpTj2dQoU0uUHSr5zTta4tOehaTqHrYm6oG/uK1iVBiQgSS6N6FVKuq4ZmNXe
kgReIvBm4BwuBfeltD8d60UGjEQuj6anqmUQgDnGcIsSaZvUjDWtqJIrHrx/28HYK21ExE98/IgS
4vT4MAFIpnUYs6Q8Pi/kM/JsU6fpDRbC0UuKKjMEoCsBfB+TOEEGG/sRrH9PvWGwxNu33k2Tr1uF
eSUEphbVukO4wwXvxs0dvl7VVNzBPbwncozBzS564e22kh9bSG08vbQUucNQ18dBTE4TCPXHMUx/
jBYL3gzDJSzVKqe/x5NeP0VxJspkStEPFq7+C4RAGLslh5g2faKXS3B6/MF0dTlBwZuFPVVgrjoK
LJxUXt9bgRHoZk3lYwcDh+P96+S7ITbfRCKfsuhCtepYb8CiUOSXFZQXxQVwBeQRX/7RA24G117E
8VKmCi6dPIVz67z5XAOENt1og0Vpn1V5eXgskv469wc5o6XrR3DlxOjCujbmhrKkr8AYBX0F7ny3
NDv3yBDFENh8RiWd8prw41t64TQqYZZmgmv3AoVpjMAQKXpGnmuMed0qOI/EY7tI2jLhke9+191g
k8wzsjOG/n/fHmyaMMIF/SLdCmwbhn3M9m+Kfp0I5rLmNwFWTsSXKTwpChQnQ09G8oDajCiJGrId
Iap6RuPsRmr5nalzd5TNBn+Z8O2PA/a+WHSi4+YSxSb2xOlQ3zwgyj24RXjOhpXT6nQUHuQUfRe4
wbRTRGtbFV0l4HOVzH/QvRnquDL3roGwYCp3Gub5p9XgFLb/Y7M14HLOpkGfC91ntIza/O7uVhEo
l6sWuxtH33LpBg+QVG6VW9K60JyJS7llXP1utNfQDa+K6ybHwjbbW0Hd9AitHQzyjUhx3PjTbB8K
fX4bTsfNN3I06m5ChLPvI+PYfz5ugtlq42ZVqDj7iYmepP2b9j10IZ2fQJ61nY0M7d4nKe/2RrPf
TPuvWziNxSTQOxPzNvmhFCLLHn5bj1q3nAurTL7+7aeurRtBAGpQb9jj3aoz8q5b9C1DBypfH85w
K7j08htrg4gb/FgEuTCYKqvhs2hPWmtq3Ppe9wLmXpnUgsvqdpY3wRAQgsALKfuawn+8QTRiy+YI
OTFRR6hhFyIGAUfA51Od8om7fCWd5irif0j8GMYOridXLVtX/zsno0RpviMoOv1OYkcAv+IHquwj
AeTVQOhlhLKcU2P3oAhTs5PMDkmkSjmtrv7p7CFP8VO0E379Qaswmjc3UBhZESrtg/XCI3EyCpzI
YknXQzJjXLGWNGFJ1SJzg94MzQQJV+Sc4prC893bl546Rw3Mb5zinnPW9wV148Chh2E6vokCvH1Z
luyvgXlsmQmnb3j/EwXeqDbGe2GlZzMB1prgbyuIc7NnujfY8THMXO+YJ+W1eXTpSQJPi3wKEJes
cZJx09yqQOWQourMn6Q9MQeW8rTs60oJ+1txvCxRqoMtTit7qAeTMGZdBj4mW4IQiimE2DLr+DAQ
arrZmIXePxOfikcz6pwxvOxXEduVkU9WpWaHP9nJmdOM+BbicY4++gLea7D3IWaMP1yV5S3ty/gr
ZQK9tYNSSCRqPqW0dohkDUIbdIU5wg4Sa+o5B8RJMwi/fXc5h72GIeIwP4QBwUPnxUWCEi/iKxgw
K5y65Nh4Oo2z8IswriX4RBXM6syWAMtDE1aOeqqPE6e6JHlddCKA23Tjx88vghBrmo76npVWDX8H
TSKU2lz5ZQpzbwa3weXfU/DXwwtlOQRmyB5exZJ7qEFRcz/DF1M80lWd0tjI9jEiqFwrxhwIaMhN
aVJRHERHICdKeRTp7+IdyCOsoQ0619VlY2w6z8MrJCUAT+h6B4wQhaRLkho5MmHgTn3yfT/77kvT
/T+ym5/w+7MtAXe1DdXbCZPnF2MP0QfTCJFrasaNIR0B45qFMmrze0g4hvuIq++4RyXrxJAv+MAG
D/WwMAvHpQopzltFKjs7tkcyvVRFRh88lWCA+PVGtB5KW+MJGCTKqWrowxs6EBwY5Nw7StmTD1Ul
eoPrh6S9WxkPscdc+PXZWY+dA8pqh8wTe0kqyONJ5pNHuMWpFHIzWO5y3FUkNLQYHa3FB32XJkr+
DJQW9mtU2d6s4YW1R1SwyBNPrI33X8wX5lu7jtPGQss0iTqMsGMoZtroRwaqHBJrA4ZeB799LM/Y
Ev+6GTmD5qkJAaBUby2aLv8CLRBHmu2e7ri+hiMEfqQSIWFFzqthLVKHcE803gKyF+EgooEFrC6o
D5U+6czog/xp5vV/4jBzbiaVsRR7xPEx+k+AUiDI9SBi+IW3ozLoth4OpluTNE3jbqKeJtSQ8+9J
hVwuSLo5vlAIkXPbVqRM8nWeVOdaE697Aa3EDcaI0/CM6i47oF34GFO6g6AHGMHzUseKSSvPmGQX
78tH4xtn7ava77YFB6mTOFVH7cDbuRJ6YOxRbgcyt4VTqmc/EWP74C2TtZWoHb6ajh5KrFtEoA0k
7bjHvFn5X7znii/K52Ec+TtFTNqM+cYyDXu7VZ2ioU2ejlBWcrzJKdtcr67BIENv8Rlg9U+Ehd1x
DMGCc+Djn3yaDQcPVWLQiH/FWUX6wU7JSva3e2mKIl8PNH4fr5K3nuQ8BpStbysR4doxVj3D1Ikr
nm0+kNLeOatFta0YjUyeMqrwSXtJV4Xf4gnReLSxru3u4zJemHXvxeZ9vsbfJfRRDGX+zK8Pm2e0
dOBJZ32pt7DCqst7z2CFXcUm8PWJsrg6nrslCLEwRIhcqdqCZSCM3Lc2nIZ0QLBySHtFjdTuNVxY
bLWq4tw/kpFhYfCrVZVK3nJehtgOOiYrRiK5kZV1e76VFWygJf4gQNU6JY805iXT/gZKjXelr2qI
NX3mkRnrRllm1EU8yp0sWpci3s7Sn8rTDTsh9W2tR4BD7eKx8QKZfbfvmPN+g8cJEo81gprlzxyU
bPmXggIV4Wpm8zoQUvQ8pbV1JTOhPCzAMlfWsFJTZohBF1yh3RTkpygeh392daGdaf7G93JpisKv
akwzpH9tlIYyuEW/dnyUUWuXax0ze/Ooj2FObIYEHHPN4W07wgCaLRHNVF4sxIXnDE6WpGm9PZ0F
vZXEUKMcUbMTuIDoO0BH6pr/fhSYHb99GXEwRH7kMMNRvcyEa5GC1XCxmCNKbZISirYJP7ueVnsC
+ZfbovmqQM1KywKAKfsfO9Az18scuq9bg3/IzaZKfYjWiAoK6xtJR329AOPokG7Ilpb+L+E8Ugr6
x0w8M6ZrlHaHPuSIevN3+Cg8fNoBCYlQNAHmbI6O5/kXxzBYfMLh0leLGL01+SpYR8FXsL5cGBoG
BQW5rU57+0+dzF7D0saoEUzdHh5vjPNx04S0NTml8Amp+GtgNQRwZvrCGe1DKpv++4o8GpQSkIGw
637i4MPdhLQE5bejwMaGbJOhl45Rvue8h0Hppcd/8wOUROSPPYlTN0Si5s/zT4k1yOce6tFNforL
k7sKEwpRFjtYGILufeJrk1BlkSGTFL8iqrFdaY8WtVu5YwLoLwcmprDROPVfA0iMYYbUIzZZz8Fv
v/nxWtPQufu0EGCkMMnmnfKicVZWQgMa7UtygGhCtDXd5fBv6HIjS+yq0eniSBvLDYlSQwmoHQ74
MOBfjRzEQCtdSeMPevJl2jYDkdSRDhrTADI2QCjDFOO4ePuWU7zKTrON/kmEqGlO01RLYr4yTm7e
dMT6NrKQP47pwGbOPCR9riMv4GamrXwLd0CmNxC16D4D7BhvZDqUBTqozEF3XL+aWY4t3yBuf2M2
QYGtKp8YRglH4gUev456lhyF+3s4iX8NfZi82Yc8auX+hgSaXH8EbKphWB4Ki58zwNDSoGsC6M/y
RRd6uTBv9dE5Ofeefn5pS4R/y5SAyBZyHzZjvqoU7jFAdhSy3CRdL/enMViMHM9dQOl1HvMPvAUo
ryrSx0PpK1bPFOhqLnGAo8IAMLW3nwsUouDekE9yeGHNbxVXtB9gmcUn2+MmgNzNTdzcZFoNr5Pj
mUYhld32rpD1tiLrcx/L0dsz4Jp7GC+/Q2oSMo3zWNdO7RrcOI388YCyQ9NlQXFF/hnycONE1crC
Bwhe5zvwjyr9XfMBCdVjspRNB3+CLEijbOccLH7zllkt2kdICbzg4TplJ9vhJKK8UpnRRhNtYRwh
ClIgA/1Bz/oLTvP/D5MJe5Z8LFjyO/Uf3cSSd+0HXGHyWn0Dcv6UZry3ek9Hu86u/wr+o1HM8FO0
1UOvK2+JvYAQR0uPSTWOLNklo/JEYAw4M+vWVa1b9A1wCy4LbPsYmpbkeSMFZ1eYQwMJPk4j7inN
CDSbOZxPsv9PVg+OVDgapqA7b/+l72J2rBKIghw3QTlME9UBHzqfSj01R9qdNxGn8vYLkD87IljP
XmACK7tmaXyM09Rt4pbNelhDgdth0tIyzEI3a0G8HG+gjbHCkv11PRBCOmmirG1kX9q8HYLXnGka
A7c8WF8AH7JWsi3dbD3RizAzXvpyhXZ/mxZD3CVGBnisJf/XLqH75snb6YwBUlcXp98PzBaRS7Eh
cxUNxzDod6tTbY3ReDqLeWMiGN1GBIKil3EoDjvPu5nD/h9e0+NAk6q+qN/SCGOMPnnfn7cy48q3
MIVWSkyKa98TMO7CiwU1tiwNz/iDLKCZThqX9Ua0b5bMMywp/LPew1tzuiFvxBxWc0rlCz3pZ20P
NFCusrH0sBHje9ahyDhVT93ebLSILsoOI02DDY//o6RzvLH0vIoPSNHJF5gnjjfOFXEGNJgExYS0
sOARrVdKF5IXRgGb+b61rzqv78T4GOfF2rJ1EB4gVJzk+I0vnQ8rKVTFINqQcAoVwI3Znw7KqzDz
XgiMgGlTCIgrQRUqVDRLLcPXY5yqKMRmKriGU8JUG+7JNegs9Ttr112k3FaENIwD3ymcoSCIIS1m
LtFfoClGpFOR4qbTsPqWTYEBsCdCjHH6bwyU/SdqfPwsANMUGsNepvNTdl3IdXf0pplDEWeFgmdb
zJufscN1B7F4aov9LeeeqYryXd1reiKiArHkMh2Xpsr3q91CLNchYJOXgBAou6xkj1gyQ26Ko8IL
DIOfSNWHXHZoeLntGce6E/fbxZdD5PfoUVYqE+9hBf2g7VXN96Ix+H5D7I+cJ+poOBl7WBwNWBe4
m8XCrsRL+vrR2dWGvC57l27rsoKlnx6hPmXtskKoxf1vZzAK7qXVqwao4IyHzqsHWgrOriYulMhI
W5rz1nqRCcVrLZKKDS5BWDOskrGNO2oPYbpCMFQXaF5ugOfSUVjmTVtZ0uIW7gsaW8I0oBaIUSH0
lyxc6tEYXizvapoyLRUsZnOsRGJljntA6hL9FJBKgXkGGNxuL9qXaziVh8/YXXf47t9sm3IowgDE
F5ifYL/yp3m47CtAznIs0vcBQAwavbFShAHVGk3DVN2SyglDdgWjmdQtwebVbINib+M28odFu9o3
NL86ReFiOq2oidFldip0eJtmedDYI5U/4RIbwXpbrj1ZQOt5aQYsS2FR/8WYKHBzrTzcwm6HfpoP
0ktHKRYVPTnKfTseN8IkFSuUKfVWzErvw3tJSLQ1Ln5Olmrfr1f0AT0sdww4H+qCjvV3OODGyaH/
v7N3kA+O2HFmE4iG6nxrBOQe5jbWiAU/6linkqg69Rt7css+bcRxAxuGMkOUv3Yxk17aandkyiSw
OFMcHkXu/cwfzNH3FCFpgD9fknvH0/VDGS+oDGh0JqyLIaZAuX43FPNniTU2waf1Z81cY2xWuYAK
ffO3mwbLzDLUSsDnwDFatlqNqNDjzK61t4zAW8Zb7nEuVzrzykopuB4hItR8hfOvLWK9QWY4PBzB
fw3l44JaLUOU/IHz6tRjA0guArXOi93E4DRlN/c8879B1PRE6/9EwqiAR6/QOyZjc2padi4+sXhW
aDf8rQ3ENZMPV5gM/QfoselJgu8bTdOWZiNZlgt79Akw18PrmYCI+VYsDseNETbJrNe8waI7aFzP
zfDK2n5o6bBADt+0NqfXCTRJFfBJ82WVF6BsmUadmOT3aZHO0xNBasAg2WMVujeboBCGFLCD81qB
yD8Q1bCDv0w4Hle12/hZ+TLXLZMSWYxGmcM1oS08BWeCF6uE2GdPPDDmY/1qhEXOiO/ebb5jt5+3
/J5VdxV7Z2DaB/EoUyjbkWYz7h/9M4b44KbNy3YhePG28qi7WDy0AiTryA+sIFYr6PFu6I9iYx6t
CHSwZY8uWEmQqLJFiD5Vo9LlYlDaT1XGv04kF7f7O1z09GieSegXhyRmZ9dwLxcLMuFFcCUjSkU1
RCn/1I+IGjfbCNvei7tJCIm10SedxcnlbSFkZvJhuTGTnI1MDmflCiMfRirx0AgH5+1Yie3hWH4V
q9HLpkRvsUFVzBFZ9p/ycPw7YYI060M59uEoNpXuNTifqqxn66Eg/6sIhiyLOZh0zyAY4E6xDPvn
v95rL1igi9aVWeUTSUJoz/LcDqrfIji+Ei+wgd63KRnAElodBfx41j+fwW9c032ms00TjFKkjHvE
JfTl0ZtzCIWH21w3Q8AjQ11X2uWZrVrIC90A8ub/1WwpAlf7WN0GQJB+n+u7Hyx9Zw5vc5c7ZUnY
sG0ChpNF09Sw1BfbSw8pvnM/ZYEX/+R/dQ4ptnLwdHF7Zke3WUB2hxfhxrXP2XKZu8gWsYRp+N0Z
so9Z7Yra91MLfK2u4YXI0XdtwuUtZ5MxRl/IUUFDNQJsiQokegoDnByQ2v/QS69/UplUDAtcFgtt
fOhq1tVtiCthoZMyZGNXkg4lLulUZYVvMfrDAQNtUyRqRmvoO0Si3nqLXLCMyZ/DOUJ5sv41f+32
AKjgs5G9TM/ikOXP6zzznDB3Bs0iOUG2WsUM1Z+zP+0AO34c480YuSUF8Oyb0fuhhHlvcndLAauY
CRIvmXD02d1qQh4tzYx/7LR7yCP9OD6D6od5NYiEkeZm8X0yWeftmGNhMpog1poauW4gV1YKjxL6
Lu1PpHnZqD2OOyNkd2lImQ0ix4IQ5+i1Q8d+MQxd+ZOcBHC3AZ3LoGntIRXO/gp4l30/U1YpoK2E
fpzJgNH9fLag9HHNLrDarmu2zmrEVoOL2mCUSkeSFQjezmlJ5NbWZYsiBqrs+SaJ/Lk7JgR3R+Z8
rk0JHV6o5JtBamZdxCucvpzRih1jQgSTRhiMb+xSKOZ29n/wH8JnPrzJOySfhKy8++9gkHIbHNp8
tg4hopXe1KwnKBT87sFJLe3SJC3qDxCD3XW7BS7mFPWso6qdqRzr4k8E94wjGkXo0aedTkmLqm8b
aUFhWs6jKLJDmU3WV9eQTCIJEJWMZxEOvlUm0fn2Diorky015v7cpjYuujHTYZlFO1N4OxEtjmTl
04CthI4Kelp3JuQmI18s5cUGlrfzTFsGhsXzjfCRiX/CVHFb6U6P0t0Or0DottD4anVXfEvIsF+O
plRPIOENiUpnP9yRy2wNFvPE0Zy8aTtKd7hZzJlSCjfxNswQSOWDuUheZ2Hs4zC+WtkQk3mM2yIa
d/Fvd7oi/gMXBL0n/eTeCilbRqmn4atjOHeOjbIwPD4Fbv+KVey+KrxTa3ldAzszwEEwlsUbwmHr
HUnT+v45JMaxTk0oiFaDNBVDXDfpu1aQWmbZQtnGKiJoftXlyLl7mXcDeAvlpJo+X1haaXP5ChgT
+SoxeRYNUPGMVkVzx2Te4XBz/eQQYENDu4g+j42mpKARUGz+kaEc1i9vkbv/EyRjT5IDI3im+f0X
qYSytaZZPRbjX3aIToysn/tSBrqonC1QxH1lOtdxeRWXIFvDzMJOSBgrigI936dVJAlNIzabCe52
nQumPXUFc6sBAodyn90v9kS/M1uyyD0YpR/oQ5ezbH5gu77MwBMqmUEvieDexfCHpvZxhO5w170O
4qasXkDZrpWGegDW21O7CQksUA4PXRy2Byzx5WwGJN0aM2WXxe4zrSewX9/xOiy7pk3TUR0DPD0N
Xu6sFZ+tZQr+JxYFljEkkTvy8m3Mtk/Q96xqSfkrrpwzRbGJAbc10vlww3dQul8VG6UVmd8zNybT
QVUxDMY0Ghm9BuXXjEvqrv1Gkz9eT3JlgCQtRK4hh/3qPopwEFNZEQwdE+Up8jpmTq/jYAmXxIgE
8X8fFvUAz33k06/hAQAPaJX4K2FePSww67rnMEXWL1hhQ1oy52tiQpkH567rzZI1KakmDZ3ZXig8
cJ1fjcrJPMbILEbmQ9w/+QRa5qLOjEGYBOjDKjSBCJ5z+JIw5VUfjFI3eEDr5qeipVWxsbdbYQs0
h0brUnd6N0dp1s02EbohCUtSytt1DsqTjjWoHanzafgiczfINdFUlNvVDRkN2DQv+U/2fCW5D5iA
M/sdy79RDcC7IWaQZ0U3DcWI1z4N+HHdrx0gPwIzdC4ucCkRdU5lKi4HSFWI8JKqFtF6XEwAiWdx
q4tiD9BB7KgLeF19rO3SaQmFY5bMSX9haZc7Ydx+aqFE4QiLC6hduTqvWwb3Jtnz6WfftyGB7no+
uvkjt5U/cmZQ6oqbdLmoeM4lm01gRM6VhRaxZ6H1o2VyP4VJnGHRvmIm4DpI8dqQGnmy4rUE1Avh
5lWHF0saPYu+gRb8JN38lxAjLfAO4ZERaOTwZK7e0brFQNTZ2AtKrOL4N+m8v5uHujyX4q8Sfl4C
Zm8NaDmm0ToK8bSqYWg33yGSqkaUREP9PvIhNfe3yM22amIVL1RDvQYqXj1dm3Cxn71f4rc8vhVk
KJt0mmnahCvvfFJtWFJ2eGNa+U2eeGcoI6xGMvb2zkwlGb8ddiZi7wRaG755e81/EXiL6e/T3Tzq
5Jtu7hryysm9vGFEmTOPfSWRRqHVdJEQBKAoQUj85K6cRxNOtXJRjphTnbh9BTupB/G+dz2W0ILP
UDydngSTG4rxY5YeAiTqlhnYO/SivGleGY8PZWIvFC9s6i7SDPdpmVIPTghkqWU18NQAtzU4pS87
Z5d8LXwLZvJukhJlpXlvjFiYAe04/kFMiPDYRi+F/S8kWnPy0bZUUl6rSzUtVq8UyBjSnXIDXgcn
VhrQYochiL6150hswSf2bZCtzFlzj5xa7hiuztndFfqpy5nOuWKewx8g1/yMsSStQ6E0trUslDk0
Cob85fO/NxtGe6MpDwHkEqBHXnhxZpHwzQMeYBTY6vk3vsDhRgQOIxzSg/DA8Vq4vpI+VDdrqB7C
v9Nd1UOA9AlbJbYkK7iAFdy6J/QU+T/dFptS143fPnYj4JOU2WDnhcM347JiqYHASJRGR88isIgn
BwhpJh+yf873QtMPs3FvnYwqSp8ttNJzuXSOuuz2f8i6/wlhJ1sbhsOyZ3soYT7ufj0OIVEl4JCZ
wPWCikhIA4SX7iU5MD2BTz+uUwSc5cJSMtOqUOVqaOsbnizDh/GK3T/MWtemBNa6VRy3mrGne8jm
uyGYxUYtdB1BjVjO/HyIfBHKbB+l4Aq5nfm53zVcCyXWw2Q1bFgsWrvJ09mYICS1QsCVyAOdOQ4r
d708HjuQq7Lv1AOBMdeRWqD64ULW7IenIlYWn4BcqcDcvRGRu8w4vbME8W1MmnuDXzC1hpBPc0TB
Lz9XE/ovYQBXe5a4V80GE5wyzfLzO/2nkvk/hM0klTq6jtcVrmGmJ6j7wpgtxd3RnggZ9zh85Kgu
xSXMEQkv+aSbK7PHLV99XBOCxVkbaGENZ+kz8KnzbBxCWZSvUyGjBUQxz7GdnF0pzUMoBDiFEsiE
p++EZFi9iXA6Ls87j3nQah0oFrnEnVKyRCDhaPAk0KyIsGEOanKNrSleVIHZO+8gkUmxOSvijbmA
noUuKtZ7v+/uuSZApOeanNP69yCTBV16fNfvhXdYeX2KSrwMIm7jJsNfOYfjJc8pMFoQPlndeaWp
KEg0xSUDcgNt1xVh3F0h+JJzLx2irW+hSnb7dAw2qo3O5mDvLfJncv528UzlRKF8smcEoPWT5tIa
301udChD9A8q6RsCQWTEG+B1ST5KHQqBILqJAuVX6zXYO4mjuvFp0AGFx6VTWIBvMids3+ujfujR
PRdlMuzAg1g9PbiGIKPffoEBRh5Vlg+wv/i+zCY8L/SW5I54W5GWMof5S7ID3O8arbBaQ+uHGKiK
2EceZsK84DoYwn7qpRXacLfxj900je8+p1/RUGaPxfZEKp4KyherphfSlFc54Qw6D1nlvFnTDyKR
GuZgAP20kodQFCMGkQq2dSnNwdFvayer9/51H+UwIpK3iDxujwmDlIfNRh/rhOCsSPJiAzYfrwML
vqFGLESkp6yyQ8YQ7MkS60Cq8d1h1/1KRPxM9dkzmS06CvywvThvN7O6g2Sra8xhFAR7/MM0PKHJ
aVW28yBGPpQ6tMWHoeS04CyLWFI1S+EVHxnvomnL4ZRViOEmixhWiVAHHvVeCODX9US2PyRU9lL3
UW12z60YlU1pBFExeDd5Z719ckZB3xZsubE3SfSAgnCKIPlIS4SnlsuSVHzkK8keNP8t8/Q0eTbW
Z+8PQD9QLyV7fTAP7b3lzDbIyDQAX1P9qXka5HhAIeAf/vhflNPHPR8Zmh5HdpDHQlBz6plW9LsK
A3nc7pjOZgGeBUo1Nz2lrk3mYhApYA5palhcNdo3mrDusK1DgKaP/noSGdtXVEzFdfzt9qwAeoNN
mInMzizyRMN4yJF37pVkJ2Qutlnul3BaVOKSrnqPDO4j7J9aUlCMpQbI6fMTId5qD4HPf1EMP3O3
DiHvQ6WjNMIfMjTHkSLjB8u1BWk6L7UTsvVEEarPy45R5zI4o26IM2TP1T3S3NkOFLzAhgfuMO2e
l3j/6EP/g+LMvIJpBkhDxAPibos96bU9nNIA0p/4pIFh5QcTGCtqfJHLVCB0OaL7yJ9+9QEsmdaJ
9dSYZaRRgL3PlQ4aHVL2X9KOuavr6GjYrRkerU+wejdXmW/3Fg7nr3t0Bs7hODc7kM6pWwdxf5EK
5vlhBXYLEZGXsZ9sQtSlsyEX4AjT28zF8e4tqie8BFOGTmIzp8IKAK9VD5+f6HQG3b4LbsuCHC4x
hiysZrztfCpWTRCnQoSq4o08cOzRqj/Ar8JWCvR87iJZHscOLyQHxZXCLFgmFPzvMUnsapuG2jde
Qg3ZHiLkLrvIvQnE31MRHkE8DkkuzujkHkaCkCr9agQ+aBh24yYWIxRbo82r0q7UHFzkfbKWjbef
8TYvdhS3Oi8Q4VugopIbpxgi19H84xPCb16fqm7Nj48xXi8HeoggPDPcMWQNyC2Ol6Sx2P0fJk1L
+o1gV4h7qfltr6fwwiRYisbo6yi0lxtu0DR8Q47I7GhxEzd8r9MgHID7xkUUZsqeirlu3WoPO/AP
mGhsBlE+/7YfyN69Mdb8wwPsEqo/JqrPfKeOjlYzfuimudKlYLwcQu60AFuEz8lRFeQPP5U+GtJX
ZdJFyti3yNvTH5oxc5ONZkN6E1nxWGPnLACU6vPwLVSox7SxUP3V2UecQ1Y61UzZLQYVGhLKgovx
9Y7NScsBkk5a73HOCIrRapvk1r8uYaF0egGRojqOQTUlNF1YJoGWh4PitNAlnAjVzn5z8NQBRY9r
H4DOsVPkphs6yGfuuT6aSbmOk/mhTijMJxlFbVzmrnibH66fbNZPlNdq3Y95nCaqupl9XB84w0XD
3Bno2V24dCtu3guvtX9LWjD2U9XEEi9u2ZnC6E7tNGiDm4HcCEslql4FOZ6s4O7QM83PFl5QHDmZ
zcZ9SDWG6RiYGRlY6H8dS+zcLKc3L5ofZpnBjjf+/fGJ/r7mGlVDzLAvEFa8lZP1bubN4mjazK4P
FzK3otLfFbYVjjAjQTCCMZBQRc9q1oh29DNpIIiShiPPGKy0uYX2iOF0nmDOqoapMg+VxLYsMyXo
3y7KLyTd+vWDPYoa3su1bNGNnaTlrkanLXIw0xXZZ27YkUzyBiZi7VandzxJ1O+aJ3Suh4sXPVFC
99JKdEOkMFA+ZTJlQtJr7BnqF5NsDxfPem9Bqzk3Hkf48JrdbHxgRWuG/FCxnRYBpD9LMTBqAGR7
O8glBPFa0SbylvtgKjx7zjXt5ouwNt53BHYFdsZKK9L++uxbXUMQaImwgkRLuw+sguE/Pg2fneF+
q586wLDleWXdqvW/KbVTk2iqkNXC8a1ZK2PpyxNv9rzsdOtjPO0ukk+8zjyV3WTU2LP4xB/iTsg0
FSdWmOsowXaASYFkkYfacPn9GliK0R65P0NfLzaAALtFJPOKYRaKma9xmIwKzw85qDZNVU3Bp65c
vO5CJkP4Ta15af+kuBwftsKyIBXhHrsozbjbWti/eURHLEm/XnskaRwyMu5JTE9ln9fi5kHLEBmA
1typmGwRNyRm0svYhifIGdLH3J3s+mdMAYEMdQnN0erPBfLxCgmVH7/ZOu7hv7mQBHK92tYOqMmK
Nt5LXjTbfmoW8UUEQIhXa/uKXwuJkb4FHkaBSS6sI9V6DoO0ifkbaCrtXGQUqQ/9ApCka83FzweV
VyGcFvP2hg5OgtjsaNjQ+a9C0/GBN/HjYvIFrN87MW9X75EaBes5ulqlqoLoSS3b2XuMOUrqK7yd
utSV99dr1kgZuzAuCLwWCntIYUz9FRIhtI/l+prvy+Ci1x8pw4CISB9d3ZiMcPQpMDAJy6ITzjFv
Zs5Mbi8rGKYHPjftVcowLyufIFUStAi/5wTEE94wzznSZp9Pk8NT6Yta3I3wtuluXAYi8jXeSCJQ
/JB62M32rikcLTZMIr0ca1ZQJlvxhLp5hi4Ov964jsCcs8u9h8WFJUbWV00e4HImf4Ze/9QlkyHn
B/3vteYZ0wNtQ8B8F6SowVrq6Tt9hwyi1Wp++YRuQd4LBb/b+da1SSH9sIejZmqeYyjXYc2PjEuH
GBJdQpyzqBCKgbeC2a4FE9qTw97J5ZqjEe46E4YK6SYnF8rVzkQqiIErFD+JGv8/3ziPO/g7c9CK
EDy0x/6WSO91GXc9b+O3/4APUj1e0csSaGxGnjxjVpv1rql5QXjG4IM2qJd0USJ/0ffwtwHllR3/
8O4Pp/COj9dtYYfvA4t74DiuGvcWNSHwL9/rqWe2e3GA2UEJLqoLPvsuoAFcXAmDZGQSCKPrnk8c
9SPCquY0jlYC5oXQ0BWIeO4qoTVXYU4nk1Ui/MXqivxexC6rRhSl/9TlLaxHWL0wTgloPoKuJNh0
5caCTcvpTQUy14DKadF/DDylSGUVHaJIXRXoo5TRFxfYa59CZtgJ5eJmSXcpAh6LjrxXxzf63Dbq
eyJ21UPVXM3xfmn5RvFzVqdQQ1S9Esfmh2f5elvdA26tpcOQe/ePTzWXZjOgoei9mdfV1XnmhGBT
cueb+R1WaQDhaaiXVefH4NukxU6L5iScc5OKtjJRW0IpACjL63xVg7Jlpz6EGsBAfZCLpK/kilO7
RYZY1VM2E+7PoyAP+RtkMLeqXkDiZ1+2DbI61fc36gxrEFDmAdm0dywRRpSVOY++jBJEVC8jIwUM
rn0shbgE63T0a2z6RrsZ6sgpTb4QdWlMDbr0NtxSnYlTE9+ILSC5/vxQhbNW8pYRmFJpWAMySSWc
ffiLmblNS800S5CNmi1uD/pOlN92zFJBDkcrz9XY+8magxCn2CBvmV07HqtO4sJXE9jGFP31rZNz
TEP9MtIGAWjR7upOqNBypI+7Er3ayqvhdtWIVeFuDw0MBq3S9e73hiISxsk26QbBKy+No5P3Y2wH
JebbM3jwWaxisE9R5ggFP1h7Z93pvEqetPitY2VXcp61au5l0il8LOA722ajngdcFhJf/kM65/aF
w4A8gnpXJZZGDU0i2KMyqGqJNYPlyK5DqkH/PZQX9KKW/ClrRHj1sctNezPzbiU/Z6rVSzV/GA01
jfeBlYPG03fjizpsfNwIYDCYk0pnxVd4g5XCyWG9qLPabvZnGaTIiC6PGlCPT9xztwb1x0KTpr9n
jTfHxcK7U0V5cIjav/+xvJARv1DLRpC4jo7o9YYwALc8wl/XTz9XCgYlkl4RQpE5q41JsW5WfP+z
bWMikHF5sIqUhmP2mvpuOsNs1OVxKI+TJR5OA8fIM01/opTlMnlLCKLspL/8CGL+CEPNf0ZjWjHh
+ILVacqQmxr5vdESUfJvdKjaARr0fjIB8wlS8PKoPS1jmitr82E6htq79zuymFL9ezRFwHEV0fPm
MSvRoxZVuPSSDtHJuuB4AJErZGlwJqisBD3mPiYDyIRSEZ8oZ3aatpRMKWayKP6PJkSKs3pjkT61
+sqAhNQ5ywJWZsjMaHfvD6QZn9Bd9pAk3yAUxGK255e7zJ5E9JPfW4tqZsma8/5ZY8s+WFNU7Xr7
MMcM5f1N7Ec2dtppspyn5bYbaHHBawgZ4hCgw+GmKbSWa8TQzNcBPJ70RU0nPY3CQgoSabe0L6z3
AtZ4x2bcokFG7qSvVY+zpza2lCqY99ET63mgsWTPrehdBlctLJ3LfQk58C+PhbowADnckNF5kBeY
vvwmmD5UFt+DCvrP9vqFGONBx0lop7ojttVkWiSGHHec9ZZkPQtEgPfaK+UIzlz+sh/rpJnVcvXj
Ven5s+3dl/ttOsOK0py5CUyn4gcDZ807vRY2UNQmMfZnijFo1Tn63RBIHKZnz4qE+J0l4qJyyHSL
xuME8Cn2faokNcd1/53qJ3LaVREeh24fkRv7BHciUjSEtnb7G8Heo/25c6VEoypIOjifRq8aOYt5
nTzBmiWXFm6XS7d2EAdft89RDmg5fYI2VSxVW2sfxEXqrNplQt6ta3ydDWQJbAhRzCPSgatcsltk
mPyfFXZxWkLzK2bXt/nDzKwLHSOwaC9NHfPlQVIyimTrX11ExJ0Vb5I07ddi0pyEy7rSmKDJOUNd
W+8W4bFhkRCDdUjzzHA3xEghrVoRN065t2v4lCGYYa/moM9Nv5W1GWO09AAqopFAWNBrXJuS//dH
wpyqXip/sr8gtCOkYKEMYZIN3Z76Q9ekDU15jSraoGp/g7lS0LZJ/KTCcIWbB8vIweZUqbIdGisb
Q1POneaXHtLIeyp4yRax0IhSlEWorj8AqwK+ZKIxeUazwUAi54erbnOKdnjJ/4j/lAxLuqmEgx/E
mgza871eKLmBL/bCyWPuIRPrPXXD8sNS7gw96Zs0rjpgxabQ4jSUZ94rL3EQfqDPp7o8NZ2Ziiv7
6yd+MiRDy5rDemJU+gRmGs8hPsNaU1IBMHBXYUJJeGe193dGoXZimSKw65JT8v1YoNbwnWq5xpqO
IjEGpyTy2Pf6nt431O5rwoHpYwsBreDZxc6D2qESltLmmAs7sVdHogyekgu1BOa5EPtX4olky1dq
qNkhml1A4IDAeGs8AIqtaGyW2Dbg+kDPKc0Vb//b1clPv2yFEUnoIAPlR6zyy4POKlkPPQPResOC
tJ9nbMahHihMOz6XT4QAaM+LGdS253vLmwj83TPY4CH+RwZ/9eyAFBKV1xHD6MiIiJfE4fffvegz
MUhz5GF75ky91nKUJ7fesHYDiLQ2giFKGcBSr7Rtag11LdjformNcrFHQrQPaFKauT/NtFkE8Fj0
1iPku02yoT2nGfwPH9mREXcTt5BFD7tFeYS3tZ5DXywcMZ5SULkZWsGrKCek5CAalh8ESOCXykuZ
KnjX++r64A7p6q+PZIaCOOMhUKKPcbhw7cApg0sSXeH+bssP5ik5QnXcQJQoovz5+7GcGYRSH+sw
Dm9jVRCTfvEz7e9Hf/DjqOfMC5jTtKVWWeh65KH3rIGftReFm3RFeXmjJFzbo+VFjkhkdxuT9kHi
qih64SvbCNhA/JCmmeK6C+NR/SCJdTRFpR7WHeOAVOURt0FKFR7LkBVxGJCYbYuv2HP4Zz3HJwO0
sXsf1aSig/loPQ1X2M57acN29Cck5ed2/IHQzURna7/cMqgV4/6Zvx2Dtz1qVEceDBSx4fNK18Ki
DkuCJPDT54XgUiPmOAav0RNtArziV4mRmZq57Fjn7yKn4j7KDeWRJOjmdfdkZpz6H23fbW6TAo9A
gDJfdp0bO/6APrOiZ2Ero2UbZEQvkXrL3JkzNqYf6LGL2CIbY6zIZJGL8d3iIxD+sIsveQUHuU6S
zqkQ6AfZLyjBQ/GUJaaKIPL/lguKaoCAdcjFcInasyWoatLVUH4rN6HAGkxeAXRId1xd1lmue8lx
nWhBoZn+vYWSWOYocW+9e36osZ6sWZyjW6ARHaaVnNb6KwciCzRkOO2NdiH3/xupAF02ENJVwLtK
LosvWeDu3r5p5/s3jWN6whPXxrmMLd6z7uAYb73yMohHUxNazV05edhAwrVhoom+5Xlnb4YvV2EU
atYEqMroe/VruZ+ZrPotzi+3bJwGhxkTujKWn2EkLqe9H+0s2yN4p1SUVPHcn+guUbMlicBGFLgT
o7WZlbAkn6VRleYC0zx207rEEacanvwUePfDewmKi5s6kUonKUWgtlJHBggb2GYMlwLMVXNFL+z2
LXiOsd6+GXULCC34mM/TgaBjB+IzwELkPsxfjZWmq26epZ7CxQI/5ClAoXV8kYR0H2gRiUP+xtmA
o3V4/gyhwtyw96d1GLdgVtlBw8x84+Lvq7hXH7mlvvivquM0YKEn39IT1cImVgd6kjxOpwaXqtSy
z8q6uOEFXVN5KCQ4BRXSujnGxz3G1EEhqzgwBVcAOHzabNKgjdWB15Z4OuMYYpMCZHNIli0mlmEi
nX8jmu0z62FdqLIy3CU+qEgCiJhfv3AHiofSlvD5DNveQN2N196rTzmuTsUG5Zy1xU9LqZkkCRsj
WgM95gNFBM9a1d782GyIuF/0cjQGWj7ChCoqwcH8EquW1huqp8MvGS4K99jn0ETlfVJkuMrbzk6A
/Tpp1+NPAZ9btDx5z6xapf/v39lx0tTFv6BnhLec21xXHK7j8I4e0p47YSlf48zSTQF5uI5WkHoX
3uVc1u8EJ87EjizlPLqm2RYYgWKT1KpKkkgHq3DxNIung9HQJ44KUIKhdQCNmJgSxXdD91E1vdMf
V0QWNCVe1q75ttmUY0sPowfZiaZiJA6ez9Sb9OwbQID3so00L5aHVbPfpY3bW+UOjRBEGowWTr65
1RXS/WmtV4WiPN1TE96ZoWd4IGxwOw6aB1+23Sk7Yavj8pKYnWbbcorrnQLF8Zgxlp67RMLyJa3F
FAJYbekKcFjpIqBmZ98Il2+jHWhR6eNV/LIGbxKK3/njS7YGM76U0Z8j9MrAktcbtxRUG4r8uqbu
SaHpBIUY15qLTzaLgVjDF3YdqeyPsIHrhDI4ZDK7eG3HYc/lwkAM93uN4iItuCWEeBtsRwoWnzuE
yW4JPbb+ws2sYv1bJwav7oAXyjWWBl4a5fKVU3SZzTkyoZzBu7/hHBe9ha4djTf7XmVAFJRZQRGr
nJR/fRPzdP3hBpUY39iyEvX/1KZ/aJyvT9tmLErDbPk9Tk2mjDVnq7S1cfWuqq2MtV0Dc5ZKO8Wn
W8ty1iqt+x/XqFUsCfniE+eAoy56Jkld73BLbZv/sfJOMV0Ky2UKvvF94HBwWbGKU9Tk5hoVuoc0
Dl5xmtXN2knWcugHjeON8nLvDkkfn92OuVBkhh2nHs720Coi2rExAQdctbrRgAkF+YDlWxVJeVQp
/fLDfS9YH7rq+FQUsSDd5lpccPeLupD4rx7hxbdYBbCKRnfUu3lrM7BCgpJePZCHi7nvnmZ/KhVD
e3TnrAJigTp2+VfLdHzn2RB33Z5U6lYkKNo6wbZQb4MmcREf+PIJeztcOndhaQ8rBBTDbPUZHg8q
CCaQQowdIvR6w2p/dzmFyiBVj/ZeU8kEFGzEaGE3WgdKPQUWw5dvlJ2B4RiX1tea/Rb++WnLOM4P
cUOzRKN+lQIdedwyzstKvmL1kJZWD+Hjy4TtR+cyYmHJJy+I6Au243QLmdfQtWufT3pAAkf3lzX7
zBBlmtqnbfMn3RW3LYFfyrnxOc7jaqLP+RcU1igyHRTXeEMxBGeTj7+mfVX+G/LqF0yVRnBxIwOo
aYvmwBJ3xPiv7Lw8TbeUPuJtJSPLerifw47X2xfvrH0Y2fDfDrBR6V73YRwnexuzQ2otN3cPjoul
2WkMTofHDaRQZvrAkUBWKZK77sThVVxkqc7zs79gChZylKjkYvvCsu+A/ijMLT9/POXkZhxnVcY9
L1UALImbKUxCR/Q8CzCXC5s8z/rxXKH6MCsqKO/hUw+yZTXiHOm4H9fCQcQGx4yrq5lwpiicsVs9
BKlfDSfkn8ihtgwRdT/YdsmLWN7TSt98lB7m3ZyKmVbOl/2x8NewQ9p4AHhv5XUS8I0JoK0xUkCz
r+vt0RX+VxQ8g0xM5pdew+FdgGcHMszUSHwgKsdd09HbHdEcjMME1zPhP9Oyy+JcUM3QmKpN/5a+
sJ815rTi5hcMfWX8WOgZ0xKHNgl/03YBtawCnQcZZ8SXDFZhwP8yb0JP5WZpcQ7zVwRfcK6a0qeD
bXfnCl6r6zqljfUrqUcw23gSn21LAazk8AnJJFFcvKmFBZv6ZpA2oOVj5Z38VOIs4Ct3oHWLOwHh
khhjqVq2Ex5zK0VX8sF20utqqTBao9ve+OS2J5kCTDoTrSBH7a6kVmCkUqw/WEGF44VW3yPivDdK
6dV2z2UuhimUGOPdSl6OeuHsSwqWgTg6KpCmE0yIBeJyM2RCLmm0971uvzUtQ9KgOVn8SGh5MoP/
CCM9H2h40T5T1EL/mSG8yDjMxz8XCGSZOjk6CmKIoeJKTk069O70tCjnR6F1vPkDINxeHIaq3Amo
9hHbha9u/wb+ae3qN37ziQsumNuTO1rUdQ7BXKi6H1DcAAacFALr9k1JFodmWTQbm0OWa0vJkXO/
XHjAUIrSQXl6RQFQOSCdLG2m6R0HAnmQseRMQ+k2W8H4530NmX1CruBwLHmtNR1QJhdlVpZsPKkO
fQ/1pBjR237k3mzwwYgyqR/D7zHsiuBnMAx/dOj/YPYlK5gDTBkgPuWbe1F41BM+y7mlIjqXWne6
dpiPQaWtg9T33b3cdaExY/PogcFziUExaHOLmV+XUJaKZpxg4sudNx0jydRVHGa3f+p5kvsSVMPN
n+2wG4T4QSyDcV3dUQt1CWzEizTPdHcJyttJIq+h9PppkSFwFy+2MoyGPA5Ulb8RanEpFfANsKhM
TMC+uho72HDCrHKLkapEevxz8iU36kcIqe8iI9wofWsQ/yv1TM2QSMiamURJMIXBHlpNKMRfcNq2
wSgPqTn0pEbzKRagF01XjmVMaemgQn3la+UFqMXgXwMR0erJ+2NwpKVUJJ78/PXDtkUTVs6k4Q14
FUfKyIVA/q76RGzo2bA3LkrI9o+o0YYaNUzRcQ0IMBG23jKzMMrFmrrPpEECrYC0ZRe0lZbcGiz7
sf+D4ToJuDprejwF+Y1ZFmC0yZ3w7vpJhRcNP/ySkUA96WZxLzrQnEY49CEj9/7w6axTYgcTUqPs
UGi/mekBTxgOlJJtxpXu4aM4dLgp6XgRmuFG68WTKfAaXAzg3w5S/zUAn13rifWl84xvWbM+FeY6
nTyjlqsuvhi4i4mXWDJxbKGpjZ91zOqm5GT9XiFHduwEEciYp2MN45gSRdDT0ZZC5cFB1+pmoOrU
WEeS7hjDN2EOM2q/d5Ikxg0i621DPwP2AgVtdQkTnxcEV0o3m0nDY/sb/Xkw0h847CBgfgh/fVN8
UoYN4g1pqKsImznSBIV5HMLHwX0cQKUjOeighZ2XG6RLnNQhXpJexyKQHS99cvMGtmQRvrto6r9S
+0OOZxHN2RbTHSm/HNOoe2iXO4j85O7imOpJZWBuQMswyTIAc1rMrYJhPFej7INaXaGyi0Jbnj7B
kT1cfb/5g9IXhigmLSdyhT8dKKS1MIUx+aSSd6z+pj9mxO+POeKMdmgoB4xSxF0Zm4Am0nIfNVUJ
lkxQzipSA32+sEC7GEQ35DOOlPyp9NvRFPzeEtrqzvNWPEDojD6fXTBK+aEiZ/GafPDRVbJ0TMIH
MWSNgfqw/NHEGTFsdRWHm2KUauxEDSjG32mC9rp+q5vErgiLteAAkqyOU0SOK0ZrxwU4lDSDJk0A
xOwpdC8G73zU2bZzR0BNcAOQ7g5ZfVoq/XE0ctS0FJfNik1gnWJrf9y4b5/YTPp97fCxoKwSbyBV
t48ITODbsPl2lJLxmVjPl1AxNVSV/SHRbNlPxuPF3Nx/3rCIMsa1/gIWvBrprB98V++NEahPk3sb
EqGxbjx614Ym7yerPUil0fkOW2CtUVktHuZdHxvJoQmyjT6pHrMZ0d66Zvt8KCakCklfBqZz3syl
QqR4xrEeL1VCE0ra/gTx58oKA63mN9biXmH5tcJ10Jbw2hJK8P7/jDj2PXMjiVlf4wSDNdMPi6rm
lWjz9R6jO3p9EWwAbRQcEqJYU7Yxrf4HxZ5moFg5Do1cjas1R3wIZ5wEwuINdOMDIpCC+0oojvKl
n/BbGd+Kkp1VK8A8cvloz5ulx48adf4XuAmHaaMqW+Ex1ktfzGP+rtgow/QKOzczKC+0OdLBC/MF
ScmfwC1MhY4O+ipP5b4O6PSPPhXfmR4/bKU4QmS4vBas1w92AOI5xfz2yS4UWeapaNNaZ/l+qtCB
a9E1dzQIPJ6Lx1NQPBBrgt3EZqcc/S4lViuClAwLg07oQmljxXpNk7Nnb5S5lMEONx3w0qAhhVx4
dlwqZSS1Ve6KLtNfPK7ZuKZIDaZmNLeQFx5TnGrQwTsU0BCIdzYOcF9errO8ja8hAtkdCh0GLAPk
/DQRbAlEanxc28nMYk2LSPlDwsDaqpBLglhpNnyCd/e56ZFdbX7ACTIkkMkrEfjPRHW9dMzZE9m3
0jsJjnxvP8tYEui6/J5UbsrmCOvWfx9RKxnfy8pRhy1eknq1zDAEMMErHCEO3UTnNijSrQdo8UEk
gpVMFTAHxt7EihvarF02RoF3k7pl+QZMs45mCHa9EuzlDQAHyakncjEBlEyDcRfKj1FUAu+arOgv
5BosYAj7r9QlvhNJpINiEtIRMHu27Vs6awg1ShHZEIsryzFjqC9opQJspbk0bnZnu3sCLh2yuta1
IJtcxFq4Zj5czigNPQv++cGRGnhZNxB47lZhT+AbAMXH4LjIAcjxpaSJB4ani7xgmt2rKBrOFDXQ
V9OLyd4CM3BNCOnboBD5V4AGMGJ35K+QBoic6NcPE0UyCLhfzm7MMFEOm7f4YvfxdHVIeheCREQ3
8RWrSDeuYuO9qjiBU3blswIjtVS4L9zNB7UZSefRzlqS+mBAdYwBmpz2wJMzMpD6CFQD47g3E+Ks
iUe8GxL9ZVJLe1vCpJYcS20XF/pxWyehn59teB9GSXRZbhxQ+Eo7BoTAFQuZwX5wuMiceByGuaoj
eLPfSQqJ/je12qj1fwIOsHtmQwaR2pwl+41Xd4Pg4jrXEyKGknWmf8Ub24hId0O0eJnnMu3Ex0Ji
fbeT8Yv86D2A3a5j9aa5PfqaQBEePqtf576Szy0V4FO11q5MwEAJhSMUCsy+eHIcxEdcUz3Ie7J2
L+u/Bw3AScg+5Nq6A15HBAj1ED8ecgnGUokAgPuiSb9xkwwCUYt90HBQMGh0UoL/4+zmxX4Z9vi6
t8tV6IAHrx3ksiTJOA44yr65lLD7GtYXy24GQ6ILk8XRp6yb7IxeTtjt8sIJsEf2vb18SZh/UVNE
xUQMO+v6iY8tjlojDd9mVhr75qu+p8VO7FR6fXt4RcQraN6w+XFJOnuecDeWfTrIeJOJ4vEMgP9F
xN4pnwIZGQJLIOr9hiKp72UTAsGSc4IbJUgYYIhIm3/K0yIPRQhHyVGsiMBDBQjHvg11B/bfz+4R
mNB4vI2JpYEWGoDs5X5BfTLQ51RgmIDojiYb9SAvMGBf7rdekBCyYTuLjf4qOGrHMNFo6egLPVF9
d6N/8ZR6c9wJnqalbU4WYZqqpw4gALl3Kt29ikb+4ETY5DjPaJjQAitOGOD7wJjp6FzjUzaEVx46
g4/ZF6/cIky1/rnCLA/TGchreSMazVZVe6y5Ph6c6c/Mx7yZYa1exXIr2yXEDTCwU6XdGRd+PdOU
KiWZNHDb+OCQ1IZBX64dAfjpekndQll8EivW5GilJBpu7aiCTjPZskghlHm1VYqCxzgoSrp/72OA
XH7eC0u9pWFNRt3NGD2FrCnsshifbDCKwxfW0GVuqxmRx2vaAehv2jMeJ4r3GlZi1FMKgQ79H2l/
tCmJs6DgCbkskV8sVJqZRf6nX6IKPpMaAAIoNPxbfrUPByLmVBecXrmT6UMeU3ysnfqw9wJaqkjf
09WQyES+u5RTp4evKCZd7fXojD8YjoSz5+kOPKUFpMI4V6jsoY6yvg9a9pYIJE4+CA0KO+NAMxEk
eNUI4sKEAv/MwEU2wjtnkpLIW3GMXiTBK7r5rLS1AvVskBQdCZ7zvEXZw6pwtuu/NG81gXMR6coI
C/Vi5RHg4PyYCcgoU5jAFx02gyAsYo9pNBVlnw7hmJmX1ygX6pbTI+j9KqaLjeqReTVn7A1YHtK4
JeO738VbRIZgBY6XyPy2qkkdMfQjnXLTgzvf+rVW5XmKMPI/4UBvL7dc9DbzcMbsc9qIGvC6JnyV
F1yFX4rk53H0YHPEGcPnjiw0u+V8O7axPozrvbNPmvtjiI49INGSmeoewep74UKa+vxFoW2DlsjU
aBNgb7SQTPjLNYJmcZnK7Wc34JTwI6+DCop1xeGx839/8nvjBr4DV229rNtBO8QdEHiKml3ExILZ
S8JyIplCc9PASzq+Zd/iAs+atlHAEQpCciclru/oVzgS3Qa7lsF0T5fka/SGd4PzYqqDwQfb2Sg4
4X5SRuHWFfgngAuNKWmkj0avbvVytPz4HK+XOjyKyGbYZtGjIBdG//X0ZWgSzVtFIzkC6A2lLImQ
98WYzFgTS6bF5mAfP0C0ixWKna0w58TaasfRiIo8WA9dvPNtgFpQ2E4ztPYiSrTnb+Jmjy33L8wH
ZRwvDrmF4nCp1bpJQKOQd28nF0x7FaHOTESEGmMkR7YDaW23I3mc0H9khT5bXHyvUNlfOhuljlV/
0KAuIEchcXEGgF9+HwUgjqNh/Mn7Yj1pnRHFUPARouiE9SJ101GV75QaGgJIgmYu8467i2HYCR9O
u4cvoFFE40+KrIbFrm+6C3PsuOK+SNwLYhhOB5GK82RXo+iZX+7oAUPZs8L7Kr9pK2u341tUc+42
2J+UqwA0B+qZzP6toqqZ9O3aGzKJ57UoK83+64tm67lDRcKrjT4L9SlSAC9Kj3FHFXkj7lMaceF9
PCKS8bll8gie2y+p6n8InWzoIK1404NyY4FcgipppbYp9vKNSM66TbTdfJPu+fajdmnY2fOIg9VI
2pIhTKwbrVhTCMf/6RE8l8WPhUpcC0JXsyHt9t7euU6W2N0uW3H9cYXfMEQ/7lhtlRUZRPqzQvmV
RbZOMl0CPSt9VqTGIBZ9ouIA//EKzyFuwo5t4ex0wAY085ZvJWMfN8cZTxCHpdH6VSPybZSW1VDZ
9cICjjzAfwU5IoU0Ztv/0CxnjLDlKZ1FyByvdyd1jLPc7DHn3hW1b2okGOi/9bKEAmy2WXQ52Ru6
pMLOq70UlbBqA3ulXXgotm5xJQkGPfPXGkIrRXjnwg95wW8eGr2UJZN2lJlwygtcxpJ8HoYcB7Ow
6T4GiGEO9xdq8m8xXguSqXAWL93bUzP0naD5N5YdC50JN6eVgqwgDLO+6nvjVCLpLxIgyZgluYb2
2RosOOqy7rlPI26mP+JplT/QE23Nxkpv1z0ZW3PyDupFv36xF65iFjrAx+PPBXJLSBdSrhgBnvTG
OpDveD85He7oo3PKPJJkotWk4AuEU4REZZyz48sClyjJ4/B18nQDszT8Kr4onZTXDUPTTjZM3mot
ATtn3zmTP6PiO40jSyXO6G6ZyEfteBCTmvH2pvTmxwypM2u7y+0Tul4ul8QCf2E22NT9IoxrUQxj
B2lJQSNvh/G/k+l+u0HWsJzP4oyqbUhbfVnhSz2TY6YXOUMUqTlKuCiS1vIk1EUQDI0/SIYCsz+f
Gq3lhBVvLtN0VSv3d4IABUYlD9dkWRX6sTBmt3o75r7JI0ebyr1dRxHoQBTT+ut0E+y6Xt1G4ZnC
qjk7mgceOcvhYQhixrUwYFgISntc1uacCkM/ABLK3CV01J4BXzx87EqxVkFVNKWRyStWPv8j32hX
QBMT0WRIOQGC9dG1Pq2Bh/jPRCkRSI6coxH3P5Js5HS0PHnGQ3ORpiuJUf64dMB+e/bptrgPnF2y
tP/pg9/7v5rqsyvn/C2F//E1oc+HLqvTbgj73ZxVJscyQfX/zGgIsEE4uquN0Hx7u2GLHdcypm2O
38ywGOkYc1Oaqjh5XSxdVqF0/mYy4hbhBRACycORA4r9dJQD0OwrGSkegwXzyK0jBbsFFaCrvP7H
zSN8/jqt05FY0qAm3mkf195unyceJZIAAwUdR7oB4fOpgwbGCqrlDn9znVq5uZJdYWn0l7XdmwSm
lQzv7Aj3rWFXNJnfXN76jW3AQBmZ+RqzrUt34AUMIYMGO4emJsVfGljoHt8m9f0Es84ogsDpsnX5
ILh0ARkGz0/VisdUNK2J9gzZdEtQsaOS/uY8fhlf6xkFXTNCSs1hKiHGQJntivzkzeTCaxFkTJqw
jbRMAnyWGD29O/Q3vgOFIudpLw8OOVMQ3h4rLSR3ptaaUdTBklSgfDgqNa9CkRIoWMobHU75CzHl
ramdUjhb8O2Fi1qDoiYd0qA/vqZiazveVMqY9eY74v4uycgXXyxdfekxNfOr6ziXwIiSkLLSjn40
/ULkNFLmnw9Sv5Qw/1AZ+E3TyQxyHoGy5RmP9KzWg3rbFpVxkfc+8bXhhpAnKJJ/kDfHv4cgDH8Y
k/kPId5ayH7xjaoVzM7tYDhyZRUlpZxB5kplLlBbCCBhDngIpaO+24j8kLLD+olREdvcI/SoHiOI
lz+2JUzagtvGcAKGNJrHbJbunG8i2CDm58cs9sPd1zQogMZYBDeO3Gra69Sql0tvdEM91KPN5cdh
/p0kL1TTc3qld5Y43/MOkKW2xKZyTDuf1DPFaZ+7fkIIK2N5ox3PwQ8+FUxO2wBXncN9ZIt0h3J2
Vu+8tEybuUw02GiUhDLmQoF4TLg34Lq52HsAE1HIseBkypHja2TiBUYmVI9+wSWk4AZVRz2A5WWT
4oieoqwUVRyawW6FZGqo3oELZTJg9nov0IFFD6Jf1EyKKgQwWxtgiqstFh3pgORN9DKNf+ztUeqN
sBQPZud95ipf0mVZKmhYAXRo+UELJsigj4SIp/32rf2+oPtyxB+XSk0gdJIBqKiDT6l/0HE2p7Lj
aremhKrGJQ+jrO4ZUnsRa7kL4STzqTcSlE0HZrEE6czPRmzT9gsHpCXBt/X9PKcxt09GuyTgvqMK
5ShGP43ve5jUo7XKtupMtU0O3+0SDuriK/P+nCj3WejaD6CfnKTARLhbuVGU2PdHAvxWFOodwpvJ
7BGGdIhUktpzljftnTvr3ZwidkRx85ZkPkD4CjJnXrUJ/x9GMOPVQM0UuoTWbKm7iHwPTkoWs9V8
JKzUUnoc7/ChMUWIrdpPSB55oA5iNjtuoeFKCnvplVyPbB4ExHQqJSuvtOh3GXbNWv9ITZH3IfUo
I55uyHdV0pYB4owjFFE0IUaJVR2Sh1eoU5OkSn3OZEim5zH0ESxUOE5GmGhKaDALV4vnCf7nhZWw
S5oeKnzbbbX3bHnlQ2r7w8BBRRrWOcNES/U6t/OTvUF2PDNDTGGYPTCHLQohg/lTN0dRQ5Plwjiy
niFKUQLaQsc8OtOTRhrevJ1XViq5PsPdVlHqTmy+cbHimPHbk7kRNXH/3WUVf+apxv0eqzNa+ius
MuKN7aoDs2D5YaQtyNR0wYeE5tEUW8TbloziGM5yQy9/mSXP7ra4z1zaUCe4YU9cLEVGQ4U0g4YF
JYuLKx3HCJN2BFkkR8LlmDPxqEzL/jKbd+Oq0PXs++zrd/W4lwYXJn6mBboQNj6xPTpW6WjqEbg5
PqmY10r4UVwaS2zPtoxRLbRgGbA1jAKiQ0gEtsTI3cH1xQ/35CSixHSRXxli4xUx0H1WaZQ4/YGp
n0C/y6RTWLzX4qt+hZlWj4kfkiNnw/atxlxmQjMjDdT5FUFSmYcq/lP9JaOrhIZwxTMP5r3/UQZY
GKeitvhHerLG+BeTVmPuCQEI6PavMJHgmf7TKCl1mHyJz/gkRSA33K/0HQwJq9ZY091+jfU1Xvo0
c3Kl+6H0ngFIGQHFwYrE/batHHxKT0vHufuvgaGv1DskqxjRH51gkky0pDShefdSXt4EBOIUbM+9
x9zrefBH9u0Af4r9rS72G+g3mNkPZGUPdjOkvJaHRnKiKlTObsK0jpGe/CbK6zhd2X+vAs6iotYv
xXk8f0JGrzLN0d7xyX/DUX19FSSkb7U1cztUOHvqFzpBXod5osZL2Y/adkZpD5TzgSgX7FfaLTEn
MmcgchRMS1dTEASqXcC2H3a9QBTCYUImSW3Rv/B0cTnsMSrElsFEu++zNJbTJGZJr3FkcjqjoAAo
mPiPGsZx5z/qwIYaqUgvNAfwDWOd2F2AilqacMahrK3qSai+AV9r0jooz9RrP8yD8IN+NgtUB/di
Jdb9zUzjvOq5e5otvIig2mHm/4It31I0+qgg/xOcoAM0nqkez6RDk3A3DbQ3jLc9W5IBugr+Cykr
+xQxRcxy2K6OXra/ycuE5sTHTZxHYXGk0yU22XS1z5BHppcQyFq4XOLfiNMqHoWwwHHSLtSpNmnb
r2xd4vxfCY/y/LkMfV2a5mf+FMNX70fT/N+fERvJJE89bOSVADnRB+YR0VjepyB4v6LJSfn/3y4H
kXXTM+YTzZ3wL6JMOlvzrrhn6UaBdmXVWLTjc9bIkeQIi/a/9I+8/QIExxKmSwFrCh/S/bw7QLSX
PGzGGgmM1KNTpcso5w6w+V6ukMpgWjDiycsjc86/zmpA/jpBPw+M3QHiYTUUZPoPUMfirDeoQl9I
75C4JxOE4rTHePs3Z36xB838TrVCGVxgGYs7IMwxZLcee8x7caJnBV2KY7dzEEzNgGjyyfnd6HZs
jQqyTKpOAA5aL+OM8vLH2hbeEZ5rBxOkVbXt9yrIyxVxZpGn5kK9cv+bpyz/lQweFmAha4iJJ1to
aKIjw/Fsn5UBXq15fur6bl3ELLzrfR53R4ltbMQ6/eaeRgrzHkZieFZEhtQq0ZGTGY9ILI3/6Zjj
uDXKEdBtJUwQiJ2EDzKpCj7GbaL8JuFGg9i/bOfxyzS/GYaP3oCHW7q+cCYvAclSUmEdMzjACkEJ
qSs+ejmn+qor683pK8Mr7j9WVjTTrbipAcXqA9IQvmOrkmBQME8DZ32FS3TbMyaYfWHrJEbo6zlG
JHn+V74uzcV67RV9/DSW7xlZd89JLF73+dLeZhFsQ7mnmpvwLusKH0WTf3kUf5hF19M1yUXi8aLv
EWsUmsOOYX47k1ggmN6j8XqGUc73JJeJq0qB1Z7TC4Rmo83rhYidpHU38ipVh8bjLkr82dNCUfVJ
LY72BlAILPLrJA2ZIzGlhtw+5i93dOteHIu6hXlub8FUz82mCNlXMmLDBR7FGqfZls+s15UqFUfC
PkguCaQ9co2CI5gPmKJz9GXWwVsJqLR0lTaYq4eg5hC3UeNHmGETB0SAwPMtaTTUc87wmmu/8W98
HSMPnsvXXQmSp2phXQ4JiKz32rL565jbbLe4XTtRefm71b8DcY9lPQl4183h+kwlCEuqMlMohJZx
BhuwQZbu/nq4+8L/UOQ4yKJBO4xIiL7x8a/Pu/ozlsGW5lYzEFv6NaASygF3OEuzMCv6ec+t+g+V
jkCPsXCaLWqgT4FssPuRNpFa+B972CnZAspbEYVyhv9rzCRMGG4T2CnZ7DtZstR562UwJYWg2hxY
c9ytF+TLueeBpXgzU9OoK9r6XC+d/wFd2rRddQKG+u1O2IkTDPrYQDzRdlirm1pAfILqM+L6Bcac
IOMwpJe+EcV7rL5qNrQC/YfXSe02l+PHnWT9oreB9p8NJ6b0kDRUfCwi8EGhfR5L4Zd/enLWQDCI
Ng32dbx23WBAWnZEApGozHoRGad4BIqRALBLDwGafDjX0faM6koQQwPzusvD/hko10nWMFMoih8l
A06cWz03ioUF/Lkyw9BpSEfsH4JAkG5AEOK3GaWThE3ev3Vm+yF8uZIrlm0+bx3YEl5wron0M9jd
HA7pjw48znMwZSKbiEyl/XkA8FUZv4gknHHvT2WmqbnfFrIJvM1NAvADUqmoPzwMsdzP2bXPUNGM
4gjY7tYZjnpyg5k7te1ABHykBgpqipeYBNr9iccmHlAe88caLtumTLAT/yYCVAUpS5uQTDY6jIj4
R4cC/SQ6ZLEBS3qsPF867kl8JtApj2gW5KzbVSOak2EwFeY7ZgYPfp4FUqMJiGlp8eAsKRrYPRoj
33BykCUYxBYQM1VGdgqgAVuVNstyOWV/BeKWxE/r9RZPvmBpXgkShEY8qXqBfDiS3kayBwJT9Q6i
bzs9IjL5J5/D5Fm9+gAvg+fVuoCQTBq1e4T5UNMYeqeqeTAhWHcQ2oUs3MV9G/lPx/sz3K7UNSzO
aMSRgwN3SVU8RY1SZC3Do89nap6Ul5xAIHI8475VJRyLpfARkxGj9OY0Q1Vrpv9yBk8AUeQmlhXv
gOOEdHsaGxPaI1OpoV7bTS+ZgJuXiAq9pWNh+UuDEgo/5CQB2BUhi6hGcN4962kFu4ikc4z8m3lU
zhwmODHsFBCkUbqmJc6MqL29VNV2cS++WJT/8ZA43TXXHXzkFsEWmNjkmem4ir3RX+ikSO2+MeEB
kpZIr/3LoGzR3uZG9yjQJmsJ0Tf8AGz+2mrY5q/EwLzN5o2cu7hUOMnlu9GCCcbhvpn9tHijITni
YBo1YBf8GEAJ9XXH1ccBXCr4IumMST0S3JCTKvwgPEJZeXKyh3AHJL3gH+bN+XkwfEPIXK+K3tG1
YcBGVQTeK3KrNP3opUss1HhQiaoP6uChSvk81rBHx/8Q38Y2FqP5QC7J10mErLf23UUz3+RiHVIZ
SgZ5neGewCVXqexMMrq4MnHyJchMVymtYu2rxx97mAA97Anu7cSKwKbG86qSPiZXa5dZ4xJVB9vt
HBrP3T/P6IukYwAZr50AWDsZHOsjeQ5Zt8LHPHVuWIM1CtXYCHHYXZqK3tdLL6z6f0u8TTiRWw7y
ivxVtEqsLE/DM5FmPk/jR1B+CHjMZEbIxTUHauJ8fEZHy7g0Eiax7Df32hEP1mhGY9lYFyysI/vf
yEWLW/cjlvg0M1Xqnfq2X4gas6qnuZC3NhpvmqHLD6cwmLmjXucceVESKpskI8KmgYyZH+TkTyb4
FhLejtLe3ywyv8K12RA4l/8/KgWW61P4/j1mnQHSPkPhhKFFsXGde/NTLgbk/xdjPXxcwZ4ELKT9
BblDnNv5QEMVkq3yrvmYzIjI7Dxzl/5LNwvfuIeEgZ4si6wZjVXL8wlcu+4oxZCgKuv/ONlz7rtQ
uixesVASbZdrV8xOyM3Nx2QMCRVBZF0BrRX+SEMYTMl1Bp00oMGDGyxGP0t9PhNFt5+fAUemfoaO
I/k+VJXPCaSJfIj8uJJ5LyXC0yX+VpUuT4674poFzZ8oxNBt04/Be7x8bSDHED9OTQF85HLbPTOw
2d1CEc9o8UZ2BxirVUnMvi731mf/6pFhtCJIyr9J3j4+Gym2x/i1ozYCPEPjM6T70CpsAkQdo5qk
/SAmjbuOoZKKUdQruf9ordU5zTa88w3QXK++Mu4Ru5+N3anQON5j3supY4c9f3k8SduzqNhUmvyb
kW0Hlvp3ko338Qc7uyrQNZ9jOyvRW+uxhOJQU/+kGooKyHbW6OysojzAIBJfShCziApIF/QcpkYI
x0KavE0h//k/h8LU7bELcyyjVs4d64PU6AIWKmtPPTgWoKg9VG9+MXcHJSoynO+B0p7B4/Ogxjyl
JiczJVRBFta906131+YeM4TxHGMOqrh0pvSwnzhLmptaLXIaM7qr9MJvLYRZSpHKz9MZ+vhUX453
84Op3gowgt3cAJhu/gc5GfpWaOyuptwN42mo8NS6trNA62z4teLYfMBa2y1cPELotjJ572Gt9v7+
A+f5ifSFS4t6LF5zsPk9YAWb40Ul32np+QiqEkdtqGlYY9n+0nqHmwxqg2G5WYggInpTuZCbw6pt
6Bd2RBxFPrWS7ts2eplhTTb2OlzhUrHERAJDsA2mekYMXtPozIkf49nX9+Nlb1A2SFgEjsBriFo9
CyRZ60plrMupGnVmDHVCDNDdIDAgBbVEHJbbYQV8yy5wCRZATSGTw//zjj9qq/3wK/lvSXNJYr1N
7RHj+Gkd9m8E2gHlVPd46l0LkOmijigKTY2E5kplKtxBq884luwMlXOW+RnE5vtM0N0ThNlxeNQx
dv45u7VzalrwnMNL4pgN5dm4lsg9EcgZ9GU4ElAXBnzKnhFToeLHZ0R78sJTg8CZrfkTXxjOC0tq
xz/fOKowk52OdCK2MOG1jZsRDA3kJAn0PRpFmfB3aKrQ3MWZwTE44ftRnupKRkPS91N4Vv7p9EkT
RQ2tWo8Tr1jJsaXxnk+IVueuuPjc78gELsygm2Lyp2H4lG1pguF1o9p9/g8g20rsSv7Zp+NVBq1f
jyZ4IJ606YVLfXOefB3FAtinaFc63r8fdwG8IOIu54y5y0jerdhS0soWMwt4lUZC7tmNIR+elXPR
+y7ggq7UZwudd017k+Wbwi4Ybz9LqJkY7cXkU9AU33iioSwaimaWpuiDQXV8vd6GpZ6MvCiJ3SMJ
JRsD/oqHlW3XQaCZLrRjI6G1h+yDkQ0SRGvUBXZFppb1oy5h/bsqUdqf10XB//pmfoddxlEqTWgy
LbfZU5oCzlKtrVahF8CVpe5bZrdwstH6Dv16Q/b1NWJ18DjC/tGoHaAOFDkuX/8qRsQBwkJKBO7s
3e9RFaN2tXyoe0DfDDwKLWCJTw4zIc7QlbpN3tXVm29ephntwiyY3D5ce3MivIARYHLYIgCTNDSN
fC5eBZeEK/LCRboJSEN8Que5xGWFfccu+/TsD0WV7tcQuLEdhpuQ6kotVfB75UZ2Y8MfV5cZj0lu
MJfysnAqZqDxHs8/yj15w5NY7am+B84GBbY9hI+0fz4oVw8x7ozxnkfGAvpD5bROgjO8ZMkvPbFT
m3kIlrw8JJwunQ6BbWIdYU04rxNNBCiut3kJSerx+EtWMmUE4vZN79gVfO35QJ1VWYbhea3UxgXV
Ex9i3kgQz4eHYgiC26Vhvxn+dk4VBVwPPI+TaETH8oRJM7uWQKOC2bZfWj6ZWrmL3F9WQ26LFZLa
OK5cGrwJCnG+qcynCwEAvziTf6ObE/J0aByJfgXS/lgr0TGodLjCjzJS9TjGtNL03Ly9c9k6D0rF
jYtgTUEbIlcn4eaojBxcA14AbqdKOVBP2Olu7LwhHYXKVGv98wWOdxObZ2ngwERLytcC9LdvVAd6
6rx80cNAAuxKIVmhMHPjumLtXXNPD3fDnB8DvvQ5iLCG+7Fkiz+totCXFWskqWd9XGjLqI/7g+Br
52CPJJw6fjFYlr+V/VYLen2BOQ0NgqOIm3p+ZmlHhjGmnWfom3pHF2vetE1N7NPZ8knq+uVe550E
OIdcNposAEoeMK8McbpuUJ+o70jlHvYDdwgbZ3Y3S52yYF4d/KtIEa4gGkk4B2eJtaavPDVtINK8
aIBK73A1eN4cmj7t3o0GsuRg6nunQSkmHG8Eb83l9SQjF2eJq88QsLpeAbJCDG4fKk/yJkFTsY1C
ArPHFrT6dznXR4AF0ZdmD2l5BMQd+TF8GL3OICkBcGO8+AbmvCovfyING+ALHXCZ5CAohmYuRAri
rWcgyoH7m42tr84Gwqb9zWKI0AiXyVzstMJRyQzaTkEeO4uF1YdPrrzf41JXl/1nB0xmjOP3UppH
g8ADRZHiwOIpdCobv1SGFl6g4hysrR9QmvplK3oN45RDF/TgpvP5/TiGIZ7jASArzKxplXdDWBm+
I3kF859DC2PNmB/W8waqDsz7SUeMTEoDWGUg4GtIPxaDJ/rycU80pSa/7HHOykYodgVZCT5xrphQ
t0ZXeLr4wRUKNSP2TiIvH80oqDkwvItITkHT7h4D6FrOzm3TVqthFpfH4+ltft5TWyg5iumD6+68
0sDva4PhGoEHbmArjUf3nmCROIBLWYcUQgtwVnX+34xs1xU+tBcsNqkMR+/iWwBgm5JRDno4Au4n
vU3TesUIaX/jInGYsDZD8v7hzkDOUsmPIqIAb2k6S+1jPuxUFSzcgd6lcxkf4IfAppIq7q36AP/I
i4DUVpqONJUAguKgDZTDpaFhTMYti75+XTPGSZJQkcUkLe66aGrpYkIVhtNPsotJEoUVu7elcvx0
DrAGC1Iw27qfzYqjok8XResEMF2VhozK8L992d2R5oogGWVyUIK8FFMY3IzHYjUl9MYSaZ3JmXaf
1dnnnHwam3hc+ybFXQOyj1y/cJi/HutYMtJP2meNp+s5jx3KgbOmMwLKwJuMBLfhAJJ7kN5BJLOV
3mCxrlNGnuTShIwdk2ebmOUsdldkoaTuSJiTd8mG5uA7LFjVf03XBHRdGr7c4/AtVegdFYT6szuw
94gqH7boQTEUcMeK4k7KMGCFl3XMOcVIdn9IfKtQ7JdQ3ivODAZAdBOq3ay27uh5Gq1kSqHB2cep
gkOkD/7/gI8+Lojn4VxPGlnQu8DEvYsZhY7jpioALoGFbeejNCUHi4zEdVccQUfeEZkjlARIFCNb
CSVvh18Ebjl93jqLEqlHarmREAjJF60RTWi0GEOY//TVVP8A0wLMk/p9XFuOM15eXa0V38WVkrAD
GtybNzmNr8jCt+KnN9XwaaNTljOcA0GfT9EMSR6OB38aNV8KW/a2wEEClr5B4HzYpKcSl4eMAqL2
vR4Ja1WEKddf53XsJxKtMNbCvQWiELc4kqF8ftkv2NztG9KgYAZ18V/fw3AjNRqS7R2EBJvMV6bC
sNVV5980n8rV04j9U8AylJTir9DyU2oSxmIoXpXR2hd0dbAx4OsQ2vXNaDZmENUE/NyKSLF2e1Ba
0I3kAhTuD2iy0GwY0f00Uh7FlCIPBxe6Vo78qTZadtCdQrRgHAlsmKJqwYkuj6jpT3JPAGrtyuzr
PywcFCbXYIKi8VRo4lns/6P4Nn6KRygCZ1fRqRl9W41Wax2oeU1f5TZBjzqDIBsEfLZNB6kQi5Rv
BFQFxr4SdGXMW5dnbloD9+G7sNIiq57D5YRLY9NF40FJY44PwrG2Xs22wWRWCyzjAWGylDxZ7aeI
3mgooTijcDpkY2Xc6T2DiMZWQedy6EsxTL5+nAZ3yNhQR7GC3yqkeRA25W0kma/H/z6j5odXPfwi
eyVdKH+TB/3kjQOkkFDArtgUIovgKXUiElfTSq+QEvk1Ok1VKJ+VOhyO6dmuh9ptyyDcKqGrDWz9
QBHeqcPxpL1Z/nV/bNUlAZTZirW8o8IAMJXU3PudW1rYZo7KFZyHNl39jUZPkLx9HMHu5uOKiRk4
KeR5n1HIZHLZkUAlqLoYgg1+2nocnoZdW5qL4/CUm4fYuZFJkcz3IaX8r+HcYsQbgxVfutp3ZxRt
4Lc4tLY7YhDrADMoxC8JoVpbo94ZBJ/S5+D1iXpq6Cu+h5bZ9gYL8dQLyuE4DK8ITArTwjGiSYMO
nkLWcs0wsVe51svppH1egLks1i02gdxG3sx4tjU8uJJyre6qj/6lncUMCfdevm5HlQZ/5TxXSZXM
d0IoS5uLXgCntNw17cUY4bdbPEJUOK6fqv9JbDkINtrBlOARACEBIE8ohovkrK2A/A5UU5Y109U6
3sIXTm0fGgPCZiNsJaMIgi+F7CH3+w9bV6FMuLR573yByxHf7j1tM+adrle1JL9ihj5yDmT9FSbz
2nednCIvzuEnAuReGu1jMWW/aMSGI8Q1U3LqB5Q3EAQggoGFt1aH/VKEm+xoA3TDHhA7ykVXu6BT
WzHU5Cn13yTsf5jpOD1ljT/X/HD1VDbXU2QYYbPwKu8V24SAaTyrF91RTRSJ235PoJdu6vu+MQ7A
aig43RMPAlN0M6Cga3QdKjKzFcVYlQ9SjmGCNbte5D/1S5y7HZhhM5yMuZsOl20oRuZlY6ZIJ2OW
u60Rv4OfMGTKqDMSygosUr/fm8Jm4066aVK0dbPqlzqcP4ET8E6U6Jlc5TjS5LaI9R37N+iJDFuw
wqaPOXTaLWsKkcdT8/KHwPL5UHSiWyrVGBjo8fAWsaFz5MqwTBqIVf4P0HUs8fbxGV/wP9AjJQGi
XqFYx2Bx0FFJ9ZjIejbxV2gqgf+JUVtQu96m9UKhBOIecoq7/OUdl/gkM8Jb6nVqII2XOFqWwaej
gsvQHDTSLXO/qyIPngF09CyjWbFZsDQyES1e02F8E5/HeikyuzTINtU+DT8Hu4RMiWiFWzf81AwS
f0pIA1W+LPz00EEZbAZ/RcjOwebseWlzCQ7qZo4X1R4e7O01OjWBuHay+4RQmkkQgdVU1NqGnKUt
2c72lBgxMUNc2Rz9wMBvoMrkbWAYKMJ7OKjrn9HaqehoCNaIrKJeuoMi2y5E3PzZ9e8SjQUM4wYL
xcLkGEmZUjr5oXAWkRW0v5IPUq5ebBaFngMSy1uZXiucGSgazdpn8X/W+6O1T2KQJUlGYkpN/gha
aOvHB5/N3vUGsbTmwhRferFybGlfxfiAdZT9mI/fCtnkebz9hd58sZQSZaS+VujvgJRMvZiAldx2
FfVJQvBB2NdOIx36uJiyP5a4wSHocVLmIS5kHovbfeYh2rkhAyzkfen0p+0cpfOXfuJVO+Fh6tED
azSSZ6lgGAA0XdNPLON463TyJAj+xsSP1gV5/9D++VHns2YN6TmBQtN1px15MndE5c4n35dT1n3c
erYa2MZ9Xu8cKjnqEXxMXsJmnTMTNGqs4xS5OmimpgNbNB4Vcq3rBweSlT6n6klk49qU/N/tPhiU
LHoRaTM8VWm7Q7L5pgxRQ4RlYZdIGESuuwGLBoABX3S6+IYUVdoDdkck6A1Ek5WxPMK/kYo8hRaV
3WavMUdDF7ZZdWrSkaw9ZF7GDTa6MGjvHN94KGz3bfmVR8P/7QHelEAfcglsD0Iy1a8Ae2+/o57M
G2HuWMyOW+eOQ2W9bpl9SMVO3KTEHDQ6JaBLfPBAgkYnM/0+SyYL9aAo/lnUf17N6Np+oH12KACY
5+0++K28/s7FFSIappv3DoeWuCLXAxMhAV5piwtRiQu8X0v8qBco3X7xVH6cYTt2BN+6yTUR0Fdt
BqxXoDFVmcKf/YZqoYzxCqdpL+xDxyvKPsptcBMRSaT7E5ZCD3zqMPFEvt/B5O5lafbwPdxCKvHH
fub847F49huIqrbqEvZg+9Fkp7QCFzrT0Cq5fCY1Y2F8ds3rmQ5X0ucXwkz605FyB0VtMQFzMmJl
U1xELfyZ9rnCi5+rBt59IiQIXmD3kdZmWwDKGHqWpfmrJ/l9XmufZFCqhiP7BEBFg6oxB5x3EI7a
/2DWaAM1vhLYS0+CJYwtmvD0DZeUyRL6nImw6LTgkV4MlOSXiNkFudGVjY+YGDKo92X+CzB2c9l9
MV2TB+PGTd7DA3ltC8UISyTlqcOKnxvriyMJtbFPZohBtQpAg6vXa4KQdCKTeQMClWxJXJ2bmym7
qW52CW+YTpxtEcpxSBdeIXSWZzyoBVdJ44kvH4P/BQRWvodr9tbLYoRW6VlirCuLugUeu1EJMJLl
CsQh2NW7UApSFWKdOlFIpVWf5E2A37J5BARbZe/zuwWK32mi8M77X0r6N6FBVjLtbWLbQyw4k7n3
i1QnpMPzatCrRqHgK5ruwH7AYWhdeyvtLWlWdDJW12/GnsvWvJuj5GJgsDo62bL3tnhwajAtraiC
ZEZUEflCXR2lkYwIv9VpKhmkFGM2ATnWg9G5tbkS8fS794K7/lh3u/GEhjjhuMgFz6xmdPvVaqnL
gvrTvNSuNjrTxqvd6W+pPjD6uijpX5P++8Ocs3nXw4mlLypAeU8Fh4XgiQKQ6dPDejo+uv2peAZG
k7fbOwQL3fwIsDW0F/N13ZXk57OlcWe1loWUlUlhnpTGDvvJmcxCVHzouBT4l4yCV98Le5/3eGMk
Yt0aYKpnR0EZZ1PI8jFRXU4GT7UpoSsFeUlSNlBx4RbvLDDDJfnzCqCMYTsDO46aWK2H6dvQnt+s
wiuVkQLklUiY2KCFcA6278RTopZD0APMKNdHTAFrd4Nn2Y+wGpIy/ugO/gyaH6OVEXPHNtoSDlIu
ngf9oVdviljdYNtpmH2MQbDGHLSrjQpyH49yMZ+2FpLUTJOP7oZ2h54xlaA6vew7XD5yKqB5TpJI
9qjM0++1VzjHNPcW8POtGeOf5McEobUFBx7t7O4idsv13s9sFBLpZ18bWTiDaGd0Q1GkL6DhCSeK
dUJc2QRqklTKlyzgrgHlUWHNpzR2P1LWQOzxQJLm9XeWZ+8pUQ0D45Ig0/ZWv7OZjKaGSB3L7eEB
rcKYWSqzGRby/euOTheWqQCARdOHT14tjiA7IVW3oSKCQL+R6BF3QkAn6tYRXAD//t1ZM575Uknk
eBBQGZtrhBnbVRb8CcmEyaZJzcnAlKTx3jZYDtfocsE1h0GKm5S/HkDNqg2Rc+il46lroR4pq1qx
5vp5Az0qLkGcN0g4M3xK9Lhifz2wZjElnc6Ls1sKVUr9y8DDqMb7k/45c6PUToFCd3raj5WXDARj
RkVPHjbf6FRlr8RJxf+SI2kwdc340T5jepRX2GeWYVnxMqeyovxGPB8hfm630LRl5SafbTNPVfge
brEwRfcTadZN02siaaBo1uwuch6wU60/z2f7/JjVimQldWDb59Fli+FwTtRW2sEZH1ldNRu+Dik5
oS6Ey9ve+G07lGgs/ONd48Hgo0pg9wCyaYqK5rYwHwYTD6MVv7tnHEoHp/kQerMEyoS2QCBOTWRu
iO3TnjbDGm+YpzbIB4W9hIuTue3F2/CNqy/mHYy6ooTvmEw9Bh0QF0eaACQC6MdiMZKVQ2NIbhQN
neE19uoi0MqUglQZPbYtkbFXdITFPn3GQkjHmIXlmzQEpm+Z9+PXz5zkru+HyAsZ75hOzdMUmrbO
Tjb1/HjATlh9HsMXBAS7tQ1Qcw4WtQu9zhUOObRhSlAKaySRw2kA9G/fgpKSVd1D/D/5SYEGb2Xi
mVtyYELevVLSpyEiuhTiYKqPdwUG1ZL8sHaSJN93vQ8tNAdmDYEcR+PDJJtUKV35BjLEgvyDwO/+
4JuqvVyt/ZuCVJwZB7RXLqTpaSOczTFF9NJkRA02tEfhxkK6vY8r9tq64gEa2eytzGap0ZiAjyUB
NvzLJAirxRbSw69utasAiKQX6jzB76VwdHkAUsSQMdGd9uwQqa5wa3Ud7bgsrEDcnoGlvg9qSlih
wD2pNaGnMZo8wxETiB53P0/ULtxluXoR2VbAh6fkVCwm3Z+61R06hR5sHOZSsTcYJL08lgWnjOat
WJUfqf60p9/xjWbBejcH3lCF/JgOK/BWDuYAdrEaxH8f7AlIAm857AVct092sBwA48n1BCxg+pd3
nhbsue263eu4dLsmmRUVxedsDR61dmsD4/8TqperfiMHUhOZH5eThZWuYcDpR+b71PHyXgudrsti
AeI/865sFnta1HLZqVWiszOldTG5AisRb1/6Ay4elB54/28O5o6L/Enn70A3ulVX64qrB8/2GGoO
KAt6jn0qEbRMJpohhChInfulfuFHaSoqmJDrPaPuY6tJt6kCvowdJqhy6jqgFxHn9yDblRm9t/GZ
hOiba5AK0IP4g47d98Z4jK7KC9WGK5dm+xsc8C/LmTXDxtLvh6U1qgDMI8ad1tLSoIEWT3TiuOHY
2mFNVbisUZKI5+paSJ/VaoWenmoQ3VsVWbQHmRY9AW8RfLKbyF8pqRgTIMUU/7Osk5X2jBWka88J
xR6QxqsMs0edwyLZt0iIvaxBiA/MD0m6W50WdPj829olLAAfLvlnvDvqIICMaye4n4CsP8LlCe4W
fO2OLBzUwj1M3fHZjuQUzLHG9PIG9yx++Fq6EBi1pjr6TTfaqJpMvDqtX5R48iNJufaXe1eDRPYg
/JlGRZNYjZqW81xKeKq6CbXpszbXIIqE+/Pox81OyMxT3No2E+akCia4tv6Dd58EUzjzxsmju8+M
qlOkg4Ar2ASqPNE5PjBZcZtORVVr8oJS8ttjMK4LzUe9HxASNRFyqBZB1ezmJe9gMNM3mVbDREy8
4jJif/MwVaVCLuIgr+kuAVhjhxzA5HMN0/dIwVOUxKGBJubTJK9Jl+awqKYPTjvpUDqb1yb8E3+B
MambXyidy2tOy8w6lELePwBqYrqT2ywyRvu8DwbOOWQMHiNS9d0kTzmzbDuw2SzArNHHmIMPzJnp
w42S/BERcYddFbJbeTUbwtDPcbVsv4F68PYMsnnvNKJEyKI1rQR121EzwpKgXSxt3uyirWoCFDAN
KSWoY21fomqzhHhTzZUPt2ewPpeMbcFLGZSkQ/eMd1lSf/STcmtXB9LPvDGEnJd5ILi4a65k12Qd
SOsmCG0kE82czBPs0shPnzWjYvvDe1dFobi6lBYBFCn5yQn4uRa8FX4xSWB+AvW7PgHkayXWvUV2
j4cm/xTLStxYtUfsac8MGgjCvHGba5iB3mVLPP5KWJz9QhfCLmikLdAkVyiwBQDq1LI4rZUJmECW
fAa7xGaLG21zmxIl0HVkDV8hS0hwLXm8ReiSLgBa0TrIZrmUasVsbqYA+u4mjdzw3KyW1MqsB7aK
xKj2rPXhjCxzN/BTbbogdzu6r04sSOQzCrh6j/bat8iDM5YxFPXn1901qM3ALH2tQ4+M5g4Q2lJb
32CVih0rBfMS4cEP505IFSi8x4N0vEYouaFasUvWFgD6yOtHRIYNH9QWvkkzlkfJsaPT36XY0JV+
d4CsSKbH+KSQxOe5C4kszSJzNCejSS/vwvvc2Y+OuQUQ4FX3bNpy5FcmnRUJcxJHSqEO764SNgDN
6im+wnI7T+lIrEWzXI9MF28/8kCQuuF8DOZ95/G8qCzHK3TFftYYdNtYbA4TI25+IjzuY1WCpR07
dr0fCduGkZXNNCXeX2gF14jVbsHMmF+XGuehfUeMt3p2Rs5m6xz6axxc/DZl4RoBC2tMiGNLzM6x
kx3+9CdktztuT9P43k68CFSqspQ3RUkgpY2Vbi0HZy7rfd2ADg28rdBSDK8n9c4grWsRjgFEogST
M1+Za6Kdbscq/z8dM+QmPFoLSyYNIG6umZwgMnoUtFaQdvohMthB5VfsM/386cM2zf1d1wEkMA9B
eCo/ouLcQtDogI1bv49/Tcy/Nzpa0ZlbUgzXC28DHzV6BD9z9WLXH+IuxZwqN8U/6RX3vROzy4vN
rXc1ZfnHtN0GvqPS7F62yMqnvFz/IEBBnSVCCX2EO/lUY+l0XAAfi7NP5r+Hi03DVu07F0L7BlOi
e9ZSv6hwYPEAXqhKVOizdFgowkextzC0u1rGAcjdJydL8zOBT/COo2RweemdtDkfnmCqlsn1kfRi
hD8j/Sz3wyXukxGdJvgqLFc9IjSMOM1fZuifzy1YddXGYeWJ50E82X+ixC5IlYtgUusONTNtaiAZ
UI7YLgSHK6ZWGXpvzP3oXn9zl4cxnqUNV2UwPNlTEQT+4hmil7PZxXPPTcAnE8jOo+Si6F5mVbQ1
atpoOSYf9hhtn/SQUanS0HlLqtxkK4FucqvfxVJnmfxgXQUfpoF/Du8Zs5mWz7GcKmKlZqe3E8yo
jo0ilINzoPJ+8sg/B70HuMFUR6SZYHqnA3be2yKmi90iJ4vaxMjTZV8cKW3k1aZlScbJFEnw74pP
aoNibdC4XpsbXP3nZA8vZ9GOgfvjs6uzUw8UdxgkRvm0HVMx/xZfG7guTE/e6OosiAa/+fhsE1H6
ph+6EhhIc9jDR/E4CqeufLUwwp0XrnWBYjd/3sbXeaE6aLFesEHjWdfa6rLjuRZEX9OAkq08HLNc
R1JhBNgbwtReyMhTtJ37sEbhi+KzYoixZhM+MsYCurAjHPs6VcuKlj6P+Xr5l5jWjmYinbEs4sFc
JrnRdMdvIAqLOE7t7jM8HQ82rxtHqEiSjWIIlF9hMG9Z8kJ2+MNpd/hBIuVWcLiKtsQn0kbZ9CcB
OaH48cPDrjzzxk2p5vFWakq3q3cfNpEmuRZRtuRfaVDWEfE+ZyIm6mDx+WDHyqBiN/hiruDvnLHE
YJhYvd0ExPeI8y17cCySs2bXslfsKuL9UZfxt+0bWqu7jF+J9ShU/i6uesRJOTXGlQL3sP3VZ9ni
u4K6NUGn2A3XL+6a47wXdDZFl2oUWDlHt8vTrm2Zj/pduV14S5up0klCckM2LfP1ItmnZSGRyrxf
kI0q3/sLZnaLPxRG5qhMmP8ODOrqHefyrPS9FpG8YA+XjPBgEApEZpgCU9M82QrS2D7mnH09lVKD
AKvOGp5lcc5y6R4KpGRKm5S86gxCOb8x91Tslw4YVFZtOdYNXFJp91pL3Zn7uVn377+mwjTn8JpG
VB5ywrH9MNljMNV+sBElioULUkqEcT1cTv7XqIoBvfVJuUdEisl5nn3sVy1qO3mdxBZvDTEgL2qI
MqO4LOLSyg7aVQTqmTvb3rYr+AkuXV/hToqGB0AlwkOz4E0MEg2etUr0IJ/kVCzgw5fuWL+Kk99G
kcvGRVwoHWVGW6/Iq9AgY8Dzj/cPv7lXJdzucF+DMCVJqA8pfoISeCnudstFyqgkcRuRcH8OyAAj
UXVIsSjxSXza3ee+jG6ingBEnI4DEmX7U3RKm9icSSvaZeIiAc+4lV8KQ32RVu75bG4DF/dQKYPo
BeYsB+EvaE3sNNS6qjM3xodd8cb7FCUavWS2WKC1Km8RsF97lb5UqE/d5fDZQfKTH9YZIIgx4Klm
ocLg7o67k9k4ikVrZNl3VsAJqPytrRSMKMNVXMc11PMu6WExh1bGBe5/h9/mi1grVA7+YYQ/JJFg
KbBSmO3C+Jo/i+ZloJX2i9peC9EPZwFiKCqjk+PR9BXWLzSGCDtHQ7XRd0Lg4kfktdmSAleIkbDv
n6Hd/xd9Bg+z7ny/2tnSeq5watQqm9a8U57OY4Cru+djScHFYmwHWUw5pMKocdjZ077yOMnYFLB9
obbqyZe3B/24YnLADqG9XA0W/TO8uyoLUfRT7yCqlnF1l4NK8cuSL0hWOUMWFYqA9hZxLgZRHBmt
oR5Q38WtJnd7O39ZUU0kzHfFviNfs62J/9bk2D9jfWsjddfPoD1w4WIxtr6EDGM1xTdBJWBTZ+Y1
AyLz8RUgZjA8QPD2H2Zaw264cEnLt+KniZFFmqRrFKOzXcO3O7dIqpHsLpy2j254hpmBwwMo/CjC
kZHt5rEy9B4HPCoPQdms8g10oxZFO6/ZPcWe1KdZNeakww4UnpKlTSXdhVcPidRmb2gUxisVn9y5
l6j7K4sRB3rq+E90MsA3AGbCW2UDigcXcdNLuV0Z0mOYjvoWMlu6DrR420a3P25QXdrYfhUHvt6l
FTohwBLjeyFqxOoql4qPBnQ/21J4dIQ40nQCMXch7VoJxyTmhrXfOmKBBfDY5Hu1uz6kXc3puDSW
7ZUJ3kpqzJ6C1oWc2kyNENU+buwqSAs28pMzbCoVmzJRVbtHXKMBkL6ZlCfRx6u+zmg9r4ZQ48oe
11KuLxBruPPMJZ76w0yBai2idvVkrV6lZ8hvcrvsdp112O4lj6aEb7rQ3RShrGLJBPNxYAA+0UZD
s7ay/rz49Yq4NWEiR6bUi4klpLkavwmgCaLve0ek8Vq3svaf/Ll5XLlwrp5LbqzWMIFimKoK7QXb
dyjl4e8XzwWboWpts2qAw6TGFujlX+Lv3bGGxnj327ohbZMVgwLUFAoWZOSvjo9zNApT/NBrubtQ
b72c0dSi6rdFDCZ3+55hm3EfkCEFDzRO1wcS+pkUa8J/PLQ7wA4Ep8OHCZbnHReC8FdPGe8H+CTC
ygJd4S9etrBXZKgIuqklewpJ+0EwiV5iikyW0ox5xKe2ShF7HB9/E6EhI091D1XNuVHGOCOqM/3S
smekROr7UpMevKF0mPSnOSOFoP/OWMH396IZ1vTmmvyFFE/JLIfHNfpNv6pdm9G0PytVWBAbqNuC
ccTEIzLdJO9wL/zBBT+E/huWHJ77z3fLv/Im7EloEwmE9fJxTMXFJK7GE6JeoRadEbJphX1RKpjy
2qGwHvoemeA/iClEnOS030IioeJj+oI2OAd/u34eKhwqfu1zHybYDzL818V9KlJ8UEBvlOBVCi0I
YuB3pqeIzgzZIKOs7cDSwGvQ4/3h5pW/Ei2K6JFl49pc4L0XXg2b3QQmTGpcSMPmAW9HFlC23/NO
ltZHOm9mdr/5aRfHdYsDuGq++W7tgtjnJ2cwZG78HYy6WGWHhS50hDKEvhBNveKZfA62jSYbSS0j
Mkk+mU4kvMqBIlSKqbxZIZ3VW40Fcnke0AQH24zz2WDZbW/5K9nnolkKxIi0phNG7V+s0E5wl34p
37EeE3ejqOeQsWMb56bp0CHND0inhjWU4RDIzRpAaAqLBk8A8azM7nAhFQfjkUJtA00B8JKB5AGb
GOxOrIqw7YS3H0+FgtT0y4u6tlJ6V8zCIAD7xHrt9oZL50YT+/j4fEHWex6nTFMb0GfC03oN/c/I
j7e/mUwG9vJawRT93x/2JuNjwByC+XRoOeMQXgqQcKgvwPJRAO+Bm0hGe8O7oBILD0wFXVuLv2bE
Ljmab65SG9X+SYbDudchHdMiM7zX+IiCBDLHd5Vbq7kzGKlujkKYOJJpwqQsmi4+6IZaXZc1ueIS
QaRjvO6cRd9MAJ4zR78y3W5FqSkKl7voHJ/IaESshsSAqecSsd6PnD4ypCKU9Bj76FRL7/wBAs+K
RFwDBIs6Erkiqq9Ct0MW61utn/ipBRx4y9BCbYB8/zrRY8EfW0zzOvWe/aC8jaE/ymO+TU5Tyjgx
5Xfu+HR5ZpYAwtL/BX5b2c8pQgnwffI8IYEm6/ZoQGTQd4zBZq3TTOGhmtMsG2IEiwOmV0Zj+SrO
+MM9/KU+fv8v31U1NOvHwjIJA3ilinoMZ7vLB1KkcKVZfBTgrbJkoOfna4w/qFNLsD6w/yluRbF4
9Si+Aa3LwkDdOMO63dJS4TQ/F68ssW0VA8mdHXdjl/KP5/jEQ/E7R6wKB01hNWpqpRo9qwSeeoqe
5pbF+Ps4LWTTpk+eaEnXHWfZuHriAM4NJbm3+0AKMZ1z8Hs8EbCbUO5cu+fw6eaRnfmeXA/1tkkj
P1BNukrdo6pqWeDRHHMAJQgg4tF+9wzXa9WxpeBMkjTO2Tvslc9AWuy32iBrfSxbGXYhdd30Zcmo
fdKshPjez/thDfRj5CDrNCCVXbRo+X9Bw+rOdW1Kd8zknrRfUWTyDR6QlHt3ASsClo4OZ1bsdN07
2+GEgqVJMhBULgeIaEI6RiU8rcDSNul2icJsdY7mis9wbOd1Oi4PYYUXlDWNArwq3CzGMXOjQPbP
xK+WbfTpH84KggbZEzzF+dJx8vOo1PSlAyUDnXGQmZy5GLZ7AlaOEa/DVLssy6CFQpqCWRgyzW/u
fsDjVH+kWn3IsguRghQRE5zNGj+D+FNcYx2waO3HmRfO8neM7rdaMvDUbpjDAEn1LL9+djo5+yzz
QTXT4XG6jm+3zv7GFXWbm4Jw5p64nX10kIm5WnoAVrNPUZqrKLNSsBpg91IoQ9nsF5Vr633R/QY4
xdOT+tsbXQq2q+mT0si7JUdsn8BYom0GUwh/aK+fOT0s7/Ud8n/Sb1L19TXpZMKJVJ6qjRrdwpSj
lJ3zSHIvpRoEHrxROjzhIiiLQBFOdwp5E3TJo9Gk3FuuJi3NBWNVNv5I3l0ACVvFwhKZQ7KBE/oD
Pl+1bpdxaKnvy4Qh1InLxNX7oD9Yrl4qXCzFZ7A0En0+49eR1AWFtJRpTpJrH7O/KGk4OHF4ku2S
UDeNCimhEFeSQ+e6zLuQrIdknLn7a2OJOX424kEgoE5D41yMq75WXtP52hgW9958V7BaQgJ82LQU
bBveIGyYyS2FygGWD3MdiSOFFTQdP+cPd7cmZYk3HuB3EvRlSsxPF/dB0K3CcJUlKqckJCGzOwdL
jZD9nghjiXwvauI34GC+OdU9ti8hTc07bQQTNgMCR5h5g1ESRO/fZm+XChMjRt/RBF2uUDFgMqGz
pm20g8SkRDuNpSLTscQbTPY4egtDO8BvCVn0CLLszIPvepOx708iQ5Adj94R1PrVERINTMGhzxqP
QY8BRySdM0nR/ob3PovGBwz/R4q206ZQIrlw2a9vV0rNPH/+Jrir/tc+OuTcDF6lZmUkKY7Eu28Q
VI7S5c5yIKqFtfpk8BBQt9XjuuKAyMUDjLqNbB4lSKZHglOp7pUM8r1ZVjDsh6wCNLrM3nawnsEv
f6nm/x+y9udXT3FDU/Z35bljYuzUpGSouoOd+kcg5J4u4eIoSVZxFgER4zmWcWV5/ZREUpooPJRV
Jic2Ad3Q2EGOqBsU8rJprPEX5v7jM2aTcxKOpBP0gB0XsLXV+cQMU3mb6WS+Fka15beDNLS5iCJf
YHY89j0RxtUIipteMkfkIK62l2IDgfkY4BHnfKxQcMxeuf0jlJVxnFNnUg0zJJ0VRCjq1tFKJ7c1
+JWAAwZsYuq5eT8raLOtTZ7CIL5vyLaBv87UqW6rRb0e1gZQ2plm9I1zJjPLQrWFAFkCafUhATua
bySoiKlvk2KJSuy7MVnFzLfxPoocV/ozNMf8CmjhS8oMLstQApj64ALEfUSHNEAeGJ8HFCcyeUuX
ytvBy7rPS1mm5D9B/A/aFCweSPObdiZQ40Gyqkqq3REbuh0SXsRbG0Uie6Yk8rL/BF58Ch9XOzOz
zFGPfwCM8UD0krp/0G5FD+Juh5tzY5apj3dKK4xW4pG8svB+OJoDnbHuVE46zj1RD6PuVfa3Q+Pw
A2YiTqghhq60FPrX00I5OhHGxD1MjhaxA7vYQhoa7NZPjxrlyUHBP65lwfIQ7ucU0q1cjhpO+4YS
eOktnTbNkQlk1pz1m3JSaxgd/sJCLccjNSyNJTvh0z5NG30i3+hBJJ/QWma7G6I234SbRuaHBU3f
TFHZG65drjKaEH0BvGpfFiSHlJVeEPoTFpTTXqFB4YtSFAAiqDx0AsoryVvbK6F282XVbbhOIxXe
wQqWsKZYc130fdVHxFmfQtVfE4lAo0S3dOJr0VklTGbb0CIoQgC2r2IdEa5txRhWvWJ+XZvw+5TH
QQBh71OxK2ixMNTCz2chcsOaG6/e9vJtjhbvyym6tu8Q7Ayhfir1qB0gmC8MY7saetyepB88U2yg
ooX8Slg/Oy6qg159Pczee1phQIM05YrGaYR13Mjuz66aDQRWGUNpJHinPqb7k7UTfaF2XrIsprGc
JyZsPUwffT2VCQYyutN0tFUaUvsFy2Vd6l7wJEbZWltYyQVcV2nJeojeNwEImNFM7rWIladfsSCf
S8OMGFrunuNz0Qld4Lh5zYkWKWLuhgOfI2Ne7z8lmlfY3Rw6znr4gugkcoZM/ns0p+qGprCEy8Tr
pRfmP6S3swPCj4X5EdCGmCVxMSaSX2Uy6qt0c3qp4vFWdc5htr1J4I7OETKqv32CIM9HCGoyA8K5
PSMbBbRn5XjH7IN7Xj2p1iFxEq8xxkSuk2YDgvl5PGtpeIakolarALC3mJIaWT4gZB2Lt+fdhZCJ
Cz92Y+hCgcMs6ZL5LralRWmOC2/9nKNt75royOUbUpvalkSv2YM9lIujSJja1fyCu19KUryXEJ1Q
4TFMljDTXkFOzURHLSQhVnWjFi8IAHrYvvbQ+CbRGJpiF38SmHjO/NNfdNRqkLuFAAiGIrz8KpUy
coeosgdvv8CXdWT0u8nB3Y/Ha7/BApNXYPX5u9GrqmQDf/7aXIwWHW0OPaMqhaB4lm+cT4Brvhi7
3IxM4JgkInB7KLBVrbWKeVizbAWlMK9fbcH5bumWxAb7XdfAiIrh0w7BoYfArlfeep+tt4ljBv1n
i/H1iAPx2ExVVWvWlrQlkDKKjh+ew8jgur53ajlfmJQzC2wXgNtvvnv/+MAanoVxBziE0b6yJDB4
PYfAo/HvDUidERi9AkSHsPdUDAZeBf0y8vdpWs0satsKaGjANKVNwUur1Znj9TS37et7q+L4sfiw
r2mQl+LzUtWJlMltn2fkRfhg13Sn3+fbdfexoySS9J8PJ+VRHpLhdXwvLO1FITUxFCF2mEaMX85q
sx3Abb9w+rMtkq9/zx+hOM/0KH1VZ7xkSav+O8eOEocTjrN5SwshKCDAlON7lCld4s1x+FNTSLRM
5PHx8hnCnlYuIkIjNjmMjYoYjig/0Zy7EoeZTqf4ETTa86fchr3NLpw5nbCqXGYMzWcHBoIXA7T+
Q62fZIUOw2NMEk4PQ+WzAdY/8a8VfRXr0N4PM+hV5hRoQZUz87zQe9OIaIe94F1sOW4ABrcoZ1lS
7QajmVIoRIfyynw0lU6IeSh9mGNChMNJlWY4DwuvQ3G6G92+lsETaI2dKMh50DQcWUROSWvO81AB
2nz5SI2aXwAxjYN2sqkH/BZCBWksM214Q3Dh1py85uX4pLSPu9WpHU9jpq8/nxepF/dwsXjaZLHd
3HxxPM6on5RjKNLkrvfGVtIKBIWM1vPpaxP9PXRTyVhHhbhdPCpxNWLXaX3Znck1DrRiQ4NY13k8
HuJUYpw0rYgXb01XaZSh8u2wrPSm8vWFm9p7KkB7Gb7eRk32t0oAqW9ZMSaMRox73rjIgpSu0ZLu
zXbLht8k5JoXByEGb67av56zgGLhaCsCVGlNwnrlbFb3xq+Z69wb3LUm5umlDW69ScUGSI5k/jx2
6kh/HksDMVbjRBoxc4FoIiSn4nkaCLz/cErk/hP73Kc+3E7BdwEc9jUW+3U59LO91huLHWViSFWs
o46+aYCK/azp3uVJ88X+bhQUArAQQZXBLSlibb5e45J7rrTbPJ9WaCIYks3d4QxKGyDq6XpoBdUL
y9Z//CurnjJh5D8fefFNEL9/h+mX783DCMJCc3nTvNRNCzp+szcR5C8qyXGlUt+qPSk7Irih0XuA
vnUpCseZMPF+dRepiykXxRncoCpb+y+94qFrxh8M+JcTzYvybke6tXhcRWcZThyQhSZobjTSJJ/J
dJjG+dNm5rTz6t/2qfqxgJg/Z0QovLFDFgCCyxdDCZodx8NDYquOOtTsgnzu4ywNFhH4VQ2+y40U
GHS9paNsTu8FDy73+zJxuzU50KgDVtz8pELETLsuuEHODU7jSoZMzS1EGw4j431QTcb1KIi7bPLG
OkZHVOC0BSP6m5wPprS6Eo310qYV1ozWQkDQpMl+ISNHCJjuK8YBicY7Ttfoi+n7U0j3ITB2MR2R
N1k+IWPyvs6KfM9Mz/0j7+s1YAMWRismkw+d1lIDWa9Larr2j2O188pX7JNK+mLqkFE12Y49uRjq
06hn8YUuBQvB5Eptigfl5/YhYyloXzwdvjjKdMOK08p4YMfN7/r5+9q+6JU0YaXK3zrdAHfftdUR
jHVzguTXjqQtAsBmPbFVrIQ5IZXkX/vHI9nBf7OhSg8EUjcf+YP1dP6Jdp16UGg9LRkdLEBVPMWO
O3YBypeY79kPaW8VhPSMwMyIyQolSy+Ljpx6aI2No4uLsjb4Zq1WnQ7SauNz7L5eIs3AK3W+Z7Fm
foeifPYP8RFTJ11v927iN06FXVIsISiyX671RrMVp1xgUf1Py3/a00iCXj+g4jY4MabaH8Eeqcjc
AVRYYpLAJ9FXXc343z8Rnjwv6Zgi31b/glVUg4dyCvJDqGz1GcZeTLJJZrAF5Hxsu095RnF6JNUF
d+dfqESxjcw80n39Xr3d/VQeVQ7+fKV2mLg4RNZZRAAlZDgmYceDzwzivdVYw5hDlGZdhfEPpBSf
h4ayR9hoe0RyzLL9BWLpUo6lwhemNW9PF1/5mSvBDhxEbxz6srRtrXSaZvalWH1BsqEEDnAcJDr3
kJwkeTksjyT4BoWbRbVFA0T+Z9Tj/jrOl8DwgWVWvQp41A67lEMdN3823DOgjpZ6ET7FVPrL/8pn
A60eRlf+bLdyp/w9t2GV8hNZHp1yHh/uekeN7N7tZmR+BqgZrs03B4GFNPrqLk2bc92LISt/qGcC
a/YBQVq1rq7ZlkLPUYH+lPO6gFRi/ZcXvPty2WITTy2kA5aJG7x2xkxr9WghJ/QkSc+aAZQvRffz
JO2WAMs7VqHemii52BIHvM8RLdH6d8Y7/SyLTr7qTH4eJeNxlO1PTu8xr588ipba39nMnOBFhBxZ
BbyzzYRXy1vWAIUEbe0TJnKvvgkVuKk5CPrRKOtpKBzwUO/WAX+HvgqsoEv8AvVTabA1lwtNV2cD
lwK/UVlEfWfL+ossFFM3LZG+GBnd6wZoCmu4NhnkMLtBl0tUssU5frVPvF2/9e0kHk5WoU6IwOZN
f0pdLdn3JUbGhaGx3jPI3tf3dPfauLKyDnw5Y3yxD3vVj2/Sge4lece5oBd8f6CIGJTUkdXs6nGe
4in/mtDBjkO4mdXDl3RpAp760flu758oKIWb2eQ4FRZeYOwGHGUhOWf0F55wUcwQiVI7oM1fwB6i
eWh1dfwM9F5vEqGrbyxHgAvgFUxdg3qMct35aXEcO5ppPmnu+FJwdMtPX+rqmPN7UKEXUhj/fXev
qvJEgl7Uae07zyEtqx2dkVrrzGUGNWsbs+oA1sUEzl//5UpKGZWFNijYq4MiNolh68wHHyP0SXis
IQHoPtNQIJzSUSgHGO2yMGoLTL4uprt9XceZ+xvyKg/JcuCs8r5YIBAbTdM0i3YKcoFbxL+c93IB
49kfLRi3OeAlOieffA9nyklWyM6Dzcp+0rBcBjGYtJPGkKU4ZxFT7OV6RtCaewWK5pmwFoEyLL2V
TiIujjSVYi5jARhChesMgVUr8j/G+86/B6llYigT8uheSGUSqVbKYWBcGVf8nZd+GMofHm7d0+Cq
DfFxU71NfonKJ9UOiUoN/oGGHVcE+LmoBxOzxMbJMIzyrWzM3gEda1HFrjgzBSEvXVYfO16V4Zq7
VHNFMgNVRr0XMlozwrAj/a0nQberzQOwiMRTBUR8FB5MU9SYvg5CLHL+U2pl9/I4VCnUoaiIMv/h
B2X2ywClU3GS0qk/G9d3gGlEJgMgXTFRFIOb3D5DQcW5w1Kx5SSLcqp1SPBzRVdU+p5rPA/EgzhN
gyJrCVkFsX0yr9V6MLxST/Pm9ztIGcb90a6tQ9WP/RLtu+l/PPnR6xOO2usyK7aP5vYVv/9sNGL4
6zxJbVzzEPDC2roEpuOvJCg3uB9ObNg3jeOyBPKT++CprGTOOw8+jVVgQv8gbuLUWtiIPFDd/ybl
qcU8x2Yso0pgsupKK9R5gduTTmc1neh4/Yckv1/ZJg36jK6OtqUJe6THQBFNMO18nI6QxPI3tgzC
WVnzVUntigs0I/PKKYdIo6yYUTt9xoRckJwZMH7SIcojfymWf4CH3jJU/6OUyDU3QvkRK8JePXpv
i3z4GVL3OTU2wm3tVx5R2I4X6IChefrW/L1MP8vqzvly8MOVT/j3sbkAIAPMQwVxzgHx0PAgjUgS
3ZYON2sfpDvWqrSN9rp2LN9kNlH9Dg0ogDHOamNMkFcalbsOKjObB2ubMCXvrugGVTnOI7UjxP+S
D4BUou8d9LfYY1mV39ufjGg0sJ1VkFIJ23C2QJOWDTJ9Aqti1VHusD+vjsEqmZjJY893C/IQMDmB
AmsCf5qgXiHHcMiD3uSC9FGVBb/OjeHQq5nNKN5a7GFXPBRrnu/drxs0v4mBdh3kvdLbVDPYZJcZ
ilB2McCVArDQOouvvpZb/4lMDaMjfhHYUuZ+K0wRt40idWwY5r5CbKRcLNZWC2wZEyFD+V+sgFt+
CTwFRWEauCcWekcrLQeeqJnLiob40q2GsXkkOj5BjP6NXcbouvYCR4Aob/lLOGssMB6I7PDCM8Hq
5Ixa6WQWt0O5qQ89AcA1PMaRzVbUVX4U4MvKSocx6HOSaEDAJTDicRLbJB+P8eNk2iPfmsH+S5wx
ZtccAhJ1Kl2tIA+7BCNrdFQFdEzF6BJmyJ8mdAKpxo6pfR32XewF6Jxh+VPPtDW+s1huq85QzDPK
IsWYqjcZSEGI6hJkHbpCGKNNEdkWJ9s+9BXkeJutO3xlB5prVEAs4fDz+TsbZwFutvlojgBnoF+X
9qbFuQFaViCPA45RCfpv31Efdn8OXxrCLc6mVmBM4nB5g7L7I51nq03S9X/DFlZGRSg6HldtZ2x7
9cldywmW5yZbSOgWeymX+zr537OelLO5NKo8U0NQZVvmQtWzEAlCdcZG1rlalCIpNDa2JIcCTxEh
dyPnPygIZqSFJSEdc3ONMU34b5W5boO3cm+txCcKcU939Co1UjJrBXcGjOP/zzrLP4qyTkqVt+LE
YRNnOd3GFI8851H3IOHLrxmlILfSglLMwfYbiwlaWu5TXuDaf2BwDFT2bQ5DOI+v+ZoXuxD8tzp4
7rng48piafX4n+XrIh+bxIZ0PTb6tTY+9UPBqrq0zh33NxsPI78j9yLk23iuKt3R2jcKUo+89Nuc
eSe3iArWG++HEZeh40qDhH/e8lsKlT1upmMnWwCAtv1Hv7Epma0cVWD/QtoadLO3ciA+IYPSawP5
94RG54wuAqyZ43sJmhQaepLUs0IujGwfwAdPh3yJiKMBY0uoE/9VwbvcfIoyrdBh6uDrdIfpeX9b
IqgiWEk9y3dMtNFU65LHuZVPjTMVVd081oMCzZKJ5Amo1fO1BkUg1hWvUFDNN8ftb2XQWEM43XNj
cH4V++NTayiiuN0THXqdgOtXl/AlBSYBQ/xrNj022LRdS443UGM0wRlyk21CPSvP36y9w5vRrmd0
bl6Iydcn/Yf/jgwO743dTTClhWVxo+SiY7l4boR5UA10iakEhSC8U/5ac8iY2RroNG6PZGamYA5b
UXneaqDMPCOb0D9XMy1x+6YPfvWIKDC/XMps7Qq0lHaZ6nTNqULgrmv0D5HsuPKU3iK25S/xefln
iWQDoCHYJ52J11tTAMvS5Xzif+VloUSxxnYgEXU7WWyFsdpE3QuxdFnnxTddvuuLyxJD2Vb6gCLR
yeUA8+eHX/zz4oxFoaUPfPoHU4PZfuCZ+/7NdE62i8jguPb+2NbIjXMdrBcC6OckfER/lI7Ptigc
oHibQEll396y0+la0qapsdyD2+vGhAf5zvxLeTyUmyArrJre/KH2+ki1Y0q4ueOls7euakNFJ1xW
A0Ef4cH9pIGWsR48PGl3EobGa878b5kk3EwP/lyCWycMckcpbLFsLWtWmPIyX0FGFV0BV9ZPzKZB
zecpS5cxyD2hCz6t2+GLeTpCXoAsgZZlcAx5m3+If2JKgGGm3Zj4is100ST8Gx60SS+QUM/brjBl
nrbrjLn875RNukM0VQyPA853lEg/NUH072HP0NKMaLIqxrz109m3BOpG4+5Ulhl5qqbg+JtJ8UPi
3dwWxOcWvXwjPGcurtThSkG0UjCmYzfOm/WhDrmNRMxMnG+ARBc4njbh9COBXP4XSvN1jnMCFXaV
f9awUQaFC92zqqHCkYRQQ4nEaJu02t2knWKzxua78sn1SQm5iikPImYCS0ajoK4Cd3r57c08sI+T
xznRLh2lmIQpARDhxNhfRS3sP2w+cPGC4juFvAEi+JjN1xAN0zORsFAPaodGNdjsqmNJvuBM1zT+
A6G7Wi/gttfz/P1tEPGxXVxHmOyV+qlipoTpBEQGjavuo1AJ/mD6u7MvLhIR0QX+UAOiiWjd8uDT
RzxfQ9Qziomj0ivrkzZupSXXc00s6NI2zQk6Yf9sA8ZHmFgG2eo2mncDqheLl8KtEZTCmSQxxGM2
EiNLnvUuDqoATfkF2WApDmTof1GGrC5KlkvwcGLvTxwF2G2wRsipRWBGxjVNOiM8SJQ+sH7rkdZM
Y5IJ8PWxisV/1y3U0mrvK2IJGperSX62LB2exVwj9psb5L5TJRH128lZgEe3Qxd0ycQVXhNiQFaj
psPXL8vjatC8+w116TWzYbXJ4pGlFh6gTMrDwB6IelzNxEyE4amebRzd4/80Ql5QXb2m/olDwVk6
M32X1bidTg7LEcA1Gw5pZH8Z3C6LE0mG5Mlk4+9qidSaLnV+Utnidy6c6xYFpNlin/wkN/M6ZzX5
vNEVGfgnO4/DORgblyPwyw/as6v73zYo7ul/N6hdXwWOzA5bzgyKnxgqm4VNU2Ij2z3SOLiM/Vrp
PUI+vbFqXjHJ5kVurnkS5Qe+ApDnhBuL2QL4+4HfCgolbtlt/xmACSCqm0M0x+kNLNpLTEJj15B/
ZQ5oUVVLHozQhefboW1YzEbioDLSoIO2qjhR1wdo14n21QOTNbj/wid3aFB902uVRwba27hI2/0B
G4dIwNhkfuGThjB9BzRC4pKRiJdSL7dXAM7xQ18VCJd/Jegb7jaXzMOKXQA/ipi2ke1STIBYoy1o
5Eh8nQlCeEKU6zBtR5u5mSaJA74k9Tnwr4wGRHkYLKPXZpGrJ8wtNRm4UT0YKjk8QNRJkXK8spYU
EnfvSlYFwivUA2gTDg+qipO4FTi/Axu7u3O4o5ZZVNbi3C6fh2jJx4JktjatMfuoFIb18JeLVG6r
eZPVcmItYg8NtIohP4GO7cPlxpfxZ0Li2VDeLZhxEGbDw/yDnNbcvSDFlt0sfNwe7fkktxSbCQVc
N8k0uGK8NztlwoXkmjwpNQ01yT9EEE8tPmo1rNHnefjZDDmRr1iRPj1q0fr1pVhJDLgdyBInV+5G
OVMjkO4fzKgO1qIZx0AMOOo9MMQa8o1y2cenDx43hnk9dx6XUNpsTWZn02kz7HV3/oiixTcQ+bYm
UsvJvQWkmsCQKt+Uq38p5XoqNQlvHzdR6PX27M29OxzM6Ui85U+jrj1FC6ripCzJ3ukEFK8Z3gFI
cOVv4j5CgbY7D6fyZOe/pbAVf1OKcF72bQTxyVhb75GIc7FT0AqouzVsqEhlhmAR5X4LLaDL/exD
6smNRZ5xsyzvcS6b7Sa+PkG5SwetiflEHbxnhlViPpxZ8ahrP1jcr0dGUKa/VWwPiZNseOrntp+L
17DBsrZXAYeCQ0CXm5Wz898PyDvSX9iD8n7DjLtz/sn8BtgbfbWnE7QUG9DYuT/ZHtB7Lj9P4n2Z
+We9YS+l1xb6oKzUddwzynunSM7q50h2kZYUrjnSSqyAtKU3olbZ/1jwI9tboaw1WijABxkI35xx
RPZz80eooPBibK1oyn3tCaYwLQb815ylA+HibW8knnXDivipU59ZWC9AGsopwrgDD0EJs1CMFQz7
061Nflt60ZPITVy6qoSqvS5iwuO9BF9xx9jlT3qX+KdwmgDwyEp/lgb6F3v3EvxgO2P9V7OTwY/L
U3Aeu7XZdXZgqWEOWNCfI155fcecMSjLavpbUBAz45ZN0URYKwA3sMOgqTJkwL4X5Yd1p0zj+9Ie
nuYjx9ED+ZFBM5Ox6J9aXYSejqlomgHGtH6md8Qeplr8hzc8zozWDH6Apcn1u/NVImg5y+0KxWZn
Cc9Ilm6lh1NH/3QsOY/F6rVCM5ndqBwz9Kv8/qww38pEOP/U/MlFrejgXz8A9zxJNbk3wqzmSxQX
cPzfnoQ3HB3AUFSJMKbGmupwma/IsxSojYukwz2euPXBEO1ChQr5KsL0hv7vFiI6qFCtkhZI6yYI
SDa6YrqGHZHFL230hF+4L8rddrYSdGzeiJb9jx1qEOppnvaPLAVbkpj2BWfhC5RlqDWNrYhGhNUy
xD/fc+XHXPs3m5IGwvLtGrzQ6LWLuVV/JB8jEIMG4aNUI5ypSEDzPY031vo/L7LHiAAWrSwLudvs
b/SBrmCQABTl2VNAv/8AMHNLnyIjmcYo00C3zyo19iLqk2knj7M5KEatgB1duzH9Ubrjb2EIbZcV
oiwtojHBtmD51Ph7HHolhvb27ksTmXO4SysE8njxFcYLs4ud2AWopvcFx8TQXhmgcwLNvOUYp/6V
mEzfMAZk40dC0QhfThWKLBONlxQ6GezUS6jhfhb94h8/5+4jrtBHECXn2GSvqeirY0FjIzmIrL/0
jpk6P5D0r3OYQ1ZfomiQxN5WetRpgxtvD1ThGwzDMkyc8hP6usJft2b/toZhxoKzGg+/n8BEC5SL
flhtnLLsPGH07xcw00MGBbc4AHrU8am66voE1SmLp4+egZiFqATPjIedaiVh2wnF+U6xoUhy9UcN
MDlbsr9vB4vi+/WEpcKwVdvJKW6lMeHlxZf1TWxFDnkWrNUH3C3HSWFxWwm4vU6tPWi1wbi94mOs
+PQKR+v7ikmMHpWoCZlBDCGKsTOgHNpVRXZcpAPeyd+QLVr86371ScL9+R/Br4IK7j4xa1PNlsXX
IjqoTN75nWozQAvP53fbH5G9H9xJxvWFkfzsKNp1MOtU24hjEa//CDn1fVouseIJUIvJr9lKEWAV
guqb0v+ZB4TYDYWiJ9NfWzY2MwbuwAOQpPgguMoW0gIMbyIEhwXDTu8pk7Xc/u1/elQSQUwUTYaD
EAv4wZRGOBoPIir401tPbIWc+nE2yZvD2CC3uEra0ly/OccheObARO1wScgJBjIN30YXZc6A2GEm
9mgr96CG2J9JZuPOnvx82ax+Ob+tHtfnYo8bBuA4QZamSLkZaL5bOT7yQNujInCFCCy7os1huusJ
mBMAJzaquvpG5Nwaty3VhB2jzZXhDtPKe/7eMKuWFE6EPBjthfLr45YlYm5tSxAmchBoYMvIUB6P
cSNK4sA33kv/d4gNMHjLPZjwPEX3MVw9PDEj8lbxkDXgWPv5Uo4kPUMLg9YwNkL13UM8ktQx4LYC
Wda7MQxDLOgo9n5BX6qPgCy2a3MopNMoX1TDPR9kcQ6Lqp9y6hA8/LfEFsLVPLLH51w2Ooo2gvtd
XW19lp86Epaja8Q4ijWuoQASp/Gw9vuON3kBKrz4S52Zss3FfG4jbhbnDzWn5bhIwT46Vogziq7I
Ja3HyjoZ1s026WYTktuO3XP+nS0EFyhN7AzZKa/sVRKSKpEUi0L6dCB9VtoyrXuvFLWeIfgPs0rU
Z95XdRLk8KHH52t0CAO1v31AErTBwACkORE6c2ZhRJU6yLnCO+KjNMxQg1KeM4TW8GuSEAd6sdYV
c8JNyw5ZP/VwU3F9+TmnWxChTmzlZzt7asNQdhx6eCtAUvvno4x29OcrO3GGPlD+XE2Gdk/XlssH
lwoR04OFA3sRr+GGiktc+LmoEJtUnjT/daHGOc/e/gfrjaxsuwJ9LyaV5LiXfEHUwVDbKsXWeaFd
P6pwOMdyQVMVMzAVvfb5dbOYRomdu4RonyJ4f+tKOGLs9ENRH7VswC4A+incaDe8ICZr4y/0ZcoZ
6mDcOOQZ0FnJuJy9nFqXiE/95YDXvS+0DhkJHPF2egyBTQBsNByOy8Ew+UXAa907JJlOsdjtldKG
38s57DuiFK1t8X57SUHGVA6M/4loGcnc6xSFYyzn+s9iJhJPJoyZhJzpKkRLWUwFUHm2U+XYKhYQ
fbcirEK3GukWnKyx+e4+bpdRwl8FrSnKMqIY3+PNZm1EMoYGcWPQj9N/vdOidYKQoQiOKetouVXA
MNuncFZW4GKn9D/xR2DPugon3e9SxRjA+c+3dfnk2Ch0Dz16VQErJIKj6ZC2JQ9WCzDUkHeVlC7Y
BijzhUy25bipBoBC6ZLHXeNKnEVzVxXMsLkxVrRF2A5FBZ1exIHOMwQu5jQv+o7O0aJlMf1l3C3A
WacZ4f9KaDda7Ysd1BJqO1onWnOeN959v7d2WiOq9bHHWM3JdrApYL91svqSyaALolI/joe/Mm1C
vS8Ruooa0pBLycfQ5PsVEuxLDS/OV2psMUZUdkWL++BY9oNOHrX83cbrk6JKWzOrd5jXFcB56xMy
4hBmrmgGMx7Wp/RBzAEwlaobe3RIEbze/HvIqyTtDVXXj4nNRzWJwAOJGXTbs7UTueJ9LK+hU5c0
CZoPuUuT6vbGAhvWT1wLXeNsVceJieSADSbb/KcEQyFhHrkPmVhuWDRM80ESQP1WokWhDSUxgReL
Vbyntrh+8B7Wxfdvzx1q3EWS9jsHs0pAwNY5K56HlUdLu0ZoKZXbXagKlJVBkJnJwQQcfLhpEdKE
6hIo3wbT+lnx4ezHK6nDtwzZWYZS2PVvgYUmqKmsCoxsglGfKQ3ZBCn2LZxgrrZa+UFKurl5+DQB
Ly0At+ilizJ2xmwwSC7eXcY53KpDvDgSKyqNfxriN6shzeVFsXBE3lQZZDND0KLCW3c0akbx6fC7
hBI7f64DV9Q7SpSc1fwGVXZLJqeMrVYArvsCgo1XvqJOVtN2LT/4qCYtMAcTb7XcZY2M6Krf3ALd
v3+D5GtCe52ebAZp1+wTBPisCbeKwMFbO2ziJRqh5dOx1yRe8lDFxOtQaAid6Pf1XW9UWdrSpedh
C/W9o55Z4u3DpUeh5FIdqZfOUpGvae4qUo3nJLpqia0MZmjxMIvYs6njp6jq8qUYLxUQUpiwyPnt
PA/BKmEfCJKOmKNdNIOhiU5YucLJCnQ0RcGsVF/kUimak2mbfuGmNTd7pks/dwxiJuMjWjjRsaLZ
pKkyr8Jg/BzgR67Gt1kvWPh8+Rl2R/qT8tU0N1vOr4F+2ElsQiJSPgYtSgMIZUak/xWVs6IFJYkt
5I6nWBcs3i/xE5/N0YJ/Omk+Jnbe6wtjxjSPckqFb8BsYr6hSz47jfZ4O4F9W6D4fvE3f7wPZZPe
fZWxn1OMh9UZyfLgJzBnZNLXTyZQb24adQRGLPIZle6M6TExa8afgzv5ODHZl8k1y94sRMrT5yox
aZbdjkLHrVLzM3xIt+rjFXQ4q9wlpzA0yd+5/yrHIjU6vChegEjagEiBLt4krii/DDexG81ltjis
4la2SO7lNQD23uwHeVSNh+7zuswe6EnPHLWs4phyhP/Lalx4vCNfQd8DCWc4nwRiPqmtfZ1s7S5g
/xdBriROzA2JLh+R37w/3YC40k3+uqsJCP8EMBl0AXLT2bhSjplsggfSneewUK+WC0wvik+pvpJ7
33kwV34IUCG/zvK3A/tmX/rwZSH2fseebAEt0+9MK+9226uGcmxGjHYlWDB7TLvGQhvsOxyNURGu
NNGbT2o7AjAHAuqYpD2X4++a7sMIsp2+gYQ8vqtUKXuiDp5tdSALvwqpVPF+U0kjtuaT3AxRrPDc
PUDDoRXaN0lqQMypdg0lxHVb9SbyyaJkXB7dgge4edjRzqPtTmBZkLoY/TWRmtsATAGYLuhbF3jT
O2obEqp5TDcXw5m73bQT1pS9b5CJhN0/wi5g23xwxcfcQ5i0GwN1J3+dh3yWu8cpyGcL359U/GZV
fZLORPvSabSaVQl97DIbpZuBdr9FpmiQecKEG1vWHtuXym5BJvZhRZC5TpfYeH0/7Q2VjBxheJ1Q
lQuJEOBXAtRnM3PWbvZDnakPWdEwaxTfyWFWs6zxfGDKqmwcsrYT56iL/AZw1E6fMk3nQf6m+u2R
qj1LIBDjCWJlRKr+tS8Ehr6fwnFlK9vqFrqGuu2AwVfkifQ2bU9sYtevJJk1dbn4SwoYd5ppMHfT
oWwWUadn29yeAjmBcYkEvIZuPo3381ycPGF43bT+SrUKm8FF/iebmGOk9MoDq/ueRKkMKgtFduSk
VVprWZ3KiRkEnfzzBpVKKcmtmcmiARLeYYfsx7z6H1b2Tw8QSUnGl94ofSyZDXVfYf+0SUW+DC1l
FCh6wwPBrokwzEgOhWN2c2BF+tWoBRi/5qQ4EGsJc56M/kr+I3PX1lBT7ReYo1WwiuE73PK2wGaE
VwucyYen1DvRdq9AlvCnIzZmNGyPNcN2WesWOnmOFZTwjEOtIZ7Yh+XYWHY64+qY+QaB3vq14aPV
6hEhRXgBVD8EWZg87GIq8nJrvfpq+bHShx3Jvlad+3vk8nYbRjmcQyeJ1xq6vv20MfDKXa//UoCX
Wy2pequptDpxBgKui0g6LaFQPBRRKRezJKpB6iAxyOQEQ/FmEy7VhPPEXlGq9HP50LYX/4lVEhsh
blFWS0x35dMkQ2qNE30mq9OSwOQZ2PvVJuG4LflP9hiDt+u4UqPxuCluZLPeVq4iNCJ4IuOiQl4K
QSHV2hFzLJehJxv9OocS+BWkmGiNZ6YzMU0vv4KYmYhA4Nu7/PCErP9HLVXDeUuIlnN7GXcyyN+v
tR3tA12dseN/vORV8QHfC5ZaAMn9IuOE13FTAmY7GDz37Tt6VP10nJbReVhuMI1YrNte4QTKFMjX
qGh9/rSy4XvLyKnRLOZRGwACEo0zXUoqi0tev6JAdJrYW0xj8i5sdiLXThzqpA0Cri6DnMb5ijHr
p2K98tg4bxTYdEZveygXMmJwRbnC3AMDgKCnz4o6mQylbdntErQ5XaJhuugg/Bom3GvM/sPJZr3l
wStLzIi4L+2bDXlUAIoJ+Q8mixs1aXnxCFvdhDEe5UTF+iFlQxB6KEP97SZuq8w/K/px/bs641sg
94xr0JoCzl96FSnl8lJ0ALbiagMrFa7EFknBH3s34pFUoch9s2zNcEzXZRRCs++d+kgou+yqbSjd
VeF7k9cYawcExPpad1UY6iz/vbSqMSj5rhwG92x/HJeoxTVQRBW1C/np5OTvgEYoZQyEI7V6eKyi
Z15/SADafJw5+HfjQXWR4txxvXTVtHsCYk3hGsKgFebiUsBUOKhz6WwAqwI/3y0IdU3++YfU9Yh7
iqJhDjZusv/64PZwuboySU2iXJmrFq+E0j6sIqBKSTY0V4Z3BF6oEAMdCbgEUzmq6luWYcHTbI3h
vEd1/AUbK5RrZdB1DD+Ul8qt8u5DhhaWnw3o2h2R8+vRrdTZoNYked0rig6ADRLKZx1TFGDAsDhI
LFo3phBR3RETjwY4jXg4Gu+e0tAEOEUaR3kzZIXQviSYAJTDqpX4kwtEWRBdetHimnAHw+YpQhC2
LYMw35W0LjMjBC9u7rw1eZ5DxiTf0aiQN81D9AbL/cCznJGMEcqedbsJ/Wu1vRr8qQhG3ECJ9C+Q
iJTKIkGAqJHdL5mP7EfgNzDSZBFbhOq3wVunaN8FuLcigKYCa758BoAvDyzFWIFyT4XV9tpvzIU5
sL37gCEbYv0DmaLzcjZWDA5EYwzigqK/LqA3lhZ4OkoxYmAkod00OjigI5/C0zwoZbxKkg2FGczT
fnmPhulL/2S2XEOC0E5qQuRMsC4Weauwhe8lG6aU4EAfZ1st6GKYuw3vVIChede60Gce3xlFxU7s
0YiLErKsB66KPGMz6SMr/4Ufx6tX3lfgNZcNPzxt/iUci/bIuRqObxVopTtukSGojSM9WG9NarO0
lUJr1/vnohXfYp85hobYjDBVUlKncZl4FXV2jKrUGZOWc1xGH+7mxF4bMebShnLFDNT57HK8gsfQ
pjkcC1HURdbrl9MPCmLdwBF8XL9wTGF7LoIrJBJVMqORy8YmdTWO/VhzOwmI6re+w+K+ZrExXz0a
DuvG8bs6KLt9ODLD3e4fbnOW/VWW08BD0+q9unveAFw0t7yoSm/rVt+jEDUpy4/WxxLRomyPCliH
Qcfi8eIbaD/4zgLvYxcnYxVSv7GvT5+TWUwjqWiYKgDrhhtaKoBZ3TzrHhyTT8AEJ22sq0fXn1nR
AMj5Jc62iL6v0IqI+bLYEB6yiTXuPE3bF+fAQnjSWRxwg/FPI7RhpkP5W7ghhxvEqeaui9WQxMDy
k7vJGZgVYOkulqqBvDvEUITRQvSJRxgB5iVuf5w6ubiXhrCr8InksVdWcGx6IJxsQPSc6hrLbBYM
1sczBaflIKMfM0E/d+WhE4FwgVVqDUM/v47FuUOdyiXsCiXo7kqnQemHD/DK4sEfXNqYqmydei7l
dR96qn6YuVG9W7iXmzvwmMf+c7UZhraov/d4NzZaJKUCghJ2wd0rQGIs+PaddGtYLnL4LnYBivUZ
tpYf4AiV0ch+XGKA0FGdugJDbTQg775hSCzfMSKnZR4saBr/kAQdObN5QevxxBIbvVC9AxRz85YI
B+1lwSd6mLXm2GLa7rRL+wEDhBxfB/AlolfVvEKXZxkQkEN2evZAEtNSOSd1vY4eLkuvjS2uVN3g
pRGedGa4NhZrARW5HVxJVIE3XGOVCYUpAy4FjRgugRPHkc5uWaavzy7UqASk6CT8o4vyl999C+6K
trdqoGPQDgX1ochqK9vINlIGxqvhG+SEZ/sgN0nPRI/ykvdH+tcOKLeOYFCPM/OgtEpN1qPDFtKk
YW0yfxFmA4OzPofN+GReFvOPQGOLdAqYbZoWKXbFlGzv+JgyICwYKuoJm2KmxIW3R8zKpzUxq9cI
i9knKJQ+tZOTH5ESV+mbKJFO4MkTS26ZZX/262SLHdLmsfQtGmOY0h3jOVbW4Ehc9kMQGTRtYKk0
wrbZU4LyEO1fOsse9d+4PMH0UshjyaYiE5brQbejbEeci54txOZP3OCPsl7mTegIE9I8EnKfrbhn
VCO8du6sPlHp+i4JiAF796eWrUANaxU+MY8l/Br28cR274rr37IziR85Z7XTA+8fkRJ57RizD5lR
fKw/VMvFUGPm7oUGtjbL6l0oTllfVWI4rVAjhsworhZOro0ddCPyfmbEMW2BulL17Wi9rpz6As/d
VQ0r6NmmJqmlDsqYB7VBuNcll0SKggEk7LD/yBoTgX0YjLMICjifju62xnChsYHKAZBor7jjMZXm
MtLPYi3zFkK/AJBoQ73UtMBEISG6VDd9F7Kf5Q3W4Wkr55Wt3/N0YptLYqIOHP6g04A49nfdvbxw
OvDJMZ4y9ZJH7nB4bopJNiWoZ3R2dg4wBr46aL+Nf5bWttPH7YpF2dMFbbxyWox5QHgVJkVcAnWk
XllYJUvmhn0npmVMX5XzaAHfTvZ/GO30sFxfSVtVSx/V10hut2AwS8BYTY82FLRgvLnyEqMHH4hA
iCUVZ0OzLFu+dufeGqJv/Lc/8tW35Ip5oqH1M3ID3RMw9cBl8d/u1Uw1N8AxQzwCuz8qNUBWSNtL
Sxa60pKTKfe60Y7ogHeextNWZsj3+P5WP5foRL1RSbwcUge1mMwAtfZZU35Nhm8zJsVUJy3pS/PZ
Cpyd5kWxdJv7KB598WDN+t1C/8sq2NOv4HlQMT9CSQNbCgGZig2bj4zQhKADzztTxvfU9IDS8gDe
htoCC1F/FiVqySEMgW+Up7e/mwVGgo5FN23fDyXh3NmZs1eOF9g3IP2fceOe8OP65TQETYmqfAho
FgixBqDtX0yFH3OmOOd7oUhzKns1Vs7rbQBobu7qjyCSwQiy7AtzdgtItNQseqLicjFeRZXunoyI
hL/Tz+QsZuMTwEHR0iYfJL8KJKAhs+VjTQ+7CTC6q+G3Y7Jg3d3lwAryRotMUh+Irdv1q7cYcKOq
H9zJEcu7XQNIEMzlfhn/aXFzVi8efomQLYjYKT+Nujx7QfhDcjpHtyMbRIjV/N8JF5VmhrjKVuAt
Xzx3Q80nHf/558z5sea1pLHoHFWuMJofNiZZ6+P2rlMwJ0590LqM5HHx0Y4DDokdy1jhvTAC7pcy
vsLoowXfBT4hczWx9w8hk0NRel4xOjxpJcERZmb4fO71bbI7Mx8qSkxhatcPDjpQBZ9mkPkIUMH7
LbPX6vrJVV8KNihZp0c+qabQoCPyLLQWuN0vtBEThJNocAQm9ePDDNhyTJZ9PuNXj3T1nbyYls5J
u33fxd+9tgTZZbKwyFxx3nUmxnWWyzGVwWeJCDo0o5xVxlV++QjeBLfiILlsTAVghB/tAX6qardR
f6bTwwVFYaHwRTu4mPkLBTBFpCKDtZBItt8UEx3DjN37WjNkcCOOW5CGQbADuuYzxxW2Y46mLRVs
/AUdgVWLsAGujNKq+6g55yHs6ev/Xykfxk3b4moknCTatalB90EtwsHMDPXSQu22t4w29tGHxD4x
h+YE2SG1CwyGPaNerj4m1eqXKBfIG4RIpjLPr3FSWzkY0v3kV47pzeVS7vJg8clXXwKE0bjdSpTt
Vi2HBWR68cAA/aTApG+QB1at+bnWZQ7fWbqphWhD0DeiIL0AaZVudsHyw3FiJBSIePEICRD96WMj
Mm2hQIU3rOPSIBxbmXh+qm+DT4J5QbCcfput2vLSFVzVe2xW1umNoYqa8tWOMxHqWHoOe+GeLeEm
YuaHkyQDtwWBakN750iRSg0n9+fmsctTN2JLILk/Tx7icnIMIwYj2N0KMjp06bgePmJZbSk5ZIWD
VnrywPnUoPqf+3DaRGlylIutXqwJH/tEeEffWzXkgWb0VlVNZeKp8mxDyAf1hIWwY7hFZLhxxwMy
n23ONfeAw1B/E3rLuLzFVxXI8GMl2vKofV+mD9vYSNmlKJpPWdW9QLzIF7ymYcw56hr7L8XOO3Tm
hgHZvS8WvRMfFFy07fIeAwUrBr/es4B9c/eLXUfL3Te4Ppg4IEThJI5BtStcVfRxjpG1Bl7bmaEz
4tQd0oTO+pyk6EWMMTMosk6pBS2md2Z3S/OBm0eXE5hetTiPoKVQnBjfo65kv2XETaIIS7JlD6vQ
o0YeLnrganLzdgahNgF5I2u9LylZNVzNCAJNOwGFemeZACKNI2LgWAmG9y43j/K2ozU578y5QgCm
Hb3ubW9JBKnFLCBI6lwDSmHbPuKJf3HmevyboihHiCUxSY38Yj1CDKAfqyKkCELs9C00t/4eL8PZ
AY9nbIrkfhMqpYmfPdqdFQpuE8xF1swhcIXXPRz2fQZu0Lv1o5whJn6bEBYrfIUXhEP75+5jHJWD
YWmVQBRM2hthTo/36pairJ62iR+TSmiP9J+waB09Yj7xe+q5zqViDZ7YZqVFydvImyUPZHkvtoTw
TyCX0ftt+NOnuFo+Tckvuqs4o3jENzMStaP5nNClXIeMmEswLaILhJ/wUmQ/98iqbJYR+XB1jtuQ
fZKWi5g5TOg5iCVN8/RRAz6pftHY/jqnxcZsHNNmSsdSJok/ymD7ouYzVJ9Qm8JKu3yGLn5C68Bj
R1xDeNk2WPSl37IiAxejbaLTrDH/ABljKMu21q430U97mG/sUX915oSu/HzkcJkHfcYW/bxjmEvN
0Geb1nVLAicUsMIM80ONfTlymeQOBFGXHBRNb2ymS1QzEIJWV2N9CQq0LlkTCxVIo4hTa5qyGK3r
PHnxIIkfyendLkEW+Mam2avsrFIpzy6EeTEotjl65RucU7G6L7YSq4opJ0rI5qdecZ9q+qZ77hDT
S5am11zB0y5OhjwgVyNPjmdaipvyqa/zrLmKGXAI1a0jejqK/GJioBJ+HAnyvTVrRQocx4GxbTMK
h8MHk8K0Y+Jd6hZDzNUY6Sk/Zc+VmDT4oZU+mhKXFzKR2T821rX4lPpCN/nKF/7PoPmK6o78yeDV
sk5Cyf4Zj03cf8R18PPiEQfDH2/vivWRTV9YeEd62V08TBnltLQJ1JFxtLvUM1tFeEY4Ayp/jzfr
M/Uf+vRJtqlou5TSd1PXpytQe0XWnMIBIv7o0ZclE/lRCHyecYD+2UhPb/gOAtaDCjLf+EWcWH2J
DShkhwkwZ0JamB3JVsYa/fIiQKvL6A5HUXQALF4PAsIj6vfGh55s6HExQnisTCJqwttCDQWb3WNT
4I7dO8hB7Lq6nqP7jkwfh3ilJvydLaxQAagpPlKoDOChlL6U7DhxOvNc091oybfQXMEfgo7cKm/2
/NUyGVDdiHHgw7yvsuqg+H9MQXbi8VTDLbIVPjlH48D7ohia3GWt+jVfVyWblErzRmr1OnkpRvnI
4IhijEOYWKuT0ZOAPThSWZQPcr/KqJW9y7/ZsPzq1cTpFpKdoTcjKJLrvcnXfkMH5GNxEAfrzg6l
/dADPELWLKnU0LaSQqkmPpVj1KHp1tUwPI5Rk8/JkxiIeemxKgk4A2olvJwIKOULVNtAsUHPbCIQ
c850/+/SJK4VQ9VcCjdWktBywSNEeo/NwpKYiK3ukJV75vGYU1Oq2bZ1x92AWAW3MQLNSj0iwbRk
Vm+Ib3W7RLotAwuo6Ne6lU+kIr0CoOitPwgdoxcI0/jq8Cr09grWHTWX+b0WplzUsbPY0aEYiGQe
rZ/VBdE1idQReMoT4E0PVsPClmX5ykO+eRnAVQHSRv1SmJlu/gzR7aup+MewTGuQ+POmjo0hZasJ
mFH5L0ruxQXumK6UZ/Fc9rgXuhW6+y9eOAMGA8dFEjO1AXDRjUTxUS8WXaAtjXNkYdmV7aVeVkDh
Z4XtdnNtvspqEKZb6PxLbNfst+MBJ+GTlsBSUPIQarFLW7/YPpoVgAOB8bSRHvEuxpGx1ee6QhFG
K7F6khBkj3aF87zCDQwPk05L3WGzS6N0b8DS139KYLH2kdFvLyAyqQEkGMG0exUDKJmrtbRa4yah
gzqgFKTeSHo/bAyWvCxja2jpw5t8PKriBkAoufRtBNs1Jjo6w1BbK9VpAMD4FX8hNCC2mDpBGf5m
L3RACbsU4ghwFYPhvH5oAzhO/ppg6t1yQsuppQj9FudDyrokqZI9vA+/CCsePrK/IIuHvi9DB0Fl
5qCq6XXN5vBUMCRANMQP18gVTwDzRVrkE7r8e2Q+kngcR4mNWnMxLfZak1I12V6KTW1i5kxn08TB
YGZ5CLc0SiaT5TYBUgWyq5j1dmMHUaQc2KfY6KCW/hU4wmiTkHED8PVJ1ONv8YG7H41DOaGgJAsZ
8TjpydPuaMJc62bXaH53GR0qnhx97Tzw7OE3tEybneFDVUQ4E6bBiUwxg4qXWQK1XviINpo/JARD
FvRfQ71TeWOxyAyKvi8XWWvu4xFuAIKK2JWp9mPEvNF7yHMfjEw75KJX6Gd3Dnm/rl+IO193EnX/
X+o1bYztX4V0lL4pv2j9TmLiQclUZssXl6VKtg8/ECquXMCSGR5mAe2IXbZB2KUHJgZqzMFtjn39
tPUf8OzGMByCKMiTE7Uix9EBnXXXOspbIvtIM+7AO31SArjLJkQzdB7OGbYxZNdIvYqg6dqpMRKG
XkRnWNWWa29XtrCTVh4+s12x+94Xnsg19v0c44TattXGeEXcwUxTR3Z+ENRwJxYIjmB3Vmroz7y1
jYfubRLm4Kk+6giC4mChbjLHnl6e47ZQmK682XWWxiOhT1gVjeygnY/Fc/9/PReVDrAqKYGG/5zW
r1XttQimUHjsFQyYL5Qv+dA3Gzu00haEPycm2X+AKXoD2vsskh03poapqIuW/Lp0ns4sWjEH8ld2
5y3Ul5yoA+jXT7sF0fSdUWfbtm4AUoSYGez3RU2sXPCX/XMqz56VHxNp8geSDuo3szhTohYyAXiv
KQza0SWpGZLyiqnCfLiGp7W87gbA62jUBsOdMDn6N/3eQJP1UGbUbnsHFYgMQ9icLX4Q0voNi1oe
VAhkMFFFO/Hu5vnRbwxHHmuj6ViDztJP4zFm84uiRgAP9YFcF9J5eeFHszbF5/k7JUNRkEeS5DvD
S4gNHICrjOuBRkByGi54s6Sm02q085VSuid/9HxHK1QQtKvGg2TRbv4Wi51EI0Xzq+JOEIP0QZcJ
PHZj3tkZLrtyeSP45s+rVKSI1w0Vmodw+YNLw6flCHLPE1yZdzhD2+TTVxK7gzJFEt8htUwB7NZU
CLo18mqhflOj7f1gjuoayR3Wb+owSusZTdZ6imzaVpMmYlYvD9bhpYu5r5wlkqY43Fa+RJw5btdI
ThgQ6coW8PxSgxiCnIPLPRKb+7affFU5keORsb5DyLYZNfwjeWRViJ8l+Vcut0Tgba2VF5w0MbXT
FWL80XE1xHVJy4rHC75/SP+CmIjBYFaqkI1H7cSJWw6jidF/p0uoaiZnVSeheQdxpwK6Hz9iYueH
v9E0Onm2Aq6GJSE84N7bNcX39IP++VAMYh2BZUlkPmfseqGs+6p49gN3HnJAZ5Vb1Yf9q6mhV4Ud
x6uzBiIwa5Ml+M3whI1NF/P/0M4uCzYV+p4LhFb7txMDURvBy11mjmEvIXYJKEefDG1c0+5L2DOQ
DhlrDsTRqWh7fequVf6ExepMzCsoY18ADueNRl40by6R/nTDcjL9hvVRYIoWw9MdAT3rRIYZXwOu
WSJksUi0cYkGdWCb3DKBDR7d/aBP68UcqSjjI9tbYwIQbJMRyVCu6ogGddEBYPB6kjwG4281G38W
C1g92TAsX9d2epjYIKr8kvubLvPSUPHr7+e00BlAAPsJPb5Ban7S42JMPYYNWbNwopZFA5Ypu1Ci
0iEvHB4AiwTQ/dOBFM/RopBp09Jpk6EMitwy6k7d0SgWhZVLAR4HdpcYkAm7wi3nh9h/gdb7wkCG
QBL1zi7gfFLH2usWfv/957U4AXDznRgotF1qGrpt8om0fe0H74SWryX441vy1wQzq8EpxO0cY6tn
PYsatz5R1FDQlUM/EZpbYcfBaxtUwvHNXqZJCGTxEH0xV8zvV8OA0bRyCXVb4k7LKeI0DeC5ss3+
Z9JavOOXXT1+73fmLmR/imqo45aFdA8zbeBfjZ70qFVSZedjbwXJycLRcU0ABFFqaueNLnRmLZFo
4cGMVm1kHia//Fk14m/TYbI6S8lXRKxL0Qt9wfgsJX4BhRLuMT+tzbF4uHcwsRbJmCVuvhmYT6GX
JPPkxO9jdQNKvpymoPxi+FurJ1PU0CX70bhqEMKKCnQWbW5Eb+toxk2/d24m+vH37ltuBu+iIeP6
KxunUhEex1NOJAdNoqiMbkgwUICkzp9vbL2MPGj6paq/SaLk4D1GH3UM9YKTUgH9xmwbSOxmzlSm
90psorV98KV4R4iQ2Wf4TF2AsCWGH4SgiWSefN+cQp0B8RdJTwotc+r2kHxWsG0V1/+wRyE7YM8t
e4mnlccVHGc6AlZee8UpjPlnhSR3iwOkegO6yh8iBkHrz9N1V+MtvxcortE1+IBxrC+F3Fi1wIBt
Yo/gagXepi8Ry2gWacFSvFYwP+IjM4CQiYfDafjNcvd3E2yWkGHrrRm2C0hO79HQFqU88LuAyQIR
V6tN4eYaEPJktMaWQ/LUbcINzsixOduH76RkHiVpSyluA4bcq9vRiRHRohJ/piPQpAHCM3gErMkm
9VGv207ZCM4VaJrj/flkiblnNoCBHF1N5sAfbLpA1V5camnvYq5OyhoTZEoVUtgkkCpIvA7tI6SI
Fwsvf9vWP7E4xaEE6Ch23fVRq4OjANlzWZSeOGi2+mwp1W5ZIYWr6ksawz5uJ4MVABwJ17CraNkv
LoDP0R8TNXt+iugghg9UjFrLv+wzjO1rh+DuNZ3LwZL3EMQaDk+JmHvL6OCueXG+gCq6h61+SAZo
+P+sChQ3p88N1jf5sSYRSgFqjhLNrYS9rDFXVyA+jh/vk9N5gUpLAuR33Es/OIbdMmHaH2q/rKt+
/Ox2dQBtoYuANwQZnMwYx5osPv9alNNQ5vRxZmBJEFV7eclzPTcP63ZiDzNUzdTuDx4LeqHBQ43T
23el/9pbvyQKcoUMZI3CZWMPmZB1/lkDu0TLAHwLPSNk1mFiSglomrlVMY5eUsoX9YcnTuHwXqbz
HlFFSxErKCkHX6s8YDEoY1bzW6GtivUlB1aupgWMHsMX+NA2uyiDCBW0Lm9LCgY7FqymRBPXO/T7
M3WeA447XTVTFQbVSIH7DE6SQUbvXO1H4n2mpJxZY33DxcykcOWkALsDsazayKLq1zzm+cfQ0W/I
NzDuLHnJaLkH1duxqyPTz81PsdUAFckhAytWC3Ta6nJYjpjCDw0X9hJBEdyA/xYLKS+RDFjdk2sY
tFoISVLV9/Gbq1jZn19ks5e2kXqlXYAx0nS68hGwFL2QjuufRzDimXiS+E2fGxeMRjqsBJOiv5zx
AmIpE1G+27TWhmsmQ8KbdCF8uSNyZldxkwgoU95Blrwasy/uqkbOz+lxOjJis+0dy5p3rifOXJDN
BzKKOU2Ywm4+NLGS6Dsu353Lm8t3jHXD5zwJ9ku7+IjZuHgBKpU6nppOXJoMIqYyypP+j2RAQ4jO
E5YwJd77wqlN26cycdsZSjDP757MNTyME/Vz2yGFn4HfYASwGO87+kLZF6Jq3FRIs+VuQSPMmiA/
etCnl8muzHX1Zwm5HoJQklFskOc3wCpykZawYakoW+cSDDBLdSCLGSvUaUSSt5P+CooADZxSEDs3
AXl+VUgvG3oI7WYPZAP4sF9yMmTeNioTo2hkTfHWKj24LcHLOtPs7Ik7MJvtKTxnaidHh6uthL8f
fDAOFbFIPd72L8RLaNZGMbEnL9xOcgVRNLofHZWFhMIkwEXEw0LIEF0gHHLJqh75F3syLeB4Rguk
6idpF2dj+DGa6zweZUsDcX+xm5HFH3MU3pCtCjXcRcARqC3BVKRM2YpoNNudW8ugSBF0qYQpBslt
JHVh9NiA0PeCbdQTZfxB0d7rfljtMlZ70cfdWJHWSrTRCNgQJ7gFqZxyUoprAhEgsx0PTNzcTIWO
ztmT/v3ecI3YV9E9u2uXXMJvMQzD+sh1ATb06ZyzosC7DqjJInnZvheQAY3xt+GEXuSTAy0LmfGj
DXmkHHaaFpTw0Z5qkbNYNsMq7CV47NRICgHxy/cmt0CsZ2SwASbs6KMjHEBaBOS1ZiuwnvHSn5Qr
N646K6+Gz0GmfvWobfSXrjS5WQ4u9o69wAv8ppnlWWyA3/pqE9x3+3eToZhjIdgUVuNn50hFCsnP
bcKQJxvCM9twM3yTJEFGMZI3Sr8NPqUdUckpb/B8A6C38VmyQvXiwXvuERJg9X3HRobhmKP/pJTX
iNdCAwynoXw6/Lxqu5tTIt6SPkOpHW/v2H1ORaZSbOlzOqM/NV54fcIE+5ia+Qr95htGwfY1Iyji
65Jyoko/w1OlDDr4IGKYVCLozOC/c9g+HNewC8bsTpkllD2NGKyejMW5sdRU4yX9+f0FJMv7IBNt
QRAaPXTMQ9x3EItt50T0cXFp9ODrBwhOncxfxUWoLYZ8dZv4fkEUZjj6WPM5+eaxD/g0uWCUV/Bq
iG/vhDE6ZV5LsEn5pk/qkaz1PwXPPP+FMEkCs8FMB0NmJHsAugbmUTjHSOGjW9hsAiCCsZ8sFzCs
d/irz3y+D7W78py9E+CFMExTBH5s2ghSXa0Ir6F9z42Za5Fm7JW1OC9kKFC4tzHAuBMpnWkZXz5T
V8VCie+36JU1kGVS5K/dAjqID+ffjtLmCu4SEi6ybNLJ4dnzWuXpgNCUwc9V4/wRfyeFe1d2+Du5
d/KebmI1QBrSooekXJCpy5FzgHo1XoVZgl8SF3Bq2Nr7cOH9soUk6L1m1JGZ8WWdIYYXG0KdaKyz
eAOkDT5NcckabI6ykRes173QYbF9QSfN0MZaGj+t6rtkwpddupkfdMVQVV6Ew9A1WHOAAxqqMrNJ
zKKBbLVM8yFbblGj7YQz0OPddoHsuYosBThmo7PaEqJexC8oa88cn3sc1InuqFzkjcnN7JXWphRU
BNdiRb/V+IYoYAYjl/xBNEYUTWtdPfjJZx+p2sHPI7NmSJ+HZqqHLNAwGAvm4j7L5SFyJoDbv2KC
CtIJBqkd7uSiPHFmUgKWfecLiBW803B8Ggvrn9Jr8cvTmH0uuYCNYF70VefUOn7hDPKheLaWgUG3
mtfGwnqKLFjJHTBdQ8cNqYcJoXmQAnzWs1CAnBsNCcRp+WlPKgml0EiNMZFzU3VJdg7Vhe2Gemeu
HkFaedSfCRbScb3wE1RRw16ecKp//DTgxn6acNVLvCAURYdoevQXbiw2uLYEuX9WHGY4UVWmMyJZ
o4vzj/dxsT6YBHX/qeLwrSXv/2V6WwJym5bv3X+K/8LXarlGdmMaSuSIKlyo/xECaF6lEiwU952x
0UFtnn5uIyfwjnULZNDCTtd7PsxV7w30M+YHopl47YgAMK7sA1hrNnexj+BM0yr9eGT1rxAtefBL
fU4SLvDp9xSZ7gDCzoxEx4sF52dBT+yr0UCcbQP+1BRD0vl+R3AHzkouW/hRVSDr7RyggPkf/a8z
ar4fh5HHyBTqev7nlwgnq/rpTfqewZEnYaN7U56a87/RBGqZGwfAVz8Q0xvqvFrYURnd83rUYqZx
crOAhAv0r9XX/+nILzoPQCZbogVLHYZD4NJ+7u7CyfQ+MQm6Ft1QCnWauu4uaa3/MbMbTyk9DL1Y
ZVyu6h8PcWqPwb7957uHQZU7lXJQ8ITsY6+UCDnbA9WUMm+o1FUsd0FWsjmB9iGi748jAWXFMse8
V8sQuwNA1q2gyj22Tgxp6CVCSUKZiwtNngwoNlVmyZwiKaEZTvl/rST6uzyjljUdyPtwSr/dMBWc
0wWwCEy94ycxu1OlDzShVu7OP35fUah9YQNN7esqZGpvbN/FDsnQ74o+LQjQeENBGVHfj2sMh4ax
SRFut9icQSlFKRIwR362PRnE3xKSTvmdXJCQrUBdcz4LhIBRvmSPS+Z+7ps0fGyZIP1JBdO0xmwa
f8ZCUfBOMAcMlgkw4BzW6p59tRkZKXioQYtJIFhtYxFzE7GmYCXG73j5G4BDmKKLTWyMbl7mcIE5
SPzsiuGXimyv9mTxGVaulFoDHrUgbSGliel9kldnbivvAT49KM4HjMUNPWZiS4fcHRdPF+x3tjLH
r+R0YykuUmnnRfahFhbIXvOcXLA6FgBmW9QBP6BzydwP45TSh3VTCg3f5+lQJ2uJPnt2sVeDDVZh
ZKpOUolgHQr5eNEzR50gMfN9iCXvfeSHyjgZHmY7aBRX9/pR3MR2H1CHI5guodDKizmdoDksZKNN
m9cBSRojUqeTwAcqa6rLRbZ8RzCmRUXOmwsh5ivYEsMVR9uQBMfAtI1npxwozyZwyzfdmXeAThDl
fb19x/eGOqMDFp0nHMZoK3yMag6nVVEAupCXZnCV9EUu8wos6rTo+0YJ9nwqtN5T5C59i4X4ksDg
+YyrAVLo9tpkwnnYarpg8y7eiIDfxJzXqUICKPRMoSNf1Hu9KZV+0qQApLTmqMQXum/JRyl0HpdK
luzu+/sI2zP1VhClhoPVCqA5UFz88l+84V1X4xn7wKbi4/XQ59IoF8J4meovw2qLF43YO23AW1KW
29qAQ6iWPRDysSI6xXYiveKLhqmzkInE/01/5qrRJAu3a9u3n/wOesQDOhS9a7fNz1bMOEPtX2LB
FVfQ6w2+eG9hA8pq/S5aYaUD9svsgVUwgiiNJlFw9kFBjk5g5c3YyoinnNwkM1Ypd0NBhFTEIRtQ
sK5EIujkK2lATYWlhlROzPZZS6EutwcK4AlzCeWgdJtAkBicIlbDXwlaG7CDLHAGzYAdBIwpxObb
RdyeZR4kYX0HWoxT+R9624hC42GtSxXyQ7JEyRx/SdGSBjuQEjtuWn/qjeuKdBO7vJwqS5qdOXNJ
LGJBXwZfqjmI0ssi4IBXQtZ/Zvor1Pzn7TtWqYWkL9tV9u0zRz3eaC3W310wfMZbmJt5Ewpu7Iqb
kgrPD1caPt2jmogmYPFqBtn2Rx5kou7gxfs8zFPH2suT/p+SRza9mTJI6O1YMhVYt4b7JTFoVxaB
NawwDKqwuywK+ENurbhVDetMzGn5xHgcnXpgbkJ+WnVyJf0Dm9TCSIToXqRnLccc6JPd9swwxDFk
D3bS4x1BLXXfpMwcTTu640CNIDszhvhEhpvoqzdJPIrJEv6V9TiL3SOajAg9WLyAELujin5LalTz
kIIZMBH+HdZ63R32OjxLBIlfXd5b52infK0spYH/Bc/veLAqBNY8FI2dtIov2GX/VZvB0j3rjrjm
jcRFEfv2j9Hkkwkhg294CBsURdI5glMENyrhIiz6gBsIXfQpR7dQkSL5FpvDJjozT8i2cLCriYEu
gmTuZvCEYYsHP5qvibazE7rwmu4SXDG7yQCX9jDpcydvCfDgJF0oD/cla4xZEZ1UN/ZF7sgAI/5/
5pzNKHk+uiZvOtPV724qdROHy1gZnsDat8X/G7yU3+ldLfmP1zmKcyZxbWIgNXiJHxo0xI3ysY1g
ljQ9q5U7O2EA+rB1gtGz4VS5H2YFrV95wemg83to63MxejKyAq39by2LHk/wSrmW7YpzKo6GTsk9
FcvFSLxY0zbShQE9zafkUgV5ibu8Dx1Y+5+1NmFjhiMy9Rte7saRoVJg4zooH2rLD1bJ15ol/88n
+Emk2AN2GFFfRXdGF/cePg69ObErFQeqK9eWsNISszLobxfK7ceU3Y9WPbfqwbOLzGKFi7cdtw3o
+/i+jGGLmieAO1JH6lYjK/bWPi3JWqFRI7TksVz8vLNinBmNHaJlGqOEo+1qD4PPH/5hPI/Bgb+y
M4vu4yfACFL2nPo/xciBB5afYJ05PWs19uw77fR/PJtC2amQjn6bv34Mhsfp5O2Oi4ZKEcd3CICH
be3ddINNpsqugqfGwVH5Vva6giPYQUZB6PGgEpsPfdPXgkT/Wbc6m+d0Z80b1uLNXB3Suu0Swg4B
kmgQAbTCD5V7/nYYLhdDhlfZcguHdLgfZ0KOBXXgyuIdBc/HQIPTQ0/LcHRuTNChjcB6kSuNJTQA
iQX/2XDbQZcMtW1MoSjNaxjvoc43VgcqLMpdkKWTSfJJw2Pq+37N21hJWWMWV94IyQInsAnYUNkI
bFop3HltqnczQ9GhDVxenQV/jJcz/O3s28uxa76olZiPQFruyRk4r4l3z/zqAwBDjtbpytcWxZ4h
HmxirR8r6zuPCF/wjktADrH5KwmODaJ65DAlVFlLZftNaEM/Qn3hTb41H9EWEA78a7Pw1FDEcgVa
1KlPp5KR9RIo0CUw9a1X7kDApNxbNwGqF3RTlyRbxGu6USIOI9P6unhgAvMGgDHJ2ptA6ZoNzCIJ
GvBB1+g/0TTNMhA9uS8qMFTApWb9AG/+2z5y5frCRnzCByLhWcLqzHTxxRlJ0XWuHwcM0HYdcJ+s
qhF3wzwxNPSnFaG17tzhWsX8G/JQ9pN49oBoQ2ehk+TyE45iO1gRwvHssNlxodbJRuZ5fQ5itzVi
lJ7tz+D9XVDLDofjGo0VrvfF8j8UDSBcFxth43D/pV8UXGyydPKAD3fBYGKOTZ3nkNFb9rMp55K5
fObd7+9GuSAjYbiXe5J2FidCp+jF57MmCfGhLEuQtot4vXBNS3N1nY6toWBo7sWZBKVDysTaF2x8
AoYiSjz7ivvsteKzBWzdZCKhdP1ta1FAglRhdZt6c1X+BTf5kgEE3gXaCBOBGcMCPKf658s+xd5E
aNx87lOU1Y40ahCH7Bx/11qhPsCtmI9TpcDb8G6qEE2xe7/QB3yXGG9ABakpTSyYJz4ligLMLFV4
qVipHpsq0Z3Ga7xbJZD58sMGMsT/dQB9ga4pLObsnS8/Nzezloxr1F2dCuMpJD2C9ukihMDX0xv0
cscJDomsgt0JEzXri5w77plg5yehLCUG+9jysFUjGhI5Fb2JfZHel49SUONEjYeZqZRMA2D5vrSW
/FYA1fygOfd+wCt7QFID3NJX8BgSiB3S7rwceeAspTQVcYlYg/fDrg8KR4mK3wLedrmamCnGAvYa
EfCvlhceo1OtxtRXgI6jdcflyQ1jXlod1D/ucltzLjvyzHipgch2gjMTkWeokIi/ZvmHdY+JJ06s
0HHs+E4f4X/K1y3ZX4v5QhshZ7YZ9/xiwr5Xg8VLiRyS0iY451db2LQ0Wj+2ygiJ+uPqQDgMvvpZ
+8iyvIx55wEK/wUTsHehIOPPnE2UXB5yS+1REGzUVAt6gTH3JR/AlIggHO7/fbJa6LfyPyuhr7at
+8MKtx1ucVPREu4VcBLgKpZ08EtRgVsX3n3pqVZvPoq5322jQW7ak8Yip4+cOkRWxB+LZnpFqkbw
/gy9bs77BQPWcPfHbKwrz3zUH5PhUMgTQ3ZI76F2a+sou+3XGYA92Yn5YK1pE/+s6TmWXdOX3S+R
JmC3tV+szE59DYHHuBaZfTDCmh96Rhs7JB7mq6GY6B2wS3jGN9Uc8zb3ebCjtQ9qMrr1Vi9erhBs
1o982P6eaoy3zc4pF8oAZLsihxiJacp4ymW13qh1CQODhB4OWE9XMnxgleVuqTB9Jpy2+Q62zx6D
jsTwQgnLg+n4q6jz9r0gSW9mS6D6pxc4Ido4rR118ZeGwktd49qSyz98XYAV85qcTtLI4B1eAop9
cs0MsnOzz8n6rtZmQYkmFzLav682hs9hd9ZXr9TZ4rgAYJfs92wzRBUMEI2xhmS4wuuvUwEIKFX9
DzceSycInJakWcJXCknX+ByfVep4xNpBgtAFF0iQvLBjAXftbu9vyM73CqfxDDBy5q/2lCwy2SPj
6z+ntyZo9eEwoMsi35ApQufkOTgTLJKM4VZP7v6NLt2ab4gqvGCe72V5GMZx0lOgGjC+PxTywiGI
0T6xUXZAACD1Fy6G1F7RQDKZyRAyFcNSP1IpRl011IpvvnCKfRU2bHY1hP5jzWcjCRey96DdMqVu
4ZC1KZNvFvklR1YFcHg9PhLVFpStCyKmXIyGE+f7PWiy/ZRlTAc5/CclzQazN+evo+0Dk4/hQFJF
4avmvp8JhWVbmISS0htTEMtclgjOlB/p2owuvYXBie8MRtj0rf/d3rHgLoOoKyVp+pUvTNcShRBs
tvGINcJJ+cXb8Lc3znDYgSTuRBJ4Qp1tD8uoCi/xlA0Aclrb9Lbs89rjCDrIVRIWLtjSICMFJAei
wA6hb9Kas+ZUWWwqDv6zyGlrYqRH8xgHWsKSu+7u95Bh5FUDX/ndVWHmxFaKft3B5OHE6CxjT7tX
eh33LW2uQRnAXLxnv98DPhpq9/9ZbCsFnTIXvR8+c748UQzMUFLOaJUVyPwW2+DTQlyIuCCR7Xg2
ZTkZ+1Mmvec6hretX0hawAq1gmdU5jFL3dwZ7jK4HlAiSlgZPlTgMAG2GnTfZM6YZuPmHepJTpfx
du5JTLyCVuFspGbTXfWuXASoqC6zTHHPF+PD9zhXUpSTgwYD51kc3NZOJ6ULjNb/Zc2PSZ/Z/6mI
EDupBeBR7Na4HUDyTtqdyCDEmHZGjWR3iNHGi2IYEp/8QOdb/KGR6RLkbev1VV6e3WjQoEQmqoSI
9j/tUWODHAbHXbaBS+roBn+mvPP/dlXaae278KkYTZosfCkWL4GuLl5Z9RPscL76HQOd4QJVIzr2
3pa6tT4FciHHlLGzIpDxt97uMi7x8d4GyLrYWmsRR/i0mVZ36Y6hxo6klAdo/IzKOjYlPL3MI7pD
cMa+/sVyYVhBLQCNcqAzP5/uIl4G8rnjd0JGKYgb+w0CflLeOqVLn4S3lirxQ3F2SJBG42+jUz95
cKEXIPTG/qPySOuJVguiO1h693ZSZ/QRJK+F6rBB2vdh4w4xIFVdF/j0YrMLKdbe4TzNvTL/9ecK
XEXptpEhIA/fEVs5Lv1jC3t6e9UNA0LEFFTBOD37AnVkDvB01XOgwK7BBSYptwPakj5F6jl8tG4R
nwe+Pm8FJBRWhj46GBDMFfeCRf0oYetO8r4mrufLX6PsF/7u6CWEEnmIHtU4MsiIj3coK2nVMjq/
88h2/BbqUFi+i9NfUnxGCuKLCsfcXvVAmXJnGsNvviP+Nz1ZytksHiq9y6d1Rvxolrk+02prq69C
rCEDiPE8FdXF55TAmrogcbhi0GAiU7RY+JpyCeYy2z7y0itCq8NWEm68P6r2Lop+uHCB8rCd3QC7
5iXXa7hWdNXVRDQvNUQBERj+W1+m2Hm3bCwu1psfDx2E77CPYX29ABxVuq7psj+iQepFG6HbOFq0
bDsTvnZ77kkBl4lC8bu+RYgdDELa/G5Ah5Uyvk2HVEyowmwOdQpwTWqb7608FzhF5fyrPdBLJPQW
Hh4/cAzRkTczvlFiUEz512UNLvkzX8SBcdASVo89CaFp9/Lqz/1t1xhpE1jGhZuYe6RKdzzXRzco
f0CXi0m8g0Hhkir78csw4aiMWZDP37Dhosd/hJwtYssoqJ8m+IY94kpqYUHddoP9Mtm+U1XLlnOo
6ZoNPNHqO5BjoFGThglZmG33H0B/02qxrvFJiZV7M1vWTz8D9Az2pooPGihwbRR6bWUOUXd8BsXH
tcbvC/beJoJXJbm70JEjdF+uhj495Vtd4d39mITjERrk2/OMOu3EvXV+DenjvKQZNLdBORUgps9l
+oReUAI8NCiYiKihVbV2AZU/gk/FRgSG+7NVBYKfYdrlp3I9oI0/55PEhGC4xFUgHVEV2x0xTU2h
OSIE/XoiXFzS2CUclhVmRtUUo4VMOy7H7lj073iBPOp2NqUYjQ84HgDcmcm80QFx2RkABCpQFYhY
BDX/h7/nw6m3DgLKIBcbbmLtq1mwNAPYOuprKoIL6p3lFJUp6hB/MDlShu26Y+XSbeasu3K4DE1l
ISJbklzC9lzOVlAsi9tW7VxNrcQAkbUx2G3jGjsMqmyuqEyTBEbFUSQ02HQDnTtngGmlVoTBj8Im
ksJ3JN+czdV5pGbuhJm44m1sXEzw+YUsT3hGvAP5RLLXY/4VsRKh/CZXgp+fxnIrO38QoLY7MQOx
Ro6IKZokXT3kvUI446YLYI7pPWDj4Nypw7TnV529k/holz6/Ini7ptNbdH1dqeaZiXG2uG0BmKBM
HF4Adu/Ht7DGUTNCaZRJgtiK6FQKyGSPhS/FqWGIXxKfkGAhyLFuKm2vYFLrUDcu4SxSi5aDaOYB
7duOrT2Cb0TkJSG1nnDeLwhgs1pDI6rGKT21dpjCamXMSa8QxsPW4zuEZBBYcwugitBKwLKvNXXC
b2N1h40byjCU4jKYdBiPduDbvL6ZZucd0e2voHGYXfH1yzCWO7aXryBBfoI9XHgPf4IAMC0/YGjw
H7f6WbS6LR8D/zJktnbOPdmsJ4kIVXYOmjNlUrLHgxQk3aDi21D4qsrvGPhruochuFnr3um2SWeo
omD0u1v9Pl2MPWo+VXLY7p2LDuYln+JO+BtoHWyWlG4CKvgf4XdeuoQEG5HQXrmUA/8s4IJBN1cQ
tgjVKEpxc9fL4IwX/W/dnS0bE4zfQ+fvn6nfDrzMgC0ft+PbJbnz4YOvCvCBx/qPFLhUnIuWNr+s
WCWr8rqTDyEW0Zwwpa5mnMYB4jP9MSAMlG66/L3usZgLRsOPHe5UeQlqqGgJtk3e0GF94PETfxC/
TTMHewmnWHkU9cVpx3KV2caDVeTtfu6yHIPHvtDmN4gJ1alxFdUxAW0jLf9rQdthtrMR5hKhkyo4
3hCbMaoQKANYVpV4Rx8O/x5tGf7yr/YZUm3YBf3dM8KiSOkfy0+Jd7dGQhgbZIPH26Q9VNipbgpW
nd2xBgacTAFkzvUQ+Gq4hYfhVZizBynmjqWygdxm1Kj5HS0XkDwx2FWTAxgnv5XASRAiknN4R0+U
JNYzeHol+ledo45w0bMQjsGh2sLqAhY9ERyTbj5qOT2P0tDsouHKmBaLPmHSfvK8zDL9oXYaoGj2
i2sdrHFrUr8WKOv23LsYLUf2UaWFLOwyCROq+1dpWulbZiDjkpp/Vvvqn+Sj/6CdkYff/LmOBLgx
Fq4cWCYKCjKyIfpnemndYN8uoDgiWBypRpCmC2dHxTakn0GPssrJtU6LuBV6omdIHrMsYtEd17Mf
fU/qGj/WOA//arIipkMd7pJrdX37OYizGJxMDHatadIm+Hm0BbdJk1ShCyeb+Hd1n3hTow/InBtk
TwgJSEPVX/2GhKbi6MZ4vPBfQX9xAP9R6X0E+klMSSEvYq29RKb/shvmsO2F+AReuGRELrtk3bTd
68mc090tSMloVKOxIEgYCyuasJOV70wywuS0BXjI6RVSMLS7Z/CsAt1E9sVAoH+/D8Tc9N5u6xza
2swhoiv8vVhxpMUsJlIWOdSOfl03rllWAvMfB2WkvJ4JGllplY8MRil1EJMQ1YAYgwwa8RcaKeFK
L01Yr0zGVNrHhfNmZqHRo8d8Yok2B8eK6FuCeoEKmToDql86QZEXJGm1QKOh2B9yb+1a9bVv97UM
yChpvJ/aDGjyc1MHTzKtiv+gmRK2Se1C92xDm72pLIVbjwaZ4ScuTH5xsVhKLwUW2R+2nt4kyYcv
/kIsv9pNjsK6eatWN4C/phY+kV1lzh3FV16bDeyKrWRfnR2hCUYzpbg7eMHic4Icf1DuxZfWtti9
i+98eXNU7mu9yq3vW8DFIF9P7B70jDk4OBqmFTAZIFe+UYq2TMQIRt3NUeG2AIvFugbgnw/Vbe7X
qLtTIEgjyEvgLvStVBN/t1Nj5odhgEJ1FfzjLgLzBMb+RaHjWv5rDlgl8+qOnNiwnPFBxzGgVam4
kQChvl4HFVf7JAblieVcL3L7xcVVMQBiP6QBuTks5gRNVFZDAhhWZtmpmzRtotVFOifF8piYTPsm
r2dJmoiJBJ1gy/k/6HcHdsGnnXexoMwTMJkgDmHDNdGoFUZ9WxsynsAz/EsyREA+lWXIkF+4sKSD
Gm+48riD16P8A9ICMO4YtqjDgUGAogywPZK/p8O+kuqFS+EzxPiegXc5QxHfhSUJHtTNQaG0ASFg
mWWFTyNeO2NNNcnSgYrRIH1+dKIBTeAevRe7CzT5iSlolRqxCqNz6/6g/5xpgDrHHUtTG06ox14e
6/0Z4EnxrOHQckBKVT+hOhBnemEMsP6o0U/73nfgkQrThbGPKBJW7n3kdl8T05nxSBS6sFPiD/P6
CE8MCxs1DahOXGPbBORoqnofbNY06If/0PyoP93+7BgBRaMYIgTt0ldk9rjOV6Ah0IN899o598mI
lHyPofz56pEZxd1Wj8eYWFhYaZjwEz+th1ncex4KYMZWdi0eElg5lPkmktROxkQjmrNj/cw3Gs8Z
0koxjzICADWkqvR5ICK3ohgtxaFFNc056qawRm7JdCMcJ5RAXOnh08Hry4HZX2n+REszrAsKl08D
dukAGFfNoahyp5NOx/tsAEt/9mt6uyTMcSbfVL2eBmcYDkbKjzaWpbJtmjOSBcw4Yoki6cRsZyoO
5ORN7GRQt8sC09wPTYnAuUbfYieUto10N9sznf3gIU5sxnjc/M/SSd6Y7xdHjK3em3GZZEGGtfU6
+4UzG08thQibfEox4Cdec3p5kT4nROP6GJLQdYPb28gtFuy3DMXWBJX2IBWGoGRZ+y1GuBLAcaKE
Dz5dvr16PxnK7SkyTdQLRxhUxLFDD+n/odcSlT2ii5D539wq8MFnWRdEy2xdljeIM6FUUEVNKmr7
MurDNzPCVDUpu+9eY9EMeEu2UARZtRDMpxwS6ZokcsQV9d4ZdGYzs7ncHvCYfmukQ8DoV6rD6RuP
fpzZY3n095XABYhnVBYmMECpc+8pwMpo9By4lKcasDs8vfygwF2IeFh22rA1zv2YfudTH+YbuviV
hBTioDnKiqO4+8YMZv+PBq61BsXrIwyto7xvrOWI4NvX7sj6B5oIJGf0qoAIbtNbgpkZwfrRkCDN
JMNys0B8d2tUCorfuGW/jurJMxsks3F4zXWryRH3j1mF8pRwoCV3kvlOk7SGCr8ZGT26jX4C7+lk
gU+2At2OILkZSO21TbldWWRjJgw00RS2oa9Lt9mQVpdQqZe6is8VWcAj62AmwfBx+ezsYj5xpImG
aO9OjpxPdKobvUB6Bt3eLmvbHYfbScm76CVG0IC/Y8jeJcUVRiR2sdHyDjTlIA53N4rJy/0OvnCY
M8DMHQbLfTTVxD7AZzq4cPbqRYD+O1V+5VpJYNmAAy2bMowlFVeZAXLYjkJ3HDJHUwCXCtBDIudi
GG1eAtkuxZf1Wd5U2pKqf5VsKXTL5qKx6oSJxtuY3AkIIB+xsMJjhu5+f+MlZSex0jPKuhf8+XLd
RYCgMAdsJaS4xq4ITY4Y1+aULmz8qwrx545Shd8A+P0omnsPKPJRrL0x0ScwU8hoGHZDd76sGiGi
W5mxwPEgPEDe40gJ8+lO3YyYQmBTenh6fAJiY42kSEAdlFTJ/WY7hvrFMROyPnmYoZU32opHA+YN
iT9gP2rWnzDX2Ge8rgxNBWu57zCJSedkcjFeHwDmDUgk4HbHpBKikOcWaxR6QYe7cVn80xibkaYP
+iraDwML4p9+QomduygYuEiquTnrKI/6zuxJjhkBipJtepmr1OoL05qVRRp/2wcRq5oCQ1oy7gOJ
NspWbsIUVDq9XSYSKHloDd1u56tGfcohnM40cTYDXZevwT9hyZ7tHzMxQfCrKK1/K21kJO4/tinu
32FbxsEkKhRV6XFZtEiItyVdUH8z3FNVqqZ7IlQPAIVEb4sdbVOMcMJgFnQeqEpgFYY7U8KF6pbB
bWM4IeOBARjbSZuzoq/QXd2q9t4tn34aQd4I+BOwwPFzJwDCRYAa9R+Zqt++ngz+sIDC2/TsucUb
VxresfpDDZRXqE/axWkBpQpmA7DB5wtQ2R5exqfZX1Euswl1+Ow9KUNjfw5MgScfSdjJBHH+tN4J
Lg7yzfDtvjwiFy0M1OggaL6ycgrRmpC/AunTo+f1O6qiPFtGJUcerWqHXI1IYfHNv3fLTfodeBeP
GMO0xNPF0Plfa7tUerF275XWoHaKer+eQt2pfPjQjtlpoaOCTuwlqBER7wveJYkOASs8EAJsTNhB
W2etih2TcFbMkOUkyTWsf5H3BZfgoRJZk8Sng0WfCz8Rh1TI9mswJLU3ajHKEVmpjQSjskzueuFr
9ZzjBF5dW6dD8F/u39fnlY0D89HxnJ384/jWX27olfw/AYD+kfo3jPBSHCncZMN6bydC1abD/QpW
JlifVSVhIlEiL37yo6KB4uyWe5ekhZc+N1zIrAFdyZXlxqMBJ5ngkCMZ2fO0rAdJg7TYmUYGaz7F
CoDYt1URXloQhWqup6Fl6fnZuX+WIPmbdepj6NSf8UZcTzB8mCoW5Spikh1FXE3pZQfxZPMtX3aI
+CapkoWvf9vgZ+7GyqIS5xczQyOWjE8lB0/fNRGG/faoceKmRlmgEDDsx9NXnrdKIx05kSHYN9MT
p3vUUGC0gsF5IbmZFzgEKWDfnnZhsarjthDvpqkzBGCbjnngj8QX8amoB0/LbgR5fXxlfZ1jcHl6
qWqdDgkAVa6uorKkuwI3BAqSF2mxh8OKsC80j0CEr6DFJDIi24Psw+wmzpDY1pWOnMVQjb+TvBzC
FmCDRLVqG1/3tCysehwKBWgWCL3Csbvd05QixlC90yXV5Y83skaeqWk50tRw1g+6sYZ74R7U6yDZ
iASrQu8B4lxmrNeFnlXrN4kliTuU8tEU5XH3xDCWDf5W8F6Ar7EZldtuZJab3ole+uDCc9uY4DHc
nz5Z+qe1ur3IEV0+ktFIn4dsUBoD1mWxu81bOJ/mVQHHuX5+OL0V72/YWdd7kbjW3jYwIq82aJqz
RF5KfoSMEAMkqcRxPyjQ8JkWJu8PKWxmCYkBtPJIcxrtIxesOWGu+PFBH3vznLOmhs+k/uzMPjI8
vwKW5v1NRWGaFNVcnEnAEx0153FWsZ1l7wZ33pueav2eLjieZ4MWOXsq6n3iTrCz2HtFeKkkzZtr
e3alxCFI0e1eUbH7pcb4a2oJ3tV8n6/k17eRI7I0TCRKDnz0zyOXjOs31hKIsgTKNEO1bsr8YNSK
WRojmQ4QHzKqMb2g5UGneRv8jW9o6NeBBqs2f7lMYAFJITlbGmHyqrnaukOApdESQDw0OqRfBVJR
W/sUSpUpjrV5fGnnmvsXwpBMwAzPCnFPRk55IARlCFXqMMlGnPECReIjKr4rG5FZvxb3LM+Kuwqo
Htr0ayx35qout2ThDME0vRmWBZLL1nkyXBaXfkZ+/3Mrx7d/vlJCcB+TjJ9dawmf5R9phbTUtIa9
sMqM4kDiqyhOm130I1vi2iDYqfdLFRNrGn7Y3QVoMftesTUKZWvGxdsSLrE4t/DMEfKnfkpT0Aba
EDbN5A58KyQwT3PbWA82nHOl3baTDUbBkoUyC40k472I5d6q4pAr9q5xJH3+Re+XGuqkKvMNR/8Y
PDiu9gZapVR5wHj6yrgFEFUtbZavjy5SEvlR/+7CrnC1eS6glMGyEuS5LmoJwbcF+db9nTNRGgaq
iGaw4aSeVf4ANx1ViSOmzVtEc6G+JtwEFGFXR7kZy/S8POJw29W9SM72lzyuhOUEDMDmsY32pljM
IBQnfpTtp2Ib/qj8fFm/GIVHkYXuARQD/CwTGr7rWqbioEmrouv7SuUahKmJ6dFp4Y/Z4KTjW034
fVwP2zHcauxePiIjxmqw2EgSOA6H9W7MwYhGwb6vM6ai4qza7mNnRvaS21V7QcEHSadr9LOII3Jo
St5QVftkem7WAmRpWrDhIQoHjAW/jPIUFBX41Eb58tIPPp/z5rByE1/i9D6ttq8Df3/AQbxZZhu/
KdM2Irhg9eOqQWPkhpJ7v4wQS5LUxCzCI+Z/zYru1Uw+j8GxrxlE3nn51II/XpOU92RJjHl8xrL6
47vWjhkTrRRV6aqpOO4DAU4roZZYSSK9JQ5sg5gTxg7DTbwlz3Pnp2vwxGr+TnAM8bnDOxZ3puf4
INYeY7uurXl/c51tMKuNymT+0b8lE8pzD0giuR3nh0KyNsWvXedcoJQ8rK32homN+T0Bn1OQlJFk
lElZACNz8YAspRJ7mC0KWIFcwl5ApGpXWvNkjPcXnoQsBDc/mP6FsGBSCh5EL36/1EPGV+4yiTTC
KOiPVGoHOwAYGzwFxI4vsGOhRbZfuG+1X9ZjX5mBhIfJgwhtig0eRCL95ve+P5Bo+8d3FO1FyqRM
o+DV63EesbSj6DsCLYSYonNw0LssNSDEsUay9qb590vNac7pZAsjv2Yy/lKzCANFn2VQO55lMtg8
y94Kvrs270FH0eOqkXZ6ysu3ppCmEX+BeyczwVR15eZwP4E8rteLALgKR6JIqQyAZAz4jrfeS1Dr
FeojkY2OyHm+pVZyyN0l1L52XDjaBTuZlEhtnKQpWOtjcCwCaj55O7gcKrSMz08GPCFyTz+lQYLo
fbbF0dIWbDWbIafSe63ZjBsbM1Sx9C1M1WSxZFdFGu4sbSrQgb7YDyNxL0tSrq2nOT6Er7uSDo+o
/49u74M0vx0IkTqgCXf7Wz0/wxmR5qmyWk/IhXCKUvUnPH2Q4+XitTpICNUlhfjWll4YkHw0m100
k+qiCkzzLKHA3lUtbZivyCJBhsqgoxSbJJiAbUW2hl8iw2ZYpBKlwB8rwBugA5N8nWLJKmPm1J26
IpqjofQux2Ub4ThhlAhWaTXnTW00YUJRTOkBd1DnmOgsuGQXB2rI/DKN5ORb34QMt9x/gV/C6XVr
ctEXNXeg/YSzUJuZPRLHVR04wQGRmAG8sdMGGDX6NRzlQIMUZ+2FFsaBpNARuWR3j5hqyMsSkrW0
gJlI/N8LaKxSXRc8d51rIy4OZbXLsM6nnJnWeijIL1/LaMHV5aZ85zjZ5tXv5eiu1N8VLqLgz6zm
C05vmNlAQD9YgFIYVU6J+TTBEvox8Ppa9ix0f8Dv185DPMQTbx2ATwrjbOeKMnonfpT63qXLvTsu
zpo0pnJjmLo+KGfqptJM5o3eP57cJWjOg6KjNN3T9sh6dlqB4ncPy5pvAVkIK3sUeirHse6DcPiy
dVTw/AooHftTtlEVDVOL7QNlzgbTzexeS5Ore15n/GcbXsmm6WzFQbuiDRxNzWqLntKCm0RRbXB9
HlhvvoEXmQ6MxUkzOv8N5aO7LrVWgDAqT2frBgxYK/iml16qmArfhDc2sNfHz3SCJ6Ya7fPg47o4
g+5KRK3FN2Mdy1SfCkf3zO40iHQvtBrS8iOrQ8ILqs1BL2rAw4ntBXf7w9GWHTP1S+FrkmLgky3g
8QK0qCdFheiUuEdGwy+e1ia1KjZHBo7VlPk3eJSW+LbFWp7FQ6U5wQ7j2ssKVVLC8es/U0fP62lm
bU4p+KxIpVg4kDEy63dK1mdZmTUYdICKE/jBtcz3ihugxa76YQz0DBbbR8PkstLuUgW/Ko7yGIAZ
uHECHoxbO5+hJb3FMnlg+cL14BugTXH0U6lkG8EQo06GfnwgDjwk7xhUKU1SHvUQpuKiQKqHJ1Ee
xpEPM6ragWuqo1MraC8w5rv8qu47Drql2NPt1hGHiIM+8G//Q9Q0oFe/wh03EXFCLLseLKSMLKPE
7fvgrCdqxFGDo4F0GBQ1NOJXsJc6nMlYTXHwp42zZEGpyLW5PwQORQ4VUmcKhAuxWSkTbwggzCJ8
bm9TQMJRHk5jGMbA8YFYwi9FeWAmqqsJ3vkQhzRt5cbPUXa/4IRuXQrO7U+QeN7XF2T3jRsILQSd
XiDor3ZlmlkzrS/u4mkx8KcsoQt/ZOrlDq6zCFH2kr5iTsnZuK1n1E2bZm3XJauYpt9AqUM6SQ/q
bL48ap56flfRsKt69oDFXXN0IONB74i9KK1RIGvUy5GALB8WJVbXFg50+V+jnps0IOnFf3b6+SuY
yi1izplinxl+KSNlalyBOcSOD4Nrss8WVIItIq6AmQDL0RKd5onJv1qITQviTlyNk/LkGcB8K89w
tJQL9Gh7HMLQiGqMjxDjNl59nZMHBKFqgBsAPslkr0md+f7K7fyOLmnc50CTsubD0MHbJfpaJ+rY
4c/DzihmAyIPDsfIzzCpHYwXgOvdgo+P04UuYhkFsC0floggeFCwCh5gyyFtGEaMaNDYZz6O/jeY
lXVZ33u0oIGRNunGgjp7EaB6FTCgnYqmIqKswyQcb5C4RD02UdUeahLQCNIuj/opo+2Z3Za9Wx92
J0ejc23qu0cqezW/4i6gl8nzY15D/Qt6EG5EuGW8OYMDOaIfHIxmS3YyrNocRdyrQUk4buJiesKs
U2EEZbY0yGhkwn35r5k6T3WxhGTG7d0exQGx6Ea4I+dB/pYn4L5PTdG8XbEZXOofOTXOFR+jFdn/
AN5GebtthG1/9MPsw+lSYn3SC4h2Qsfx0HyazGTVKZuyVdzX72WeKE/zPp2lvN9Su+rVMEJOpDg/
pEWPjXTHZx8z36vl2crEMoMBf7n3Qq2Q8ZPymznrrsHHgeyNBl4bEkMrHME79+XLV9qg0aUwN1r5
BLw+/kNyMK+xEtrs7nRFeIZWgLtuHct0PwLvWraVrDVqnfwT/BtIUdbCy5I8sfGHJUZht4qOqZEZ
Ldj2Bhf1XOQ28k36iAtqUZIVFubL3GSKv9e7GpvsxNK7Y9vs1bKhw34TpMrREkb7ye1UFCc4FkTN
Gl5BzN813QstITdunNp4CYal7d7wpZuvbUSLNS5N4i+GN2/2OsvA5Aaum/SBOXVTUjQ5qKGkaYUO
p8dep1RAVWlkL2eFYt6g8rTO65xG8VHdbMlL0JBrEh7KHewu37wdMMUG4w/BgT1FPDfTT6OdgnnP
ZGBkDEVPeXc5RY32Xr0VBM9OUxSfhSH4TKxFP399JpQYel8oMQAGJ4bO+/L4tpcJ8Z/JCQWyAdk6
+KZ9cWbrVdP0NjM128w5MLmV53a9RGSRPLTsdWIloWbyyXjPi24JUWH9ALjm2XokRMe+KDZxOi3O
5WNcQwrYrsIpQEuixqazp6Yf2Ul1R6Uu6V5kI0yULtOsmPJ9rhbFUxQVYS5HQD70N+4b6oXPW1VJ
DeMKLKWi0hJDfTUc6nsfqeGRlKb4WXKJVLZm0AFlWXJdfI3BegMYBsA36XwhfcClpyX4k6KuIMSu
0Y1ejtb0lfkntLTi0LCvLg7kBXRBm6GdOrhOdPrMGHNopf/MUGRFtAzOYBf9MTl+f+DtCaVAPEyc
ePfizYGFOyFtBob3h+MbzvPoo0qHUmD+b7PJHuKxrchvaDfrY8/Fl9O95a7z9rI4yESJTzz/X1h/
BODYt6JTVOxYS6AXSkR796IzK9KKCy1bmhOn18clJN0XReB3KZpmFyP42eLfo1VyaKpmQTYXQ8Tq
so3SM4jGKJlph+3gmI1YHcR3JjNpjvVVr8AvHRwZw3iTGN0bQpMG356B6ewgPhBddi3dbIdH+P/6
Kz70ImKGi1j8AagIBCHkVkmeNtJgt9wsm2DAfQVplk70NiqkRdk9Uoi+wxgNJNMmiAHqkcPrQ+0l
jXtFcwQmoCaWnSGaZxVYz/YXxLsPnKR0tjlrCDjbCLj7dTSyHWigX3323HRn4rbi39GiI+d4uDnG
u0jIqgsBkqIdOuiWoWf88u5k9Az2znVhhmmm30de8hQrLDeyoqC3Ef6for1Sw1s7SupJijehSsm4
YKqIZBZeR4Ua8/73IPM1TJlqgOeXXYjuXKnbksb1hiIgmDkJDe4j+T4zCV5yfLIn6xBTNHhXOmGB
vBHt7uOyQzq4y2tcI+iXFrwBWAcwFVWNlquguzcapAlfZKZ8HeQvGtstRdqgeRxOEa4gJwt2liVw
KuevNCp0Tv+ZTk2081KjBcpKmUV/wZEX2iJgF+LcV/lRyC8OXzOJaGjMURF1rct00XzHmdtW0kly
/Z2/9P5jZ/I+lPSTm6ss/wVZJ4KvgPJr7cfnYUcDHoLep2qsSPvmz7mPTSc3FjHXKGHcj3jVhL+K
aZpzeRcqQAOydTC5TUr0nNIcfppcVhn1L6ZATDh/gMxy9J6IfICkN6GfRioI60CSpCvpHXaAdXHy
VkuOFWzH2B++ti3UTAOLxxKPNNu81FLgLQoWdxXTpF539/0TdMaihqGL9Q5c6PaCHO1E+wry6eFG
pIIAL62nYdAr8+HMUQak8miCRC9xo87liRd6glQ/SLYKHUOIaP0TvYXndYaBL4BnS+hLuw90rI5G
f080gO3+aNnhXLHBkhuXP98UX6eNaxZQx7OMP4zD06FN3+kqyRF/0OjTWfVjmO3+jcBlq3gfckgg
qc5+KHwhzooExrT64+PNi9gymelue7rc1IeHXuY91jnCHwGOAapP5aWkMf1xfMHSOqG1NbUQm3b3
TlarB3qwDzEa8Syl1LylaFST4BCrWMruMFNFX34P/tR920lNqUnMiCwstwV2ab34LkCR9DqEG3xa
sEbBknCugjX4u0J7CvL/XyS9wdqbg3cWnxeq5y2uw8RFZVQbTtYBz2qwVBSjehN0gaE8Khg3RSCT
JE73aaLcn7LUJOr4TcqHC3Fi/FJi77QiJAKdB5CwAdlrI4Vh2/zPiG+atJs/xgUZc2KKdHqD0NtY
x3PANRzmdsWsM1pSNOwShSJyoTJGHWGel1JdwvZTICpl67mONos371A2znErs3uNvYBMF6ipGbt9
0sor2ceOKUa7Gq6foEAx0DCwnp7gEW5MccAbQodaHqQ2othq1UK7aj4CpwYx+zxqDGvUW1MOfguT
Bv9ViURUSqfLcostzI0F0rJ0lS2xXtiWzBvngZCYknoww2tLycOiifIGaI8sCjhUaMlMocdf/rH6
Xyt5aqNxOkotwkgoEIF9noHMBJyqhdGTM4GeMmY6z4kNzCIKQjXur/6fMrOOWCY9LXdXJQ8xU1LR
bwZ5HODheloTrMP1vfJCL/VWZhFrvcvgjkNJ8mbV4XYumctPwLr6h9Kl9HYH0Ezzmdqqey+vm78b
HaEZ/5+ViAP7K82LkYEkzMJAW6dB23mRlLlsZy3l0CdRga8GyuWFM0mqEZGfyoMpT/8ePRo5y+7y
YLMct4o6p95s8Gs3yEI2TtXR5AHphpFvUyKUD4wvSTOQiZ9pwCMgrOX8yagM18n7Uazh8mf3tRib
l+fjQyD+2tfQjanKnIeNAf0BPjeWlQq7QRSn5AV3MEtx9WqnJFRClOZ/Bk7dLE/+Mu0rTD5GlP+R
8cK5egIObeXhWLEQ51KQEFLUZ+rVGbowXFgvh3mOeT47cNQW9OhXvTEnGx9FEbApU71wV8V+x4Ro
dosdcZhdHA/JhAAH4M0tu0PUFPs/Af6fKP1oY1FSbwcYp5fDAKqHtjb+UZMy6Ysw4PwvUMsvljX0
rzVYDVsaPBS7/AYJi29FeUPLNvKDtIDmcVFm35Ic091VZth75yFs7wc1hw4VHVhDKoCj/1nQXKr2
5Uaw0srIWCvarx0QlaE2y6+ZnokiYsMk4sl5/MN85o66nXP57g5WAsc7g6azU71mTmY9Co+r2EOY
FhEQgqM2UvDTjmAbgeV59WUzVl/63ta1HUjsoOUlcKgTqOspUngDZnac3xQCFzCl+vyu7lA3Dqf2
cU9vcPhsp37n7gi5Q4Cz7kUqydptOSpCjiS5SryEOQW7/HupZADB9mPHBLQBP8TeEeUWw9ZDwOrf
E0AIPwy7YI+67MB5lYmEkgmT5JYn8EokZlEPp1HJuQiuI3iDm8FAjGbIWsmxTwo76qPU6PppcPOr
v5wHHxoouHVVAxcHdTwmgg7qoNQSbI0Y3N3+bFYKy9gYnwXMLZGdE2+HXRkiTjmgJ7hjDCSI6L4z
bT+wKaP0c4Gvz9iv1SXoPxDKOSYXztB8CVE1fo44ljYB/D4vNHDqX53KNDU6urUumlLk2B+5i3TV
2jc4sZYFcmSE4yzAht3TcCaSpfo+6TOrFcblT91h3bOn8c7tq1K1gWYfZjuCmJekuQiY070fDxJR
xI+4ac3/+GQoASKuEGeq6w4u3hFpxCt0d7ZwMAtCZHmnMxp5FFgvsOztV4+Y7hDKIDOCpCtMYh89
SumnFM4P8N32Ow92zIwynSi/z1Bmg5aOrhMwpmBknYcsuO7duq/+B9W/WnbHgOCSexcMGFKh1aNi
1ulSnD1BSfMs3d0euUUKarGoFt+ViL15avV7t+/g+NSvz22wnkWCmKAqepjhcwJhMg2jpyP2pBZT
ANgjaV9hW4PkT4OaGDqDSwhQE3A2rzBBYX/XmrlJCAtBsSKbCc7MdqARGXJ97T8Kd1aF4cxTJ8eT
Buw5zfl0kHz4wldGlFvs1CSZDeGUlZE/2GYtEg1INXZH44tYOXFlwjGqrcdgUzBO16Iatar9fLGF
AgrYZac6K433rBJLe4WTzeR2aokmgBDrUHtzXeGa25WA6eWpUC4+lySpcvqIWIxViqeRECm1A8nM
QPoLD1kDiMWXP9X37AtwVlcuGuCFhYf3qrCt1ceAsm+LHB8/cG8eQ9HWF/Rdrra8h/5QjAPXSlXM
2LsNYoL+oXIxnRGfNBz2OXLjaGgKSRt5ex1rCAdon4JtzLqDMs9oh1Dzh392wXM1Xl03URvdj12V
y/loUvX873AoOkJwqH6rsSR/O04kG1H6Nsu+c2YbIxI3E4a/sb4YjuC4U26Bqy/6w2FqNkS6nvk9
OXmN/pQsVm990GJnAIQ6FHTsOPzh50fCWDfrtAo1x6LktUUN57+A2jvwNgbbElvk5Q4so90ShTof
gwcg72joPzEmKm/WVPAT/8rHj1BTwlxbReY2r/KSNdSCe6/P9tI0bg90SaW6IyZTzsTtt+OSkUqZ
+/Xs5shWs/IG0DmqYK42D6Ucgw8+YEt5IDiMStcg/w48tcET5FNia2Crah2WzAL9h7mmnsiYHHw/
PNdrZoultG/8Uo2ujcTvGw2S+1BbMe4O+bSz0dNTfLhD5hxEo/ea2qnITMzumv+AsmLYTR8KiKsZ
E8C0XJmmrNluDFq36Uxq2yAH7xtBRY4mdaEjhZ7hyH8K0dMVS/zVRlpsTOiefl7gzkh9aQbOL/tX
okHgqcx4Zbu14/aKvsyBoAZWlu7hl3g1mQx+WyyX2jDyXdU+P5pGJJTxA4NO74muI0fteFNoMq11
wbKL6mycGdSslG2+Ss/pCDPyhj+tXldkcCsYru3QN4BzxYyWJrhjOOl/eyI16s99Se0ldah91zAI
jjxxB84+XMBpnoQA3vSYC9AsUkwmRkMWudwydhQ/GWB++D9tC6wdIySNwGTF2FQkSatXGdDQ7HRA
ZdapOpKCCqa/OEFAFJr5b7QgxDx5Kr+fbWo2M3LbeAJ3ZYJO7KESbC8PMWdWYo2/1vtxQDknNW02
VvBipoj6Bm3vTSZU0OAMgH+k0lPdPATFX5KEe9KmIchFAUuo3EZiTNQiWRH8VTunw96CQljfknZz
miB0kIgMSUVlSA10OlkxCzvQCrbay6KxNjM2Bj5y9sxS5tqX0A/noLQi+DeoGfw0JcSgwnNVcTDd
LZM/X5oZAnUr9i2/F4V+m5qGc6WYSQFu+FWpAPak/7ND8wDBog8+UoxvyUF6me3r1QjioU5BBbh/
vmP2qlPcP1o3ztO0jTS9pyxKFPQM+jEnG+Z6l5V8bXPe6Uez4kEWTVDVClVFL4pJX2gB98usa0TQ
Z6ESXSQkngqTriiScdnQPYOebKVbGm3/jJBDJigQ/dxvj0ionprLUpcF7XKifzw5yUcudXknL9V8
EAipzW5JX+XKLQlk588TmCJj0gW4AFpxY1u1KQlhL2hFtvg4eqrZj5HAw3ahsnHrxU9UzFRH3FWA
8cCKeyJ1wjkm26jT4659xgjfrtBxtTmSgxXxBVi+B4bLcgei4yAPpRpfzZL7rEJgLxvEyuUmpsfC
Rfmt4XRWKX1fQcFoQfakCcWSWPa6P/ojvh6sWcUvxjdLCEA7xw5TxX+eeFJTZ9Co2/UXi/2a+Q++
P5pnKLDcz23DUeEyg6yKoJ/7Bh/3ZdlxNtWWAMV76bauilso+AIQgqsbEhAvupe1DeHsu8FYpdc3
YcRuVUpSinNj74fcMcT2Ub02rA+AKnOQEXZIKw+HNhPWRvQC/8OE4UJOcpsSCOEPbA4UfMOp7n75
4UhPsQ4+c8dzErCDH50uH36qXS/J/K+t36hRt3KvkJGrR82Qc9mr7HXMODEAZkrJvWbt/f8b5xtb
V0wCzsvyTug7cdIpe2nisFQKoIS6Ds2nXNPk5sXKU++2nirMUuxwbOCog7U5zptL339vW8UhYe7t
Bo7+jFI9V3MoH6MRB+bv9cVoaSF7Etp7fhuJyqNMA+Vz84aNO3EB/sQVYu+86ZmkrNN1nWTPZD/k
cSHecXyI5OOpI0+SdPHNql/IpXD1ivKi0f/mne2/9HZkr5VMIrQjjpCM3ZUVqgzooJyN30IqOr/y
spQikW89wmX1kfEkpDmHC8vvumPK9dGtGHtgPsH2hz4hF/QQHqFnkxuNi4siNre4CT0jTi7Y6e/R
gVIZ2j9vXpl6G0ZchdmdMKDnxsYLEGwiAnOQl81z3LUtYY6nRiqpD2Lc3n3cGAOhUJzEQaOwORxj
EExqUEwLDoY3SSA57G/oRilMYdIzs1Hhc2g0HBrTdiVYJpBGJFlBW1552xgnzVHvbzxxEfOHF8BH
df0CZANpF6CFs2Txl8RLV+RZofULaqnI4WfvFy6W4UsrMSmsrjaZUxm9Nb1D5T3kzH3X0cUjKDJl
BUZMYqctlLDtdyiWlG65HWZFTntfQAI4PHHZB0L8oDkEKa88yhD7srwjrv/E6BkK2vk+q82wlbMI
qCmOukAkiPRBcRWKrG6wTSeUhHTEI3VBiR192fvDdz5mKxgrbDSyoOWruzg3MaGMLBD4NcnMyVv3
Eewx5GWatcV41nNcj/1M+n/zobeCfrQE3QTTDFLnGlbGiP6wNYCwFpTEqz07drHPD5xnRff4jL0I
Xvtf+aNMPQ6SWkza4hNmETFvUZ/PGKqzuIdAFZLE8fltVIA7Rhudpi2tgFoRszafRMq6MBYHOEbP
99efA73RW14Hh/RSaZS4wFGCjqErJ5fycxjO+fz7uubK/eJZwvHE1Yr7Mo3/HM2jOrJ/C+t8lbQZ
ypllc6jq6yZwU0fkWf6NWUzEgsZTg19+Sf5mDvZRPQB0mhAgUlClRhRd52SbNqmbeO315tIuOeo4
t9DSCA8uqrqFMH1APD+YE51AzXeFBRRT4J34pUAwXStyvGK45tsr5ylwYgELGZwIXsy5oWpH1M8F
dZC9EyS1SFKI+Knz7BxS763b80jvFFm6vdBKcDGILqpQN7lw/N4Yg7NFRv02y59EDuZdL5J7KWua
QK3HXz7ul9EQXdVToht0ugcV7JbwwjtcYvv0Ajxwca7TO/Be4bNrP91v9ojMd092vx8ZXcXHZ9OM
3DXTTIQZn7PALQGy3P5lkRqy/hQytaEKEw4hIuXtYyA/Gi0hdBg3T3F25u/c5monS20jV/pUi/yO
WA8IZPIgxEnRafFjmP6EPiflzEz7e4vhvEmRRu6cu2tvPIdL+0sJnlwLba+im5PPkxF25qE3tKKe
qeLkTFPbonIySXzMXLF8ar6mJ/arvORizCam/OeWsamROi6GSU3zg6JzgPffqZ7q9HNcuxifwRIu
m/87+l8WQrR4QAlVwKKkynzp7Mu57EbjPlefWVTAoaK3/GETAwQaalz2n7R8/kOm0fiS387hJAEZ
0HASEfYh7IGRc/2N52cL/0N0lWwDHXqP7D7r/Jh4l2qbVPZBNabM4R68N05PFJsnq5lReVk04jPG
Y/6aGvnpka5mJvYjdHcsn89Rig89bUt5VKzR1rjh1puJZ68R651pIbyppqKKZlHrOxmKgV/ZJzI8
puePBncPBCzPaAPUhy8bAVlb2sqF3v7yAf3YV5yH3B0slEL/Taa4wOGAvpr1p4vNrb4GpD4w2n5Y
MJN0TXLoYnbXw1V6gbPEz6doaFDlvW6CRsWWfTWXa7fzu7EW5p3qYJL3oJ2i8tb6IxzVjLvREG7X
o/QWLV+ark4LgkNco0VgcJvLctc3xlRttQOY2gzBrc5QC7wsFfsYdLzo3cwWjHXYvQzM23k4vtmA
p/65yocXNxQEU40hgxnZEApguvyiQtIyDkaun9EDkJMmhtxuGRO8UC6Vdfb37I41SAA0Q+f/WTmT
dTaXPHMJ3u/j72ACJsWQUr3DSY053JQeYP78sNDUc0G3JtzHLpy3rolpc05xlMPgm7UFrIxHNm6p
kDs2Dg9WVv6ccAQnZqHhb/CK7NZVMAb6cFMD2LSNAu3ADGHM6msTDu0duMXT5Sq6GASLPNgiIxQz
rT7TKtB6DWB3g0z+o/46LnnVZOTxtsbMJJnJrvUS2xJIySs/yzRB+qYsLXvg6+rx6jXTtEIRK3Tb
DWQdz/vF17FLlR9wVXvyipyG9ItKNifKNmRQiC1L/8TgCDXy9xkeyyCaJH5NnYOB7GguqMBJg+t+
ZUZcOJriStUP9JmCdchb1+i0rRk/JSamZ6cj+dh1ZBSh0v6Jn1cNMzwHAXeKioH0WUZhywP7/U0Y
wPsHpSp5o7/LlJF6FS0zAjnsU2cLSfalgaKEeSjTpHT0VGaVmxXueSaUspniuan5nCT7aT5U7KM8
+6Wl/+yiC+G7cMsKhk+twVFrGFJSMXb2XE6gD3XHinAU2bMo22bHj0WlLkXKVSX2SeXHG7OD/s+W
oK3sI5AuUDUBTKrJosBWD8FaPPlB8LE42GbZRgpqSRDRAWWoPvylWGJFBmbbP+yTTxgL3o/f9aYJ
PoHWZBczlR3iDcGNaDunlxIoetpP2K1t4309rLmpWqjNB3JOVMvCi3oihV8H0NYAZLAzGtR45bTo
VBVwRfNLOAUYdTth6YAPLv+aYQFrbTszNCPN0IqX7W4SIOAc1gxGN6igeN7hHTRLbATYR2KNS0Yb
FdnJelv0JZ5XXzsJDpx3hytNeSNq+KCN6EoPs0RmQ96GDUwQup9sH33E/bacmZceOaLuZV10HMuC
OEbIHspzIjSMmL5qh8u3JD7umPz9YJqhzLGGoY5f0D8+gzpRf63LzifR1j294YOXiUJAJvGE7hwW
OVNiktPzABi4fu+HqyK1s9GPkrGnY7EYuECvzYrij8uw/QYF4k7VxeOcO/AgMkd0uipc37Eufk3X
7Xlwzd0DFqTcTuH49Zd1j7zO90PijRJuSOkn2I5D74KSSbUQuULEs5R0QCJKeglBSQaPo50/V4tW
qqPufyLMG+C09B8uK95vskr2TH5LC/FuKJ0rczeVWssPcrjB8yvqoTBcH3Ec03ZeSXR7zkUbaVH4
Yngnq8ranqmhlVCKPbr9G7K2XEwymVzkCKhzztExlrMQKnckP/fqYgJaOWOvdguJZnH/SOwlKgKS
sbNwB4ILwUAQEqqmw8s/VT5f8ofqwAYU3l3JcwKMHTMeNRiSFtR6HJjr08iDQkH4GFARMgt6bAqF
GD1O6xIx6Jw3WPRUb1Ln2l9Nz7z3AyG47tkCFJkKBlqXhxK9P3D0biG9y7c2Bul55UtE+41hOIYu
8oWBP6AFUHP77/2F6PSEt4JT7i2nXSTfhGt6ab4U+gZbrKTO1gfPqFOxX0HLQ8snZm6q9bE+k01N
sv6rrzJqWVlaVneymXBK8n9G1jvbaVKK6DDdQnrnqJ/ff20rCUTz8q7zTuSLke2z7CfNbrOCq9f/
b9NFD9gqBWLFqwXgWxESZTxT7odAXaTLZU4SIQgS7wTJCa2o+AQPgyYU50bUS+V1bIj6rfa+lyZj
E2M5jpkyY3DXm0dmLSsDjHiGz59RVMHe8TNwtVss9pycnXpW7aJe2flLM3IGp3f0wRfiP/8SokNJ
ziA4BPceMxcZIzuIDx6145twPw9Pxlasa67fb5zcgnjVSSIBxq1qRsOT856ZCDUCipI8H0Ie4Tqj
dOf8F+w8pjq6uPIjR8i11DX+Sqr9Zvw+UTfJjx4Vy51v6lxWccF1GBJxkazGvzaFKzwv2Pz5fHTh
x96UbKk/iUIArjjNOMOOjWTi6wgMSrayrr2DL19Ki99UKTzGe2jhLC4kSNiAdtBiandL3eybPJ9e
Ipkh7+LxSQyJf9U0wN8cBbMPcTVArXQWjnDqGje3uRP/DV9vP5NX2vY/LyYDHYbciWtcKHSkLokL
+7fpfl6bKjd+2jjtcxLmCPrFhRwh9Fn/PZXHsZMix5FBMQwCs2s0I1NNAVBGuFMQgVGZjyCSdA11
RS93V/RQYz+z6MpeKAabEqxsosG8EaxvDXwfD0GdEDkL6GPdGMRr3+Ua/A8NxFYnwkG+let+B4e5
Fp16R1TRdMnDI3HgckAazt2cHpx6h9VsGSRZ+XIdRinF5zRcChoOE7RXXa0LN7aU3wm+NhOYtrX0
8vras/H++20rrvTxzS0X3+gdn+dGmjZfPiOoF6txpezNPXGp9SOfLSZ18BYxpR+o/3J4ozbNqHsi
Ll8TjM4+Z+8q6rsBkWHddHjkLQ0+N8SOYXP5hBXSsQlmgxguEZ9TkiNJJMJ5Jg7DVACIDNv7Nh5f
9diQ2hB3LTUaKKbcfaEefO0vQZQIn4atY0WixKsJoXoLEfX4vHHR6R2pET1qc9g4ggcR8rEfTgVJ
qBCXFQ27KJdddIlhWFoOuA+mP0JhG0pL2LuidVq7GogJP58YcEPBJi8JUnzw51Ix02U9TLBX9PuE
ye6j9tadwSrWGtCp4Va4oxY3XomS55Zmzpk38WTvSYdB+IIfg14wW99N4CVBixspgasND2CghAsf
TEVh2buMifa/fZg/MXqb8BsUWzCigwp1Ny5fKpEQ90xCqvBhtvqwnVo48qM/gH9rv8oyVZJtRWbi
46TqyL30qqn0pM4VbUIojvTRsq4oTmhB2cRpWM+74AhsX3oef3qo18nPep95UynEA1irHT/bYA+r
PAIkqucqlNo//FOY+Wks/FEZtH06dEi6vVFT/nfWlJKlYXCC9Y5bDwbDnFVB1oEs0B0YUlQSwbYr
gxqS59fraSZj19gOt9WDdcxAgMPDqtoZl5DS4b+c5SiABWxNRWGBpqkZM8wrx+j0RBm2hGvroqEh
PPKXkRX+A8czC1T+G8dWQSikSH8ISTlmYXKrXBkd2BMUOkMfHMEay//2Sy4uFC7cVh50FTEOf5PC
PtsyqBPZ3xdJCOwJmFV3AE6hBL4Hg7p1cpP56t7wCCWAjI3umM1JORYixANrkRW1wJ/sJZzEyhRe
kRCOJPWlZHxVtYhiIp8L0w7Fya4oaVxJyAvlk9pzab9JAFWfK1BCKe1QSm6Od8avMQJFGTx6Tqkg
UI/gQkaVv+fqs9EYT9Hp0IngUHHY4FzVeciHCA0vzkWfS0IZRZQEG0ssEirkCvZJukRmuEqend7o
dc8/1A5PEqcsAc3DsICjkuDy0GDKAgCuSKW686s2uhTdaq2g0kEZc14hO1xRXscM6BX5Cu3SxEdC
mAmYcvTO0SkmFH+GNioVHVBUsiKghzBTrBZJdjLlOYoTP0FLYrqXPA52FWBd979ruuDodmGet/1W
bgEkk/nLojZJlQNvak+vRb2hs0DwNhRAXH4nLkAGp+xSe1wR8peM/XLfkE77gC38LuWx0avjp9ZH
3KQ63Ctae3J7lAVlm8TmBXhQjpKYomn1PwSdyNDnqhZ7ufLLZVdMcsW1IbV0hLwu1z5Qx9L6tjB3
4wd+PIgeVyPU5yeJ1zwkMgu8O/i0YLEVITAQBY+4menHbDEe88g6FNSIgjqJuep2meumi1PR3ahf
zHcnibrqzMF4Y4xsQRn0czKOTavpZobLVa+rhHMDe+mo4AB2Iyu+uE9qgbNSXUmxQS8gL12Yahux
kxw224mDsT5qn1qXUsTddtvb6sVjxnCYZFSkqmPMWQ0CDKxHAsf78jPuxApmjJQ6OPIGYwdhXxBS
EVZggYItlXbfHnoNIHADJ0/83AIE/97DFFDFsZej1qERO9wghnby7wCFy4+5u3ZpP3zbS+EgcsNN
rzoVkUl8ibD4lkmcWSS7q3ZbZFPdHQ7rB2+AQdpCQ9g3NTmhx63Euv7Eqr3gunyQSJ5fyxk4j9d9
jZArjc5atzFLY5av3FxaKbQ8k7W1Pe6wmMahtFFFJdvF2IRsBqkznkQx665ymIuBgeSz4rc9k6nR
kw/1prKD81LHV6kXFS35jWJs7B2CSHKZXj/4VJa3ljyLS3OgU0MqamaIIzCXMluoRl2aG55EHSz3
YD+hQG05Or0sigPM0mQm0dPCmbpftSSSc/h4aOoBXb4PyUyvXqOKxfNVALxaP+CPPaZFY3mxABtN
86RhkzCPK6lmI4AfLC+WIx000R5+BlCH87nWlbLsTNZ8qyt+NFzw97jFHgnCxoY7LsD1yJmvIxHf
FThHDy5F7nvoZ4Nnhp+mqDeEKiXjJnQc47/6uwCp7PfaAKVxKRKLAoUksyoAa5cVPKLjCKoTs4El
IFL/aFY7h50Ka6v1l6oU4Ofjg0WBHsZlH8++5owjtUM3aEJgbObZZadL7sD6jVIWYRC6gisXOcd6
MhDbgcREfWZ2dNMd2YqPeOWjJ81vl4r4EpzgjPJu6CMKzWdCc0apHiyispXVVPAuUN1Q8G9GcG6f
82DO0NWfeMpKzvaiUXCTpanKLXPmO5SUvAMerNtRR+FCB7IdjNkvZ9ewvVH7OhHv6D3GYL5vZynP
0XJRYqEgNhGw+zFj6kLeddN6v7aJphlg0WgEou+oX8Acd9bS61hzHwrzCqq962yDRqNP5NTOrgiQ
tZnWy6VgHEa6pf8t8DjtoXviFrHUav6ty7C0yAtDnYzV3kew9nY8BygP//rTN84ybSHAHDSdI5Zd
XnARoCF8XZMFPo3FexnJt45z1YhKOe2xkzP1yDnfpKlo5eWHabC9oJ/cTga//Fag6PKLPF4y3wYx
6+rjQt3cbnbkQsf87Tn/+Ul03GFVVHOKBvLQiF56vjLWZXsYfFjWGi+UQeFWvIvW494LyNEkXrfw
DAFgc5uJj4aAlMzWQ5W8uzZse3bP/voOsvzLYx/ULB8cq4odoSv+oIDjp7AEAM6ZB++vdcuk6yaI
zdIDsB+OgfnNMhOZDTpuWTu20oo9FDjQhrVpv289dBvhLS/hgNr4ZLXmZJBRMrjRu1S78D3Ear5N
6KFlsU7gU3GbTl+LN5F7ynYr+B4SLuvqbwXhXLudrbwklYOhX3iJWoef9k71/7t2GSNYFkwNOB37
3Q8iW6sVzI/97/Z04ub4JstUVbxMXlCT1j/KrI+p3eMwfAbQfgceHdsFbuC2i6hbGzbDvB+vUDFg
Kmo87AAuKdjPKQi4/dTAoNS3QwMARp2mlgkZYBXLGWnYRrDWWCja7d/T3VKxMvQ0AIpuJEyYPw37
Bev+t/yxSci4QW3QqTkVl1hqdfrkI1x3HKIgWlGgqtO+rtk3xEo+2todrUUc0lN1hVtOTFCU2LaQ
yt9Rc6k0i40Qi6GjAmkd40WR75dce+NZ/8agLb+YlMC6jmUlOmIEQoidCZnAiS4LHit8GErlXBq9
4Gzegmhxc8sshBEzkfH4eHVWmzs00iHQHEVoZuQqGysmnuDdLnu5WrYouLyazDFEJ2n6mSkFdlhs
j8sqgRQdQrxX3ngLmD3wWdfkNj50CE6p1NCDkFXXlvdH1RIDhOqqGHXRvRqGP14HzpmBzwksLLmJ
u0TRaWIA7X3Raeh9ld1UxASFK/qZgE9e0i1Y/MuNsaOYZWDlnHjovhtHXOKurPn3ilfRV5DPSJ2J
CKDpvZRjMUXAO4Taye8kiSwEmK5b6j3InakXV2x6S+HPkGoBcwbTmFBcHssYjLKEEmi5kYNhKKF2
OiE4gv6T2oJcZNWBq8FtfftbmtWoW9chtB441U6gG/vd45PGhbojT2YTrLHhb4epO0u/GME44P7q
/3Z/QTv/CP3O1A133m7DkIrznJHWbAqIyI/exNm5HQCos0RDgjHqo1lnmq98e6jM06z/Mthmfl1A
f0k6QM34IYcd9qfN9YL1GiJp2WVvF4ZrS0kjs5JSoDFaA9uarQA7iPRWxPmE5rcvOmvu5o3J3luq
lKrYGikuGeF/Iz57+0to/MI/tfLet+HpuCOMhh62WtbN4p3VIpIgR/S3Gj5qFiN1bJxFxAmpD2Wq
mI7jEBbosIx1nyablAGO//0BCZ/ifKWsN0KxWChLH2F8eTXlXRJZypgWV60VHL9L/mxRASzQGurA
vqlxu0E4lms+BuASlZqK0LGzMdZJ3udL+0TehTqWvWgvOpIM/pGKfUCXQX2bCQ4NqZ4fyadlML05
flisYdkecLomFrUG3n41L/pEcT5X3v2SxwpDFXS8d50XhhInIzYvkky2aPTNHgWj2bTphdUVckNN
P8Kw4+9ijBTjP7F7CJCdA/2vp7mYPG96r2X9YGCxBIMRd6KR0W00K86t2el9odTSipXL4C/lAjME
rxgH2raA7j2ieDRW5tdUpAYlMz4uLNiLtN/uWAaTHdYuThZtXNdQmFd7drxjUmxV2VANWOXe+GvQ
dLG7fsivS3449mr+ZZOr7E73egmWTGn76XKlOXAI3jDSGz9WMySrXZt3kCEl01PIuuh7ewxcOKm6
9539iM9et7Ty/BDByZPSGWbrOa7nIJy8vQFSiBgiw70xAhpSyPoqiSIXcB2ZELjUOI8fQ8XvQ7U6
F2UN7crulNj9o9tKz4e/nVXlKKKnaQO1l8NndA7Ud1osSOYb3hDRYDz9Vhqzv7yIvZ5G/oYaSK2Q
5+9CqzUiXydQdQ5mltPYlGdt7gMAgBqe+sWGTVbVsppH7WU9d4FwVrMZS7cO+doyuKOTPulQC9sh
RzRcGa/8VxsYHXRpc94znuzPYJDq8mKwN4IKcrhFmmVBEOeJkKWLTu0ftCiC42MAlqt1QeMTgq0e
uCaELHjfUMX40WXy3sbjz4om/0cusvLRrGBA00P+w0PfQK1IFY8Y/ALYiTadDS/wNMSlsgZiKiZB
2VqKmxiQtpajtxW2rJ+ogmASHeVuoCcr8yvgZZFwRKtSe6irQjk4NHkiF+EsqbwdTpSHTShyiPNn
UIxQw6Td+POi6E5eZewO4N53VBWMbiNByA+RKCA53GQuN4YygwoRBgTzgGpPeOsgbv1utTRjwT99
wP1tmA56hzHhTDpuk+JKUaG+q8rJ0mnUZ02XVJAq9JIYisPn78TkwSTBGEq4nt1RSmaib/tt0fgU
7AJm8kC0A/9O3ZNmcQdcrSVJo9CR3FrjKe6stOthCRnTfeA5q4+skgH52A/tT5WLKyE4HmZbyt7O
Kc/cFqQ/F5y98tRPRvFThay1rcNIfFUm/ZVfOIWveFwe439yhhOFYfo1roaH3t1mMp0tzRGEof/y
67sdHUEW6o5lbauvDG4owgY8Tp0QgZ67wH8krbUbK0wH1gDjB8RpG8U/HZtMQZAiydtbjsz4uScZ
UuodOpZeAtUYffFQ9R9oyoAL/66uOAKXgaA6ifLTWVNKjGLi47FsCGsunZzBoW2e96aEuUIIXnxk
7jpGVFVn9oGm11Us5JZq4XxXdX5PK3+xo8o0NV63SNn//kS7KwPeEQffA/AF3cm2N6Dhmit3WC3t
vMglb4xdae0cpocD0XeiNBMd3XXDR17JkJ06aXLo1K0E5x8U9wx4qyNnRurqppLpj2AeWWFTur9N
iR7dlcibSXWqhf+vBa6o1Nr0RoHEJF+aODOttemKspX3XoArhTp8uDg0yS3oa2tzWR7a5xe2j+fs
4MkZjH9io2WYJ1Sc9ZBy7wcpo+Vle78YnVmLF3kK4gpoil9Fdv0a1eZPV8mk6IDkn0pjUU4HzyhR
y0KRUJoq25dF9Zt5ytKd0mdzLqkbfDvk4Wav/P4cgNcj2Vp5Stxl2ZcR6zR3OCOjwhhGD6PiNnlT
78CTyz+VBa3sqfo/ydWvwCL1jeXLBFRWCZ+1Een1AghepQchqIriNyfi1wEfN49XQ1hb72PnbOsq
kJ1VdQNIPGQ6/PJgKmx6tnrKr5MLtseTjn8NZaP9dXPUD2GXDr8qnptqeMQM+X1As26V5nWP9wTo
I5MDUHaJvZ9yEyoCDLjD23b1iGlUhB6INXzZNDre0x0MCLXV6nAIfk5BiF+AjlLUuOZbRjW+g1OB
c/pz95B3Dqh69msGhi09fSTRUKi1AuQLXUzQzUJAv3BYJ6Ynji1fmCFvNIfXOuCfnF2VE4BHf7sH
j0pGX36ZnF4nTJncu+mFzT+Ej06PL+BDxwXDkzD1Wwg3TGD+k110RwZ2yk/iiXKi6jyla+SJ+u4Y
pq0WMjvEAZyGqG2NWqS2fbUBJzVSeZLcgeg68/S6nn+GzRzzcE4y0B+rJTaCWFk1HFlRw5r85/uv
i2QZgcRDWADNmOHgWLvd76IsZQWj8lGo/TVD0t9G+T4Soxm8LEjZrogFcmUsCYSWWoRZbMh35edo
DXJYp1RF+HlgvqRTKR97VPzvBMPQFpQKvSXr4+zcPMx+iLgnvNrODhrODoIAL7itOtowU+mtkPZX
aqDCLQLGh0Ox6UcVdYjCVDkd90NDiaM+AEnBOd442XBVxo9+NOz6qzHmaf8UYSTuTer9JE8KjaEA
Nair58NPHtZ1g6fPvNQjoBuCWXvDws5mwNYhyPNu1TzMtkI6vnqr+O6KgcjTXngROffD3fpPzVch
RIGtMcHeFcnhE/WbHbNQZehPIYwXA9r9aeuLt3VVHtaVJ7TPlcPRVL3Ly3u1DmgHLW6stQbNqwgc
RR2aVLBSPHWtu556dd0jMU2h0/cTP9Hm+pcKS+xTHwd1nX4x7jnlnf+Ddw4ZQc1QoaXHHYkqq4rG
jTlTv1GcZMeI1VPlflkqsn3C/M4upSFXfyG5Whh5LzbTZARzQAJWT7rc4cwOw7wOxJWRX5w+YGA+
fdHw3mvsVz641M40wIMHp0egu1WUUwa9LW2Qj8/YmaEh/aWa+1KWDfkucqIhPnGXeScBiuA4uAAs
iQwnDGv/tmwNxhVRNLUZtju1EZxESV1q7X8OXY+LFSlDuta79XZkSQ3No/ioW5QRTZguQqLtqCi5
GJPgcKvo2f9ga//6/injzWUGhmovu2QdeHVGkCr5RlBAbS4De7WcF24yZpN9m/4WmVsn8MHhhTso
NbBUiOOrjPYDB1dNPfBg8ZDgCIqQ1ZVVxWNAmkbZ7UhTR5MpNAbfvzgerjGDHoMLyFg+KUnQ7BaS
uzGXVxqy3aLz6mozFt4Rzp6F8qejES2C9av6Kc0T8mv5Ua330/dwAkSKX56MmQDsf9G63g8dkROE
0V6kK9yFvvseO5ZbjioQMwG6R6xfpzcVeq/bKrvQwvB8jT+yNVkrMsiVDay8BDFum0t5xX45FxaX
TNMhgR09mchUk9a0D5/jONOAPZCciBTWv/DyocRE7Wx5X4xRPJLNOXH9wpHLhezk+evKjh22nyjS
DtQU5zrf1esX7tmhB+nopPZmYJsItU3NqyOnkE0yAFwhbpIHNVugo8+AboWlU5tT6Ex5F18zXT0a
sHiwqvFeTurDa5D0NKvrnTvXL1VxzTefRdG9eQArm2GRBgmSSwyo8kkefJyuesiWSsusiyyaA6m/
YFOhggX2A/L3b4o+JamVsH1yTY4/Ek3kcMjhXgbfVVYj0kNrrYDsGquRvTI1eGAAL1Ds/UnT5FWV
XWiBJvTjo3ywu1/T6iAU4u3A8bvPNZ79t6JuAP49Em6GzEQDcpL0f3Zv4ztEfDycsL0OVTqciU+B
Qs3l0a12aiGtFG8AdP6P3o+ok8IXkdxDhl+fXSqD0w8igNdQbCjh//AouCWuBWlegL+K7aAbPTuq
7HiirCt137n9tomsbheAjMiw7JW6XnLo9OR1jzFRbkQubiwj4v+WDmFDV7oudROAMIV3rkgdxln/
Oqdg7wSY+mTpAJHAjn2faIGXmTVjyo0owycHajpxIrvJFdt5WVFasVVfaMz3MijNY8PQOQGtQptj
reE3xhYnqhLH0vwhrC0gU0jnzCPBk1gSCKvZ6aR1LArFyl1LPZhUBxydzXMm55ZlAsX6Wq+t3+IM
vCVbywrDjASsGH76h084GoWA84Iuvk/XGUUhPOvDA6L2UNw6tOdFR1GqRbocrLIJjMapK9M4e+oU
k6eYHe3GWQt9TaEZO0OZ2uHVXW2VXRPm/0Jo/4bjGOFIMDenOUUgYokwz5iboWapT/UkRLz6CVjD
dqWzPhieorHXEbolmN5W1XIubCSzhhIWHcTRfhZf/7qV3Wt6Dtu1K9Faw5DAMAUul+Bo6mYMs0m5
G/L1QAz9b3RfqUpgKAXRyMwdzH3OQJ9B89zbUxv4hL+I/vQyrL3E4mhuD1oILRYRMgJfRq28ELUN
gBRjNFNRwlfa4NJmst1CxEOEX59hw1XPA0IVfVIFtZP0W41nLu3Kbqua/dzSfZhNAeaUOINvFnc0
TDa/6rgxHM1Y1yJ+Q3WiNyXVn2OhkHgMTSUJlPxTaamDZqyHdFnLi9ok4yBRykcwobqvZqQ7O0ws
oTwEEky9EX70/OJB0+xsXpPApeYigOmuLdwwAsiOG0OzuQACl3bec4wGEA7Bcnwj2QeIyDlZZ/20
V29DitLjbIKU7651VpZL8TBaTzGGWtRvYWzHr10rwJfmRi19D1fkSuaizDo+HNyf58CY4J/DBOjZ
/IXD2sB9hys5XWgBpT842hj/rYTuRk10sO6UJqjL7+frLN5fVAzOmRXNm4Nmk5s6eYTpmrOHNgrm
BjUomJH7+TZ4Wmspb3dOM0+HDDoVFFouTYBW/nyBNE83aHkInu1JozEqriv6zXwwfMUeCHAosHr5
rOh0JG1d3pzWVulHjh8nVA8yR9uVG1MoiXGk8EHDSCPE5WWv8A6ndoqkaFatx9yTBCc0j6/IlY44
OUci+Yd7FTJ2W5F0D+fYat14jxF49poLJ4i0ePUvlGjHUZ2nAvdlWOZVY+TB0/lCYkQsiQi0phbk
W9ZdOxPTEyU0l9a5iXH8yhmItaLAt/MoActNDMio9LJmgFMjXkgebJWDru7EeMm/LtVgFKadM+0S
PDA0BnrsEewYasV4PBDy5wduPNt32ztkeaGKUKjwGXCaC9BmCP/7IarqMBpLGvLSInhZzdQMOao8
yOexNP+7VhideowkfOqmdHw9M8YPCDOwGoK933f5nGYxyygkBwudXfHiyK3rxj+vnad52ytj4TZR
GXySqjp83HaHo8lhzTZh0eUtfq5DBsD3iwOMVQsvZuWinMmRRh9aS9qC7vfmJDPYMNsNOqAYRCA0
PWX+APT49XZOUL7bHSN5T4JYDcjWYtGTxcx9yQDPigjN2qSwPf27AY4WpMfrLIsMw1SZ1moXM1cE
ymzjj60A7kiwujxv0EbOp/fmk2a+xEFxPBqJNVruMpCAY7231ayO8tfm7OuBchZHNP+Frm2Hc/xs
zXkD+UUThsEOhYZZLN5WRf36Fv+is/MJmQgdC7iK2bsNVn+AteFDk7zh6u1c9SX7ETXzyaCCRWWa
COl8iJGy3ECNY2qqiUBwu+IQqgiqq4ZLXUPvNLw+T9WTMB91l42UFOhDHC+/qydJQgX25u/oRtni
xzy+zXrXjAGFQ8Kf2aEmlnSeAgrET2uBlsyt42v46+eUBZVLrEIvOZI+hwvwxI5j4VGkYiK1zOBq
eDwK5nTNa3oC51OkCHxSwI2DqsET5UctodZx2p3/1CnzkmEMCKa9e8X+RR8VsuujdKMDgNxHTxdT
cQxzV4QDFhXQCRtGpC/3e2uO//cRAp8SEXn/pW8X/u+HgQSmWXXBc18Pcf1QFTXzq/hCs3rdbNGT
fmRYmGNEyG3jzGtw+NNehcsspGm1tVdNqk+2yVt0f52AJ+ACGkYEBoS0mH7L+EaD6nYD0EWmIdYu
1o6Wr6CeQmzQN7642FH3d6XWVF5MT8lGdSNQG88NrjTeXDo3Q6L92NIbZktpeZ776uw0j6Eq+Mkf
D92tuNyvTFigbz6kDogt87hv6MgKIhZstYY/1juDVFVkPlEGkO6OIIGJc0KZ+r1a14mON5lghBTv
2zN2sszCwvGv/i0XlcWPq2wFpowatY+mAq7q/M05yzZ2XWUVXtbOVbuqhDuJPCcHFms3KWHizR3X
H0MGQkWTTZ4ijMdmiaTFG5usoyHdbsBcdQVlJG1nuSj1lTL6fFtOO5bXeB7VR/2nHQecP1NJbcv3
if9JUAChuOVSaPc6rzKXS8YRRWi7NBEWpxD+tOnpchZ6OPKd1e2pBWmMkd6d409i2G+jmsQhMHOb
5l+5uuZqQ8QrGIOg6zCVWYejauo6+Maq3NNzUbHd4INXfBX54dxml6mZmiccJDG9uhvCeG63LvYu
fmVkiMT5OEGj+b8yTH5OMMCUfJKnZcetzV7KsX4D7rtE0OEGaH5W8fOyd/hDsb6S35JjhKTv9NXY
cdDTA7A14vH3+DxC9sAp7Gw7nZcvxQooy4DhFL8OsbSAemQeiNy8cH1gNkQ+GGgOh7zP6wBUR0xz
dEoVXkE1klBa7MqmrxVERbdlFMwbH3yibV9d7Y8dc4U+T4NEmQl0l6Y+fTW39VpdHBVtJpa95Twt
rvmPwKZe/wYOZUd/Jx9OrFFHzoQHQK6EqltUwtammKe1y3yLDC4wSP9rl4GzsED+u8ZJZI7HpDEU
f+uIcJozpJRmwh9iGPXYVKqUww0rWlSJRkb4Qx7fnYbZKGmuBIlV5+pzLVuHRf/1KgZQAQ1/zvpC
s4DyzryJrR60f8Ga6++VVdhoQpNrCaTQTzECXwuftuVcuIpjaW65GdAHm4xtzpzBXiQV1fx0Rl0B
m6k40KQeNuaPmlyvbMwK3HLUSr9gG8G/Zm7YJot+Tu9SrKPJQhQd04Q28pwWimzh10bUr04NLz8T
hvYLGD7nA+Y1BdBv2itzvlPNDll+hnDdV5x91fOszvL96SyThGNJthsEVmc/BuGlh15TN76Tk/Ze
2eeAwOUVKU7YIzF2YE0a0cOJ2PMbTfyXzBuUJ+9daeB0L3rcePpkqbHTEkS0h+ACA7vkj8G0v5B9
fmQtbaySS7JFX9ORJniUqbHz8iw9jk8BBa03lapNbtR5QQy9M1Zkj2vWQc9KqCOtq+R4LKJIHhTh
bn0GGvTS5IMHqgrfBeX/ZICEYmZ1GeWRJrAeXFbReG+yoWoKvP5ZxBwBDTxGV+vv1mIO6L4WgnQN
ocwYetv8EHAVu0kl5SI3HZgyPdGJibp+TFIk7My9Kt1YukaPM/ODQRpmOXhlUdFBo+U41TzRm4Zc
y+Cl1CunnC9N6KwT8i+53Wu8AWTnjsaPfv1tqnbq0ZZfP2mBSdDNbW90dJPTNKVrL3JgqEuavLEs
unmfoe7H6rO2pvkcHcoHWzL+SHIKrIZH/SbNyZ8ZbDrp9z6FDOAYC8cwLR1qQ6AN8Zc9JNth9RKl
yFa9f/3bWKXALrhMHODXUTriH4lMnRQ41mNLqua91DzRqZg8lFaBKyVOUKY+5upgst9lHK04l0Na
mkayNr2+Y49db7/GuqA7sciqK7XavjigErNGaEQfxPh8Cz/xKUrF4FajSLavUcK3l/eDblWHm9Dc
KAoeOzDg19Kgyv4cKrwecBwoSBwYmKxM/qupE+TZDCeJuuZNG1keLMS2OXGe+Vx84US/uDPvtXTF
Ns5P72/MSI000DjY5D7xenr1LAenVNvSOeCrzubHmZ3Bk11EL7ES0pkIzL5gQVVZQkGiyTlxGGtK
Rd9DQraNLIM4CIzNoru+25SQIFwK2H+YXTywpRx3eUCZ7ycZDpMMxjRgAbDQiDyELKDGBnB6J217
RC/hNPwACb9BsssTJOIZI6JrDjH75Mj6/BNNK9O9o3AIxrBNbUhUZkJsYIar9q6LlYBVsNYDgS8+
CllYqGkEOz9LiDCKJeRD0swBQLD8d12U6Q3+RWNxU6r28WKONm47VRdDDa/7aaBG/DBmFZGSq//u
eb6Za4nTZQsK0Krr0rlxY87tH7Q8NS1l/kgZKaaq705N8qvnbwDLQMW2Pa6zavM87JTuPZxsRWgy
ipfEytAuYYJfCVQJy215oJsQdq01RAG3wEJzzuLS6sAMNyH47gwY1Iskj5ewBX6GdEb9q0/Eraip
eFUwUboHhF/81w3Hnn9dCwLCwkOPSgZqcMD6i6zHraLyAUMl9E5fIIcc/twbVky3OvHe7xLstunK
J6OuKLpYTbUHhRO/A/QmQoNKmRLauuOPIXVQIVotnK7dqrEEu9cLdQaTTSvhUsXPR4E8iUPZULhX
GDPSWAPOX+v9bR2LICk5IhC/FA7BdV/rZiXqiX52pJniE9V6ZGD5UdxhYOmFxSf0QT3Umx2Y/YgB
hsiVXpo6IZppRFkNhkswG7yB+NK/yDQw+LAhBWF1+ZqadjCUg25EfOHDmMMYzY/TAQ/NqwJrd0Pd
t/AD/NmGk6pznxskvsqShPIUB7wKixGJxzf1si12OBIBqDYHbY46pm3rdbcVyaLJhayqmjDzC5yO
MShgQmYddsNoXJELSDtT2SJCOWkYBk5adcPADOqd2CuR93VybQ8zUsnauTfDS9ypi7/NBHjO4cEw
Sum/lwtDo8jdBtIcD4p8YuCfXbY27A4dBITXQm0/S1jCtVrQnomJu3pe4MNL7y0AThCPj0FSXLNw
gaVc2YyBw1nhKMWM88tinr/9SxRCMOCULXEbTJ7HuFX+cHunnTji7X2JbVDK0U1N5RoEYlZNMqmQ
JeJt1MffUfqXm/t53m3660jjwQZfm1rtrUXqEoYajfTe5nWoRZi0kWBtZcGP2EHHQNO04ZxaZQml
PPX0ayTOjAbgsMAQKfM+qM2vt7m7KdiP+jn+4WFXbgwXC6p5hYUBf7F4LP5T/x4mf2VDu6+8dFcL
3kOVMdF6yMeXc2tTcyP+c6IwQwm90mErCqxknMlwvbe/dRnANJVaJyPvkQQVXr49cyt8WePXXP8F
bVXtLAkDMX/L9vmNUnGf7O3aA1qdRIdQsUNDRtsn56z6diyunr3Zo+qr3e+YUX+xuByXw7nkOsy2
OE7ERVgWa60L6kSUmnDOLJPl4E5pyqb+XwZ/7Sm+LsdIqcvnmRdQub7Eb4Oy8pH87z8TAOSVQW9T
h+BAGSKmGarkyHV5IfpaG/yJL0amsSOFL+4HX6221Aydv2oEO0AwGjB2btELO/2WQ0cA/HWd/dEs
3PsvDFkfAfq4HU2F7BICxMobd4A5fxIK3C57TIMzr0xhFL6Qy+B2gsz23CM0xxXbAeenq3yLJlWp
RPEm55qTRU+OxJ1xgc2qWVlytTO9HKCxkbSqrgletDEUAFw/9sEZFRovH9nqZFojKktmozW2bTZA
hfxCRQ46kcl0u9Hg5tXBSNGhl/MR7Dk0FDMsMVw7bMTqCOspi1Ke1DobMOr6n82/he9Z+JOJT0aE
L3GrL0fXZywq7lqeVlzrZdCzy4TuZ1q04W6ylXpjDpMdRo8Cl23RPaZhcakQtm9e3m3MH8YVrQ07
hT6py4LWEkmlVc5f6QAiO3CFO/x8Ryg2Eq90CmAflebY3eGx3ay/Y0jQGUnWh9pJQXKSGxg3g/IA
JleXNvVHMAvVCqm9FXxncGqDjDuY7b1BGYSAU/tAQhEtMl938iHZa2qkFR3T2JhmqYRtzFOw75rC
0LbTT1S1zVc9vcuQvta65QjBpwpRYa+4e0Xo2QgixlIFmWZWP4rYjm7JEfpDTww1P0Rtz721cHqV
QL/Tvt0qNg+XoG2gxpmL2GrpTofDHoyKYskfeUQioGWpBeUXHv1IGawPpqyXcAttm8kD+yIiB6Ju
rjIBwvnXK/4HYMBNQfPlOUpbh3NWBPJpZGLFRI/uc2PAj5iNYbsSGN338xA9vRHKn1e3Pbvqin6D
kjBdnHjEzBF0nCjAn2hjbj3CXlw2dnwIJBdJBrz4Bmv0/PTNHrzL33vY+tMCrKYfPr0i+ZKD6qrz
qsTG6cav91Xe1ZKH0iDcJxe/R0YsJJ+i4rpsZ5Dh5wgZra/kEGbkeLmOWvGkcV2xRmp1QJdkUhni
teBVaqIKS+8+uVF1caUyLNeu9hK66XkSGfWOm+TwxnLtqyIUgHX25UTvFdiMkt+u1ce3Kr44tKB/
ZHQIgmht+TWcPiNm9JBJEGh5u8oUxG2wGN+GCXELxtuW0ZgJ9ID363eZHusghushx+GtYjv6m2TH
tFkpWBuBrATpCVjMLHDVSPECnxDmd12hhqwjuoQMc7FVa6TisVlu1d3fzceN0RyxCAgi0oseDHXM
xyaiM064PSGUEBgJvEUy5yCsTLml32OTMQaCr760iP3T4VWtKb5C8c8gfeSEyy1NGsoQHk0ZrwOK
F9RsP4bObOScW9hCjXPpN1vxS7E/zVM7AVdhWsaGTV4fOmlSb7T5MgR0+/NX4UpIt4XXk/hULyH4
y6eWayhJ0dviW4wQ06G8pLSk87gH2XDqE7iUpDMBuhKbplgvG9F0NpEfrxk66ByiPGe49i9OYx29
7jYBMi6BjE7stVHZlIZCrmp+Lw9w/dZKuyj0mGnxubEAS2kNwUcqyvi++8lOHur87RTPfOu/jPHi
Occr22+OUhAD4PYkOZqXVfqDF7lKxU3fV9yYXOfslZMeB3daH4vbkOKxeLjKq6zxugHZYmd+UUb/
IIXwmxn9+m93cIAjCQWMy9hw/zTSYqsqazMehEhw37rZCEUib/0HmwiZCkb+QwV6nq0sHNuPHCKe
AAHqJ9CYKlL5pBRvjIwyQTfySdo1tQ1uKS0DhoCbi2I70JCbJ+4WxAIIDgeZRHLVnyAL01UAF9G2
JZeKclVtR3RAkHQALp9tXzQhvOPGIcfFHFryD9zcfAy31hahlQ77I7/93biZ9Scv4tAn8Y6w6FF0
5K2MyMlEUZ5Fk13DtvvA+9kp4tQorAypwmEX1Zod9iQ82dTuWJ9hM4Wwer+WDSWTwDyK8C4Ftq+n
S1H301I5V0/hiiysrB6dCNUh/ao5AXwyG6YwSNrvmJV8zBrenZfVN9k/N7vN6a417YXg6A4LnYSO
39OX4uTHEPD/fpNL96YjW/DiALXaPtJvvuHnqTrIJxwSoaIEmMcjegEp3RuhYqKdBOONLQbSvAmC
qU94TQ/vspZVsRvNSfAftif4XsqEsRmZNokcbZZWhv06nC5ZlqLw9QTcXL5pfjrRnsPqDIQsZme6
r3yOobiXVsWd0DxFVU6Dx/3e6OKWYjZ9y7xGkr2pJhaBmNz57TS74KP4m2YtcU/gnH2RYry+ZBe2
BtbnFjxLQXderD1kuDQIoWIoStqfa52H7wDbjeYpwo4+MsaTUKxfO9plN1xxjd41+y6RXutvnz3L
0xMjRknSOTRc6Lz8apI28sX16ckz1qvj1fAuOFs252sj++Z+vwA0VkuNjGVOya6FjI0yEX9yf/nX
dYDbhuSUGo2VkFN/u6pyLufaXs5YOFUA2QMIs9JLxjqedbaA1hr9s2Z/YGGWUap3ndR6MRLqlIcY
WMt3p0dRVmlbkl7MFkXrPBiHllyM/3Lu8NckNN/G8erOf3FGMSJD6Uunx61NJPuczRCKt9zVqk/N
cNGp7Eo//fsb+iqLufxGbOHqYQcq6fmzWjyjpOrcNW+NhpIsBq2IHiFI2bw/NtJBLWqW3zPbtqf0
LQBG10PrBCvvu0OIDjODl1z8Pej4rAGkuT/WAhq7Pj0A6CG7Lhk0A/PP9ZOPIWNKKjCw34tkrhsM
zyNg2BpTucCcCM9cDrZHuB2aexj1ziMTkQipJ/Ez8cpeJXuG5uFJZ1aUcy63ZSxJ6QdjVwU3Ihmt
VC0KwloQWj0w2Am+oew0wwqF08QRgHG5EgU/6RBTkZpHUaixCGA8YNbT8TfHn4c3O2hXjbkKfagS
8WaLNLsUPrJmR18Z8AthNQ7jQ5GPTv02NoATvxZoXwQPVy+iaQ5XbQdo1E5DWjY7Hm92gbBKxwnm
/l0UGLJ3v613DFAPy9XQ8RJ5SEoZLwQXxGfOF559tauZpA1Ls/yOpo7SKdstmKJVMVrnNF8axIpP
9RoPQJpwhz5msiDWi3gwoGpE9ZW8F1RaEN0oH1kUeVhPjhzMkXKRPNX+/nmqArG5A9NPj0Gh7RC1
uyGd71HrmHoLWf5z1YngVBp3Rqcjpq1/Yg/zFH8dDerOpE5mZk7bP4eqerINgqC5WwTxu00MnWRO
wKj1uyCCi2a4Exu72TY5g/lnpKP5S2rX78BSdXygsbaEJCAJnIwTWK3KdOXU8vk6kSTIXJZTuoxo
bZ8NoZfw2XBPfkp7VOMRrNyTc62prljAJz3Hy1mh4A1lkf1kqB/pMBuEG4M6CbiKPHNtwcX5XTLc
VHPbP/++aJszXmzqJdubSxWmCYvpsiUsuYr5LwCt1y4fiFS5ObcIKbyx6L7vycj9J97/mH0sz1L6
iFGUH22giF3hqdzApGCp1pYlQZmUnCG35OsRpngIbUuFmFakh7fwqCZLRF7Fi2agqLNcJlQWbWsg
aJTR05ORWO1cvptW8n8ums2jGMHQw8o4oRFkH7ffpS2Xig2y5K67xlX4g/U0xnJHAsNlvGEqra07
JFkoZahdaUWaOIg9ih0XaJ3d97QQSy2speVaNVivUreaX/iQTx+gwqlgyjL1baNnjrH9SSjGjSa6
Kkb7IZrRaPJmktqeJrF21piOjWfm1MjikJWY55Jw5B0AxFhHBJUP+pD354KOcuvDTF2zxIVZaV/t
LS47Tpj/jplGQ/uK7qW4DbpUVFtOhRZ0oXEeWGGcbmqesdN8l1SJ9AV1muc5HXV1QAkieQYAnq5d
FxU08nz6uAW6447ADkW/v2FTIHHiHrD5SC0A8ed5EAMvXpTn94iYeFU9yxBnL36QSfLiM0XeBLnu
ZKkhgFFkVuoKXAixLZ3XjZK7AdeS/YfUx4Ga83EeJ+6N3UMrIReGzBHt0Pcow1ZVxy9f5g0ziHSf
8SbEJJM9isT97FU0UT5l9z5LO6kYA3B8cRLE/SGC+2BrIkTxtLjv/howlpE2mc+2kyDg7ABJZu89
UpPoejChQpiJaudCW4LATn9dUKXx+MNcoaDplw0+0LdZ4YN4YOxKk2eemf68Qp8bIA23WKMGRs9r
BWW+j45MvdExw061/N+uXNW3UZBUw2xr/YDOijtlRQzne3wGL11moPLsdrHwLZMfyPuz5X21XKyw
jQ7E4+32sRW4QC4v+AnS3Rpc5ZMjfkyBauNhiTIariTrOL5lxFUTUzFhmVns0ym3gl2dAzl3Uaaw
X0wzYRs21qCyG+F+R2A5nF8hL1iXboEupvtBc7IXe++lZGiu+ML0TpCR4fNCA1TNs9Om4PZ36s7W
hZ/XEQOIjXAUuai5UnnS8ndOOVNrkXBb1bLugWF/IeEXjip7OfxUDP91GDS/0iFI27Ni/3QEocpo
bWVJ5YeF7zQZ/+aWk8QPLWk/RF+YG5t6RF2rpeE+M4tdUJluE7BAXMApFxEBy7/fPpaxw/qiqeMQ
JDrP4Wnv9YD0qmEWL4OJQZGgiMHRpvZYk2hGhTRr0QA+mZXD5q2bgSMZPeOGlJ3M3y4tgkKxiaG0
vIWtx+N/wxrUatt+2LTGyEZ8PcWe845QN0Oztu4I6byyhSqSE6qRSMigdVIDgdxBc0MxDiEET5kF
PpIilyA3uX6DkT1kbn0BYgU/6YG8m+WyyV9rO3H6d4P3XlAwGlRPdHx6bV/SEm3uxNbIQ0aQheaU
3n4O0NHcLNf8c7ZfHxCs4zU5Hwca0eqm23FSCFg3lzugzYteydx9SUVnWpLq+27bfHj1omOvHxyg
XD89z1qUJjlXlplncVpaVMmcYjt/cjy88zlCtXYBCfZ+TPjIAVQex0t3yOo5a2pekqdxk2TjBSlI
qiZWiz7qR5rWkKb1/nlxprWjuOAWc/IoamjnEoI7aUvskXYfTkt6F691RcXkc9ruiW2czx6kYBNw
e70xZZ1R9oA7nNsF4Czt0i8XX6pcJGUZ08UfFy4BpBoq822KTkB8pm9XX3ifiQ6WCPkoAI+lOpbf
gHwzf51XPJvoLKP8TunrqaA0YwPKX4ZwnxXytrIW+L5T5QxofghOq1GvHwIbmFxEy7Qm3LIHb71p
6uzP4TmjlthbZbaGNJQxANJ/bCDNHYw43HbX+InwLKLCvP980IJ67LULFsMj7O10Wcpixs+aCWZE
YTeIGsAGV3WB+3uyNSezW/qO8tJ4nyjjcFiWpdV4nEZjAzfo71IvSc9zIngtgtE15FffRhhoNktw
zyos/6bkQuMtBwnp1lMIpbuqi6hGBiMPyBmLPB0uCknayFoUqyo8j45QI/0W77Z+5GqJSL7QLFAm
gSZbRO2BLYe1CQI6CkswmDvx+0Rcb5cpevgqnzCk5CVVDigEkyPqlkTAZAutBXRy1wQH9ngY8UEp
bQHiq0T45gfMhzR13uDzncF6O2DwlZvlZqvJMdioTHotQBUpqbeYxiTdXqKmBjDAy6+ym/Mzm6YN
hQLAol04SmCA/3d4IfFsIAMuPHbIqmmvbSoMPodriFiZSOCVu0pTMZDz+AfpKCDYL/JniVlXWsjy
QFSFd/vG3ZAYoHxePXuSTkp6I5IK2G3LxgHECDTxGoOUYfL98cn725t87MzSCSj/e+K0PRKkTqe/
2oDEb/f8dlnjkONYudMPltYi9cMNj0PtN0yzI4orJTaGybCC7W6fZCnEayVzIQq+P6AW1y6eXh+o
REocpLwuN/wl/orpTlr1KkCb4Tj/JvIqEAG37vPUOhHYlTd8qqmiXFdw6JoM1z3YF5111wp8qiNo
MXOQOWSpCvtywGH/jnarmMWq8w0h6Dp7nJuLlv0cXJQra/1yTPHF6r2u3skp8eO9XK9tpnnqUP6v
4Q3AJRJvwXpUmm/gx2DeuDGdmV2IWzeySiz4RJGJ6CtaY/jD8ULcHvB7atZAIb3S27D9osxZKr3B
vu0PFl5aFWoaZmVM9MH0HKwuWsAoNutz2X/pg4kLVSkXQzVBweDvfXDdeD0b9GuCu9iFQXmOBumH
AXJaGWVhfUJdT3iNKdY1ue2AwAs8OlONM46ywvcXyMboSONzdesHiPAiv3zQ4veTi58t51xi8py5
dTLFyAh0S2Nky6d6oCpzFyf8xhQN5jrDWt6bhaEEFFCgTmRD8WTLDYtzLrMZOY9kUPVAJtFbGvGd
zFWU3j3/p7w6bQ9zfQ5GOfFqA4PEWJEObXQNoSJdBUmYZ/j7siS+g92hlIRqryjmYC5to8c1AmOv
MwLchmiTPbdDslmdIiI2ViHC50Ti442ou6Ig5d6g8HO83uGyHcM5vvRcTqIu00zzjf3JMlyo2myh
uSLTVJ8+rb4x3sTEy5oudPFQBoyja5eRdfSpVky/26V9raVIzepsTwyhLia3RH3/LwuxF5OECaof
vg44Hl6FJAkho+k2SKFKU5mfHD13UidQtYlVF32FT5BBOKHBe48n0TVe1JoCZFR7ESpo8d3Q+k+b
NYl60kTSdIx7a/W8XCh/+QB30kf1f38HQXEcmfb7SrszO9HK3qu/iLCNVJbZWyjdX0loESTNoLEY
gzQEE0ZG3clKtdZsYwM4x7Q5lDtRH+Uli/9lUrkEZnPOYOcHKQqbdeng9I/W+i4wHVmGKd6c442g
uU58Qr/THUjHVFDWQzDLOtBCa2HqZU/KrHc6jyGBV/z5Dpnc3X1iyOKlebZrPSXnzJw35gdE4iPv
8i/WKA0NnbLoRmDEDFP2MSxG8dSFukDBYlxPrLKvgkYmfstgz4QheXi4VCwmpNeKWbCzOwpIzgIS
pLSRFURAeKbaO+sz9OeyJ61LAjLzKKQp0fhzaXmx+E1cUXpZIH8JNmknDk11zaVxgTKmhredZE2C
G7enmHqAmvNB0NzwvnPo5BnpAi179dfmcTEI1nwaLO4ILcm7yXZmFgt46j+zo1PgELc0bzj3r1RC
IKgVSIE1GeayteI8nswA6ITozCNBK4pSrlTqi95MDITCEc0jzNN8ZEDi8TD7LgQBGCRSjOnAS/T8
/Sty6xtlrwxgP2wly1M/TXHPDopo4qbZ8o0f15s9E9pGWQayF8Mo36erCc02GsQYWCDAEBo5hLBQ
rPVUD4f83p5yw1MVhithhPGlfTA09xHK8NnandJIF3IwwjEIGxSGMVAq60kuDFjohqcwK5eUIwxs
njWW5W3vEe/abvAKsFOYWnPzIqQfThL8HxBzk1AkdlhyKhv4AGPM5wYN/Q5mu2K2pfr3AsIT3c2G
wy0BUQFp/W24qeZpFPXMPr6XhYF0uC1TQBOMojOV11Oo4CUk+2rdubrrzjE1LBH40ZPgBTHWIRGi
bU+sLeto1qMLPbnla1HUqlUvfuXyDqnBfLVTUPy7dCGW4+EdtQ7BfdogxG89iFsBeuRMcTVz7zkE
b38ENdspiPhjwiqS8xoBpuP5zBPp+z/tDzBeoLD34mQ9KpThQD3yXxFCY5uiPBNaHjm/2uQmUuDn
0pEmhupa/HAM+TWPjK4tj9VUUsviL5D7gd7H/W+0OzMvoJf9ne57GJXuzj34vaqsXOu7ejnRGsL3
MGf05hQX9+mFuYMxUUNJCxaiG0ErIOVeTiG1CzuTmVaxa0LlyvUMp7r/p23Vn78tgy+sdZ9Yygb/
QWvemrpHDRcGEXQS7KzuiLb9ttUA0ilx+Z6bA9dTQgKkK+kKBDVDbmuAuBAO9dGFCNNhsXPnxmdp
MidpjRnfQqTRdriPRtWgeCQCf1zGQfdtxCU+qaXmsSbn3VZz0q3g+cIWR4S6WxeE+JwgDOjcx7cp
DA6moqXlOjsQTcyEt0av5JO+KOb4D8tGvcE5663W8PR2gccIBR8bhw0bAva3jgHdsM6ZwG4sJMu3
yl0TA0SjB+v1eb8okbIYGe6Y5WyOBcEBDdfzLj9fzn56WGO1uTIQ/Tm227av2wNaNJ6BN5GpfCUi
YIDOMHndKMF+VpylCkFYLZRUCWGvIQUqr6G2k8lxhXYynLRue1j5C9K8xLKB6Fy+BVQaEFYFxgC3
ii5cUJQSi6qQ3ISt3Z2YNP3MnQ5KITJraCtb38dcmKqxs1OnWJlZqFsdrUApX4QICsCIeS5kbf37
0v+Yp6yhIGook/T7uf6MIJM8V6GQj+UovXCA4+c7Ht5uMM13CUH4wdyejvOFC49UhuFR5suMX19d
DeAZZqU4rpF4tejzL3Bqux4gv+p1vHCenXG9KoJ2WFUg0x5mToFyyPrxl0lPlmP5r1GBSTFSLv+U
KT0My795WJzFTW0+Ab2XRaM/0bl0YGIok8h6fhPCiHDVzk2ShCoyFAyqrQ0fDpWrF9CPmxnjdUd4
7PJFw5zOFAL63EPhk/65Jg1DTwFVEiCpHXrorDZNMjOdcCJFA+1gkZk8PFd0fnrUwhSOv0uWWNRz
yuZi3TsHwhIYtCC6KT7QIxYUSlZ3dczYBaWG0y38qDPySnIgFHSJS5mYL7VlDbrWlXC40/+Je+cZ
TWr8rLywwZyK85vMSZRvzFUdW5Q+IYGVrDWh4xijEwPurv2Z60ZJzPycSOF6no9zXn/ZLzI4Ng5u
53HgkDU74wWwIYSilPappL219ouIM0/3GnflNaIvE8iVGgSurnm/HytdgQB8VCZhg5NBX/zRP0OR
EgBPebcAWW79b2TLoTwwIPDnA7Swz4371w8Vl7GuCfgMdpZB/+8V6krZUTnaA3kPkLzP3nv3uDjx
NNHrO254oifAB9amKtSrdZuZVX/1ea6MRUCsbzf6M0nwjx0uyYx14FLafuQrc7vlgVLRLhotcSu4
j+sc4RTcC+lMUQfNc7LueFkxMGsHxjbgWWDptOOjvXldAV0+h6lOwfa8sJsX22oFEeGV2qxFLjRF
WXcNFSrSCng1kp5V0puSQITZvZHa0mlL9xTuwMMtFUhRHDYdxZyBagmbpwuSh6/RMj7Fpi/sE2yh
eqaMPpRMhsIFum9r+L2qJp9kdOlLl6Icwjz06vVjM3rtuJNQ4GXdwXUkvjBhuDIUrrjytP9YFLx/
BHQawVEj5tNSWKF4pfnO6M2tedpBWSt44jOtobcLKnP3qZQZ4RDbXPbs2P3Yg7/ihi0mqOTYVh7P
6BwVEs9R20atD9nUdY0ok7XA31Ui80QNIoHKWU6Za2zOqTGH+Q1Pet78cQNeoEyoiXfoO8tdmlgn
7MM92Jv5OlnLM9irkMIi/jZKMq4WGbR2E19N8RgK0tJ7+doMQIUgA4c3yaPwdRdLkAW0ityDMR0x
8/fyxHnNQbP9WpAFyhwWpkSAl8qtc7fd5rA/WrMuoRR+x69wIWA5AJ1QYsg///2uU1eOfANl1hGO
OctLoI/XsGXcq5Fh/dQs5ceRwLmRTBZyg0nKbwWHwvyAMk3nJnn1tNFORSlKnlSXa3ia5RvAjAgk
Pe+5hD/isM4b87cNytdLxempl3+U25dpRsSw+oLl5Ueg70SBisl1lKgKQpG8f7Nnlnxpnwf6W0Hq
c0ibkshvrEtZJFtmEXJfEcpBXluuFUNdpsTYfUOlTfd+fEftMeZ8Ivf1PCxeBrUIk7sI/1mUHSxv
99Z0qYEyUMl2JjfjudoqbnuVf8Qoh1Ke8Xy6Rikt8W7tX52y8T+wnSxWKD7+HKYiqVqZCasP5dHU
aFZ40SIN4LK9q8WfN1vjy2JZzfuxHBaoPIF9D5xjaRmX0b1W4nLmbl2lWrJD1Jvu3O3ypvLWvedE
YWZkbumQ7rFI67bGKgxafHTE/w0/LRk3M4+WCVXi9uuoYvlPJlbA2iqhUnaofVjt+Vd4VV1zHI6V
Ob5/zj9wUJq6HCOC9EXnsHaUwMmp6KyBpsy6Spyga3ChQriG6hHtn+7SWdp75XvUo71DFjpTMrVg
8NeIq96fuU/4tU4OsYxHHDai8elVIXER8/OE8X/ZUDRBV0evvLlYhXayVG+9B0kwJgn6lwW0AFHz
+ZzPbA8pCZl6WT58ff8X5G29PzooYe/uyoR6m4dKAUD64dbrRq9t3Wfbz48H3JRgSvIPdqkGqY+y
JS+RFdR59vTSbF1T2tZs6R58FI3ESF4Qz4dIg4+k2js/eYOM+HphhNbfKBHZLS9/mqXLjqVnj/I+
spmMqImcmU7lir8vROqgCqQQfWAGGXvzLxTkSGHHH5SyXqcs2ziFGzyAmQkHnvT9ponddX6XaZ/I
aOSA9V4ChIPrXt9Tap/Ofln6tS5qNR0oxnbFvwGhXZFb9HdOYD+ZRVIXige2J1P38MBKmkFdFh9B
KM2+WkSJU0faC29XBsiBb0JzEXI5vqnCbmFnhPqUBpn9mQv319CSK5BH/GfbIq21at6kqJC5kldL
09kLlXEmcC9c9ouAmvnZrFicCkazeq7JC4PC+/A831ZQJ54PCT39WqFwxGt0Fa779czD0NTqyEBj
dMekoBCDuBPd7dXLqIm5sz/0hYB4H2N0rH38XhLhaxizps8DYh0wBsxhexMW4BmmgiBZnh9RgBoK
g0i9icSEq+ceCgfdbM5bQzo8AYcLomxcjqSN5zAh+P5svTl9vFmaYkj9QVi3qgNe+uRRI5WEDekF
Xkzt6rq1fJU5OD+/oGbudu9gJR5TVJiDxtycRPbmI2l3g4OrkWy42c7OpwX15J6L5m6xkxDpmsuu
GBestgR4XSD4LRgm5qU6r+NXt/1+XW/nNhUyvb4NC2xv34z1jshi8U+1h/VTNs2YXJRvST/mc9qI
dt3v0Qi3oKVHJxS3uZZnRVCZ1AMIN+Wo0CPEAhoI5Z2hD9wPLu9aW2XP5bYBgIdVSDI0OFaCDdPS
fTmnyxVlaRrID5AqnVnqiZwCKT0P7RutfujfHXNLTvBa/sBwg/2FEeon/KjlNQOfbJ7h/2sJ0Pem
OwlZoek4+A7SU8eG7i43ar9Zk+pyl7YsW5JxkiX8Yj5kjo1xn3rKVvcYS05BNmafgqWJLd5vUZJu
ywk8sGW8R3Rk/1uobK4MjdhtyK3vOJxSfA728dRe60CDP4fy8chxQeM3OJiyaU8HDuZexx3uhtOQ
VpA3OGEhQ76XURrlN1D+EQNCUKMqdNKvmaclDqMsRiQ7xrLF11e+s5fDgKxsVIxr6TRzLdMgiws+
3laY2kwmaSkfiuI64w7Rpbr1lVchTqEx+c0xvnQw8sNb1lf9xzivc6QsmzJjJeIkkDTHFaXFflPT
E2QzKN4SYhpKtmHn8U40VTXFIUD05Nv7bJOFt7rBO/xStj7NcUaNnO1unFFNIGLeHfrbo5uKHzOQ
KwiwapHgB2bj4Nkuww/h0jXZw0AoEwwBM4bf5PDT3hkWaNxNBAwfBG+GdbYBR0HZDGN0mBpO8gVz
T49tOE8EBY7JPfwxogVBsTm5j30cHO8jcXJDLYZbiCj5xd78rluaZr5fc1iSLkmq/xjEhB1b75aH
PoP6sdv13ZMuWAKlNFeZF3ixoM5jjY0dghuF+/V7HI0afhQLGemjwu825sXInXveaoQa7IUW2Hm7
yetHwpDea6oOyzAOWTgpWJSYOweyJer2sAs2OIl6WrRG+Fisaf4QECfIlU5NcdP8ATsoyVt2eexc
H/UchRjOvhwTCeeiRT1zGGGP9Xf5MhN5DyWr4O2xB/QgRBocA3tS9i5AFh7vQg81+6BFYqVGSNLq
fx9po0mN97/kwIjgam5DxNBScPkbYZK62u1O7E3h/FQjNz3lFqWNh+Y6GG23BksP3cOqpoqV56cc
XxzL4kbxPfiPL4H42J4Kpmzm/b9lu+CE1EwZtRHGQiVXDu4liNgpY5Q/YRYJauG24xfPTu10g+Jc
lNRcEwbC/kok8qNLRypQRqy5Z4v2bI5JITJMUbnPz6o6w/BBK/v5oNhVgnIiOHDOhvZHeHqfSnm1
b/1b8BuwGyNqsaH+gtZJyX5O6xAoC81xpgAptcxN8wpwQP+kyYMyHaVTRT2GOXQI/7SNnQriCJyU
o3EDfrjMxSEyETEv1dj2lv9vDiYXl5SY/Aut/paaVXyz5P562MM+PtSuFT3IUzkvFos0oNo3ZHMV
JHsrXIJfCDvEbobkiBHUzDFreG4ZKo4+s6JyJGa4Kz+SJd+dCnkGn2fZrpw9/1JBUN9amOYDKCGP
flPTnyOrXn5o1zZYWQjPqMduPNTt0XLa4PmRBngAezgScDEyYh9DYGO1C6UwfKzHAA0Em85LGqXy
aq7Ahfupq1fu1/O47sbRyfnNMi+YoEoy9pTzV9nKmVprWQcQGIxemDXvIxhv7GY5XFogDa4UpERe
WcI+loIeMzVt4prkRC23bEcpCC5oJWEceSLpx5ONCvtPdpjmXU9xNMMlJkHkZJaYc8OdvrVvnGoZ
AhDicrszHTyD4Ku/s/uWUdAoz5eYl45P05+Il+NHq40+pSYXHUn19zVCZsyIbcUrXwaCnN6J+Ci9
GR/+bR7XexqwMPlZkWtgWEmTHU5tPk19QrvWMMAPJjl+nBcgHlMbYlU2cIyj5oI/ei5XV/XKTdTR
AAes6wSyzDLGndGwhFirrjcK6taBkrOk1iZSK/9KxFDxHeMIUu8/Ucf6gTNSaKX4q55wWtqRTuwH
EMZyvGRkwSjBMPSYjXTGhOEzRmdWpEmuRIM38N5XDgMfOSPUW1TKpOK2QLgOpOKBSqxIZ+1ILzQ6
ZUGozLUa0SK8+hejYZWB2VIyej+Kjq94yI8U7eU8q4xjbLCVbfmuLUyaEsU8HVg16dJ5ipsxkApk
VK9raX96PLZ09J5L1KsMuf84NiYSD7Ypvu8TXkas9ThGgoQoasAwy/hvVAIW8OFRSraPD3f28YFp
RW05ylsux5BEscPawjJlditP725jgHkeWINiwXBmUnGSZraFvELJGpctOs9dwVWW4q97W/z34Wrm
qDGggzFRXyueT01C+CRK3QsQ4caEXxAhJbHt2ka9hV/BzJF0F3P8fnPQTEtTTRvF4SAnmbmsDxqP
XGCsAQG0vTN/omrh3EojFp3dNYGYEFszjQT16une3N9aNqTiUX5HHNoH4q3Be3OHikxWzMTameM7
oMeytBhkt6HQnQTWfOSlS0zFDBPY6do8nEfBpYN/PT1RVnuASmNiohBZV/f2Ho3zIMV4W6pknx3t
nxVgNiEPQWLgcUE5L8NST6reUW8h2BVG5s7dCEXui7rZZdacNkiFp706V+8pkp7YDEoHoCcDwdyG
IJqAYw6NSqvS/LqRrVaXXlsV0dzM9U0+sruOgLaJYmh3Ns0nRQvpDl4uRCWUhmmTCl4odue5f9WC
HR3arbzrSKbhKRnVhG7Lfd2H5kjuyWsOa4padCtPa1UMz51oXfqwxP/DpVzOJX+8SUXcAxPUKZkH
CJeI0Ie/LIU0skaj8JK8RMcuU/5fTs3ltk2eamNDOzDi0nYDPffJHMnIvAGrx6idt4uhdezKEZyW
ry7eal1ZTzOqGfWAyHDsk8HQ9gFwQ6ZEfvmim1ns24rKpJnmGRyCifb4hdsre29GvTDDpFcvShKc
wm2RqPrHp3wwG4Vsg3sJT8S2NBcqwnIm56EcIGGiLf8FIKiW8an23LULXJ5F3KZCjbeLv9pHxLKx
muZVmNDT36/qvjiqOJHHRmE6y2wnX5E1e1tmPyyR3O3zChrV7aISDnb8CbeDUsuQeYHm3c6ZEXO2
z3zDxJ/bUqhB6PN7X0iSAHCobK02NrcGgyssm1L/m3I6FEbtpOvCmYuwwmcxpYHDuAf8a5tY/Gwi
8GlP1ByL8MZ7hUaAcCpTsevY9OsNbrbN3Ky89JUL8lV73rqMD9LDs3PLavvHYaqQZdxboBU/0fb7
YvFQMLkp3WgOeJml0S26s7WYyPJWHGU2Km0a9uJbkc+cSzr6ncUkFl2Byn2AG/7eJbg4NXQsaF8o
rIBV+hhTTShuOIj/aNRkfwMuI/wX38hW3JBQTNelAGRJ6OEfuEudrZqf/Hz4Py/5d7G/SWxp3EWg
FQBRHe3NZ0wH7uJIgb3Q0zq2fhZQ6dAQWsRRkvKVqHqAdtZXvUwV5XwMjf6k6hnG2YeKSFPV3zii
NNKVTC45bGZsDhFWAkuv0CY7Q41WymOhUrBYotwgggIqSI5hMG45U7dJGnQwyU0OubYheKjfijw9
0opzLh363JNhRlGU5PM7+s2YzNcjzE8fI/CabB9v8JyiupeUyFRk9SbYJHa3GlVqJPTgkcByi6BV
f2hnhQquj8/gITj1y+c7pEeJ35yQckQSXFB5ci2g3PjZXokkaOJcH6kAtl5nTigr4lDGZtG2o0zW
id37vpUSYrvMonXGxOYtWWJinSNFycb3uVGbKT62OQpVSEBsbDQfxuRg3RrK4Sr2UgVZAqO+hp/s
B01gFbVjUAMZ4k/zhFGZ06Irgx7JyKqrcuXMLTUR9Wl+/E0vaGuPadQDt44Xx2Dg/NWiFSyfA/OO
ChDDNJov6GFqEHRqFkUO6pro9U01KCXmzlgtbL2ggXcGYNbfOBvr8laUZx6fqdE1rBF+BQClJiA7
NAu2zFtL7TWqM7T3elWpQb7LwgMXx2fmfWVLe9DqIDjW7q73ZfifADV6R4zMsOfy6e33H5p6YDt8
DNva8+m1EX9O+EWqE4Vq4QDWkbHq1I0YyMXY1iMxwZlFMoDPhYMUtdZjHNSK9SKWKyk+/5M7zuMk
vak9n7TLoq3+MWo2KCu+qSya/6PMmzMPK4GQ0tts8IPrNxP3ZJQv7wNJ5gS3MVih6H6n60Ig9tQC
w0KCGh1rd+BgL+TD/sCNn7VttvFcpPKO0rhk3zPdFy8W6j4o8L3QQ3O2V3OH304nnYw4PEXGCQCu
AwN3W5/R1UINVmwQOX10ITdmjw/iu7j9U1qn2a1zWqyl9OHujybGEy9wdeuz0ypVfM9817V3mE4I
+A1M89txmRmPDn7wMeLpnuF448uzqROuUvq7GXuZD/FRQlZWkEO8aLFQO0nmJiQOtkScmD5pASMU
TMAWcgSG96NoETLXCSzsXrDPaHk4KVKda/JtO7FRCjniyP4+QZGovK+5jc3/Rn+Er/V3bOUlUr2i
Y7IpL54l7yn/RvmWBUHsCgSj0d5eNDgABU7iOmTjOroP2ei7oIasBBjfnWTzZVB/5hdsKvlltPy7
ta7C+Q+ZZrKYSiJzBX43KBqCm3wpLal9KzoQCQs4xUdAAhFIS01qltDtrcHFzKSsC+C58MO5q4+0
OZgSMHo1PpEF1T25t4EhvUoRmX7RS9HCYdswlSNA7kcv733bNMEHZxlsV725hk4xv0MnPigNUV0k
ATc9PAnp90YLiAY1IHZPpbIgzcJA8JwQySJC85vLYy4wwHXaPWxb9u9zdhMcuYP5vcXer8CGCgBQ
8O/UnFXC7grix0NeRLGDpGDOvIwbb85I/KE4i9LByMRBhjqQ2rPrqfxRyWnIeei3gJo+GvlKwlMP
8r+ekw5l43OkXCQY6BdIKuIOtXxagFc2+1cP3QVDN+6RV4BMn1IhBpT5FSPpy88MKwLYPta8gaRI
SKPvuXPCp1nzCLq5g/YdBNuBm8IbzvwRwuDSIyB1WeTEix7rp3QjiyY7646VYwyFQJ22OrSR+tWI
+wEvkE3drL9d77yF8RnUhG3UNK5IbVTCcbbCaAfDvejyBWfZ+POhyufzujvCxNR0bJSK+M1rHdzX
W6aNWvqCsv2SeJcvGyrVDcsFbXNKvvBOHo2hHt8XW0uOEVAxto0ouOKZgSKdviEbi1ax3mSYEQrw
uHgHfGI5gdax+qfKBV8l+Ba4Ka5UlWSrReYxBpmmbucom++LG7YSxPHNZFEcbF3f8doYx+1h8Ioy
zPK5+W/+9fKdKuvMKLoz+q1ryZOBJuoyKRDSzajdpE/Jf2or1ZoLZaz/7RrkGHjpqDkv0ASDz8FZ
jkUZ3oi3j9B/yMNdOaDMHEX1VphbwIzIQ+O05/yOKNdCJDFWZGXv+2r+PNP5NWiDEXx8fYnTazby
ETB92I+Ju0SoDoRjLzqopXI9QyBHpe/HlHPdQ94vT82xFxPWSH82DDxUDxL8WnFUqmcMyId6sO8c
W4A84Sh/HrgL7oHTBG8leoTH8v5DY56X1MFuoFqazhughIPy1AfZGNrKAzYM9OooJBzLw/GDCI9W
bE32YvtNEuzzvI6O3xmIUbqefwO38ITksTMO7+YtoJx1Cyhg7HbAYE9kENt6t09ZZHI0WsRGgzyo
2ZT4jiqSgoII2Ewn+j3fFYK423x8KfApNVZtgger5cPkRvExl0gBmEmfLdTjhXEyWJbIEkTq06H4
EWOrvmxuTLONXGYJMGqPw2Lq2ovPFF5Lrc0G0OIO8HOYWSFl1wyVMX6qMSl4Rk3DcY1UtqKKzrQv
WeRjhLAUYiuBaSCBUWqUDW2xP2zjS7Zb/10rxe3/BuQnlhfiF4Wfo9nIC6+l2TRkr6kz1D70vOJ6
3sqH54o22VKeJKzpSrTPfnUmkhjRadM2+wAEAUFUkMHVzEUR7/aLn/nrfdwvkwRyRoLngVRUr64c
vBrODNqLj/5/NjpZOmW+4WlBcmFBfVAWMAyLMFLd4LV2F5/f9nApYLE3RSm1NcAMFDydTxF7ISE0
kN/GWX4TKoQkRS4M5ksyNXpa2eBpPuwzNpYay8p9q/pulY1S7r9egMWhqeDZQbk2GEDwq4WdQ4GF
G3KD7rmDVlwAvMK6FijAnC65ivdWdzT87c6HKnSBC8VmYbdD/s+XN/YZW9F0phOJiaOxT4ndAxSl
PBTW+M2wzcb7/AVJ90g1/BLeRyAH9SVJE1UH5H8GavOQTqrKaes1J9GgK7xzkIRKGm1vQ9IoMN5V
FfLisPPX9EIR0fiZBZRkBDTdmmuAK6p35Ox1nBvlyYvXdePkrWuP0NsoLYH2S8SnWqvKwfhtCQv+
LW4+ACOPLZ/fgqHqvUPYa4w1tvu6q4Cb+k1Vp2VlG2LvQ9pOWsVy+SVQNIlTGObLpj22RDG4Rliz
c4H8MpXridxf+HDY6u9kYLLlykYP26ntd7u0mvD/zJJAoY8mkczUl1+4h1uw3XC0IUIzA3i3etDT
cJQonrC00aRv5RUmudBDVeyjD4TZioGO28//sXibZHsf5cxUp5GGaHvR3zw69ZjFmjjBlGCRyDrW
xogIOzvi7tGJUcMmo9L/slHt4q5kRypTCGFkceslTWDA+sWKiITag7Lf3VEo2L+fI5HBPf6FjHYj
Uy7aD/oWHAWAylEj8tsYCmUx3Q4/TOwxSfo1D/oMFAFOOi1+8f85NY48CbWSlWwAJxyhRshQR9pr
jv1EJqEvi53r3KA5GdPnX4ENJWR+qsT/9Ld57OsmMXmA7MSGwDjjT+bYbWYpFvfbEprdb9jX8VgZ
B4Ydq+DPyeqoEUmR9oINNVOsCiPhwCaikAM2wAXV+ldlG5lpZGYVtZer7jvYmJAaOGO6bXrHqrIH
RYWfgjYgcNF7iFdJ5HU91wQAdr9NoGZmd9ePl7WF3GZ+J5sQTHglUzsCGvptPPp6j0cHPrbT1/dd
1/8wu1tU3Wk55NlNHE2EIpqg3AC992H3CrnSsz4bCPR/q5IEdpvxJOKnP7kIu4q1XvKG/vW8ATAx
FrNIgydHEBWhUVDz4bF5UyTMbMaPXLQGSGoSStsYk37eYSKc5ccOXq01XQCzpPs7B+TJYShj9Jcd
mraoB7Z9DNLk0Nl8w1TdtELZr1T60tl0uocvYmfxIrrecfpgdod0RFV2jYUJ0Se2/MkDo5cvyFyB
LDemt82xspB16QgWoFsfY5cBY02ivZfSDTHMeFPL2I3kccyyt+XPH/jMY8KCpxsdHt3j+v646QGh
M5E2QGlvsZw9u48i/miRlBhCczuTstUI6QChKGmxBfykG4Hiu7ZTkwEjyaqGIOF09V8pslvsLKQN
7+EgPCcr3G2g5Lu34dMoxbcZ5gEhPHn1sXqkkLUisCZHqT9ZqJ9/bfrOzTrHRPLwB1PAleTPDc5d
HUWEjemnv8ks9l7jiBphjLzeFrrM5j8B0zI+PPXBTWj+6dY4EKmJUZxKaYwP1gLNEwDn3P9ZY3ep
YtUFkLY9L/3Lj+tczl90xZtX46xnmq++AXJS9+BTcjbFxqhpnk3RzRBlLG20J/1rg63a5C/bXrpU
ZbqKbMP+F4BqNnTifBBMWWEjeU5W5BS2PMi5wD93MtE8beRSzCbjDdR5yRk7LRIezPXeooa1by5+
xa+YeW9ng3NqLbv3ZsNfvigwleikAs4YD3EMijngMx/8zHUhdlukW+pnwpRNEyraA44e6AdH7ocW
IVyxunM03i4vIzVPQ2oRr2tPP6eDRVFrdvkHFtJhKsD6/EtXsGR1ajbGD9PZcNq0vDv/US28UY3F
B83pxNfoDHVg+I/y6p/F0Klobln0fQ6sFUsZD3s+gZGR7rGc/ZZD4woctOKOTzljcFJFqByKkKQl
tnWKodRQjz/HnVNaKMrZbMYfTfvTctdmYLc7vYIBXt8cTFyXGUllKptK2JW3Hm2VCpSddUuOm92T
IWR8ulpRVORfpHGK6HqIQp9fGosDRgnGtkwQrDCV3kI+SDA9qspSIKKJukGMi9ua8a1uk+q2d7qr
PuFH90DJ+uBPhh8kYtOFtwGXzSAs4ehGw6iy9UI519UYaitm9vgOvwpdVOnBVhoO/bNeyJcCrjpA
ClnwOGr2nby83NhbRsNrfv+VozJybA8QaCqoWGJ4DHlkO7k+CTbTv86AMcadoHrgVOmZRWBf27Ry
32l1IGZ/ANdE9mL8MTS7NXESACwPfvcuA8p0OwGHJvH683egXA1kxbQLTINqpzFV0ShBdH/tdY4e
2Vvi24lyu76MD5lSJzCXAH9sosWEfBjYcleD2kE06GzVWPi6TcjSSXQ/UG3y8Hs+V56up4cen88R
0ngxdzCPN03tvzXU06TL1tRxW8v4jBB1qG6MzLHq3sb+oDuYePPxwzEWN7AuXsK7Qsc2rrcywrxv
K03F5fXo6dCjWq/1mMgzVDJUOJRe9IAzKMhlUXs9dMfuYRcUE7V+XGKlO0vj1Lnu5N3AYwnhhLg3
v9cRop2qLypLKQJn7vWBCm9wbl7vH00Vm/dHSXM1quk6T7JLpJNc0AnMnAE+lfxFVYrxYVSdJ9nW
RVoJPoQJ5sURxQ9sYR/ssMze2hvHcBzbSIgKJcRBcYOXRF0t05IQ5e3nrMKB4xNJV5o5KNSQWtsH
Vh5ho8l0utPTNGfZLEgY6saRDTbvTod9Va2tOGPssQpwfxHEr6m+q9D9aAJYlX3HZ6b1MQP4NDmJ
Kajxd8ekXVoTvmanRgUrDWlu48gWwa9BOopYJAw6ftVST4oB/lVVMJrwxmqoflSRmqSS4YTmfgUG
xp2BiMjgwa0f1zNViMWdhTk1lBtBBIrreIj01SO3qggrgp8zL3Tv0L0FxworbfPFfoCnD6lcQLR0
aUsPg422F2Ri8Ilz/kDQNZNaC8WhSJ3TTY4YYnbG0MJJuUQ248Dx8nrP070bGD+DlLc6Xf+9v0Fd
HdBFlEfP38AUre5p/tnAkcGQGnMm8+3765PL6wg5xeH5EHZ3RDib9/VY/XeM/b3l0worn/nqONWX
FkicTCFm+KjfFv7LEfqEWIsx2NqdVXYlwGQXNEuveW9xubdTZ47MOVgHFmZOvA3pTQ+qi/yr1v+t
XUkq2g7p/LTDk6D6thDI5JOV29o8DVtcbIlBN7+XvQqwX7xd/S8eqRDsZW06UG/u21weKwXjn9Um
LPdHMYhnMLaKYlJcMRhgfESBreUHaOdT4kSZ1m9OmtmoSmBYBIx6EjTmTJqq18BLfih0XLVK82jC
YaANPXbJvZp4M+U42osjIXhf1Rk6yxNr8Ae/XWmCOKxH8LKUf8LX6icl3yOS84xYcyzyHQS0MJ1l
lQ77Q38Gf4h/ldfZqHpJq7D1dTsPaL9fp8NsiaG/oQGgxER6A4wJ6nuW7/oVkyiUEZyPYIrUFMAJ
6MubD3hSNkiEOO/c0/bUFfmcz7UXtlsnnbPeO0ECPChz9QQxQshUpMg51JGN0fDryetKS8eOoXxx
BOq4So8m9GZGVgJk7oE75699IFKeGV2V2xegVBnUKJK4wLvTCsiBy4irE2Zugw7tzOVXqj3UkALd
/BTXIqwrDPTHy0ZyhWKQKPh8GzqENVMeeNtXs3o0G86fUFIn10o6owOjWcMgQ4lFZkgGzpacLzsS
5kdABUJwshLK9gqsLuCYm/VIM0yyElzYNvbIko8ROrNYj36IfIjGUn/bajtGvSNmOfFSSWEba6c/
v3cHEsIcYcr+H7/pmscEmyHLPa+OcCe3G+nhtGsa1nuqiBmmiu8ki+c848+CiZ3G2tN7Tewm1z7A
4DOsC/dZG1vs7BC9HAja5k4BFetmhaHsdVV5rG28v+U5RgDTH6gq8D8lHMK2L6w2a6h3Bkj1Kyp5
+NIBL1kz7WF4B+PxbVTgFIXyV7aQyIqxnpweZATGgvccUXT4fd2RdsdQb0n9K4E58z+nrZrkPH97
xrP/EqqRzw1mv5cElVLgCD09F9MF5UT0OR/Lx7O+7fuAp8PtNFz+gKvAWhA1rSSBqi6Tl5F27BVT
zhNGBhLUJuXPtYxLeMPNk5NwNxsNGK1viOZsppptRM0OGONTXh+utxyWSHVZa4uoS8ok3o48iSpX
JEI2kSvLFJ48aH0PdauXbD0NqYxV9zvPDLmOVKgpAgIC1ardkk/xXA83qI92ZUC2PHwDOfqdfFTF
shI7j4tLLpipklREPAIb2snRuA5UAkl2InkCOXpUUR/gy5PSv0ibeO7P5ebbudehjsa27tnZ38xO
295uLQHmWMd5YboNpTaFxKGzEACnK8d44uIzx8rcd57Ol5m7q8Lg0c0FTfgb/VUJ8xNoK+vHeETS
AxeYAmlIlDq5NoXL8554/th16K2x20azcQRZefh+iJltbI9j06Lmla00P79q4V5oUkBNaU5REHX3
3g1ykd9F/8LyhWkwbiQs0UgsAQX2GLfYvWo+ZKSJBzdnf7aJRl+iPqZhRT/Nn1pfK9mJ5EZB9UD+
QjxiZSo7Ma1LlqnQ5GJDY7VuHdy7e4BR7v8b6T32ZLkwiZ4bWvFGCTSGXF0QfgpT106IsViltez4
AN4mbnTfXHGpu+nu+OFKbP4LDlvXVEZbaykZAGzHbUm9QLWhmve5AGTOsvNBTJJ4gltTA6pOQkFv
1+amvLwDV9czO7E5CDiFB2sgsIA2fQd5IrDtKE2L2e9L3IKmJSMuzKS1rK4FgkHKVu6E0o7r2ioa
Sdh8Q6yD8j4U0AEJpdDrodeeh/2bmy/t5HYv8kvu+mTNcsOBaN0k2XPbFAtfzz+GjvY4VaBNySi5
lsqzMhm6J39aTOrq5ACJHBDCgyrhjW3wRcgCdCeKd4Ab3uPt+BIXLkj1Y1f7gEh+2Gzwq7CVLMld
hh+ag6e2PQOHv3OEhckjGtSYCJvWgzokUfgnxiykmx+jPlyDwjszeS/W/Q8EvDIitL+MyGy6BTg4
r61ss1PnsiEOrq50nGmKlnqcWNYSAk/GpeT7PPxlF0KsQ6CeqM/wKG7fefhorWnYJ5Jta0dAD8CZ
wDziH1Z7iwHL043EnxWYPOs8OvYYNPaAZXrtChcgNbvAmO+/bpLmFsROd+hNCU7ceMBjuLnPmLq6
m7zdlFrZNcEZUzVLsHIr8OHoah6pER4zlu+1JTLncIcgql9JcxZlLNzV33Fc6g9BPzFkzuba25ul
bFsHJc0Uy2CVcuOfa99gcvDVwpS7Ynr4tqWxJajRKN/2zOF+w9hszBmyTLTHKoAhx2TqUfzACEEw
mvlP/Q4OdWx6EsDjRmLmcPvzDDjGx7FZ97JIx4gp2HFU0flBlX1m89OMxFh8tjboYSxpjOuxk+DH
AgDiO6wSFBsy3u5ZkdYqJqQRpDNeFOrbhRvUdU0he4Rvu5C7scNC7lCEigElss5p4bFunBi2PwIl
FAI+lYyxc8b/wEetIZGaEfT8foqAChTDDjwqgJbtvs8a6Dzbzp30r8x2WEDaLaVFk4iHf5+YNFDF
WXKpVC9MuGkhReucIJDYJGU96m4G46UbyTCeF3SheU9uf6nFL/5PbjmyN3fawNY+sKQyziL7nsNa
be/zqU2o448bTQeRobs6t7+IBMi/DtKnsarH1GXHpwZCZXO8tKfhCG8FD28aq0OnKNcUxKvWAXF1
iTFPZYOgzWwsmM09YC0bK+DRso+4bM3Ovb8YxKSVzgMG79VkOXdchfRXM5EIFW6r8oB+lgniS0qC
tB/C5tm5ANzCjjt2eCxXleUU/aV+uYs+olHhfDdeyf6VqBmflLKV8wTjbiVXLeytomIQ2AwcTwyz
Kh4221cCzEu0bH/kAWT+3VauvP/F+zAaf7bPp9c/Nbb5opX34VWXW85y0KE9aVzpwMFwkY34vVOE
3jsRhMDbSHtwYeeIRWf7tepKVvukvCm1W3SsGMh/IzOqhxvIc4UecDzOGdoNkQMEU1mcHJhI/mKW
m9Lb6IhvrwmqrT0urB5koWnTOeRA9h06AIGsJoGRr+mzzp+niz6rb3wCYnrPBphMrITCBvCpapYT
mtQms7js3aillQH6LWYfVTTfHsft9BzIo+ZecbnDtN0G/YmbYqfqYWDIzvJgUdpiHsRTVVWLTlJV
DxTzbdx1Se35I3gSXPU2D6VLWU8bvYL88LQxTFvU9MnMtBuCagx5wi/HdJzEGmHp37q6EQ4bqZxR
ztARH+Rd6jgWjQ8q10moOwdji8FmoT0OK3C7tdEvGBpp/JYTa4NijXCsJ6j9iOO379VywmGbZxZw
8PnsXdHs97HsgPFizaoy6Rh9ftLhMY3l3xf0BdS52MNIr/gANWG4QmY+M/ApNwsp5qR5kDorqLsx
+xCGhsovPFz743oqrPFjtdDyjCw2X+pS9UmAxGv8O8yrDCbK6A2rh7SMEWJjFLdZ/Jh2CY/vyvT+
LothoOXRaK0Nli0X5lmTxCci+FJUtBLcEY9v7WO1r0KnYl+enQGNMCMyQJUj04Ttc5pn821dMeWS
wPzewLKyGsfQqEXwO6uxw7kezq0IBf1esMX08tuEGX9a4X760uGwLFdOZ+d1sQg1EUOk1fmdGr/1
qDK4NYdGA6JSLfsrUXWPG+NkQwsxEUs/ifUEmi/7jNf6HELJFEIQkuex9g/rmHU0EVJB6gkKK/CM
i1vv16w/BZzFky6pHBG3VjsuvQY+iO8dGeyS0sio+pfkVdFa4SNDTnti59A2B5DSP4AWULL5B+A/
03vlCyf1X4M7MyMOCHb9FU8h07Hwjio0VZcmv+LmHsKu8YfL7+qqREfTxdpv69K7X1WYHBEmiD8x
XWxqgkxBvwWwu4d0Mz/AtXX3zqRYkpLG3rSiI8Eer7GCq9D6fhRVMBqVX6y8GJOM2jw1Ygggf2AS
ZMdA0LU9xnD1FntEj22hq/JFmzV+Vlx2KD8mA7xoFREja43V5UYy4OG4Jy0V8XNKn50QDb2S2j69
iMXBf1PH7qIb44temlifB5QXq2IGmI0WuwnK/MmQoVonqyp8TCVuR8/DdY591gYDolGYP+fiHH9p
TbVs+ngxRGcnGJ5mkEXaMT2FYCVPOzgFojnBQy+QZ6rPD5eaQbmrRgNunSJHpE7g8hyixj1DURT4
oJbyS9Lf1Iey7/Oc0Zw51paz1NyXmSR9RG3LgNDvm+CEBi5gt/UgOdJVt/Qg+4M+awFTpYDpBZis
q1ryQWWtVzbHIKEZVs2ZEv+5vGVPXKuS+7Pj8pIM38qPpbIgIJhCKZSXPXKOhQrsptwV33OhYiLn
eC5YGd6v+fMrleSZk8guyiX0ykGrje1I9CvtXLqNAIQrmKVC70Jj3vvGDHHDY805cLlGBhBk9TXE
048vkePufQDwntlN0bjjjZFHqfh62rWztypTYVqd4Oy8FO9uMJxu6P5uL7LOh1xVJY5i6H6zV55Z
97xnl2+gvsyYWMagvUs4o+dgS8yWQHSMuXBfj67nbd3Y6/Ytv+bAhe/PvDePcOBkljT7/I4cKTWr
xoiCdEocmNjr0ok47wi6FcK/EjlTaLBVDUviqICwVNBJoreT3qYJ1fNlLA0vh2TuMU2evlF34nWI
6DtUyyl6MTyKVkqNGxv2qPHRD5u+hRqVZtPfPqBLmvYzvHi256+2rxYMub2Mxp2quqTLPCYBSjwi
JrzPOyg0ophFCsME3nH0qu5b2QJgZxUXfre69cKRHAdlcVmt14WqABpeC3DZZqliX0yasOBM8y+J
ql4z2klJmzv7RRqVaZ+IoqCcaaMdCRXrXT15QcAOxR4Dsq9jiFIFzSKw/AZlWhlvSQR2k6M6+OUp
mUp6N/1OXzP7yigHHARAsVhANI3srzMGIKk9pjzNWSIclcSQ9YdC/oyBYy7CknoyZ4F0wegDgrAR
PJp8v/GueZXUJUUO4elL0oy2TulphZONEeRBSQChdaAwsAnhKHCdBmgEBTreCbOGsh1e2Gbl0DIv
AUJKl3Lo1HgupD3ec/8wNFr0E78mBRGP+iydePkjrWgrEHmh7cD82O+4+KEI19LXliWR5TcVt7hR
PhnXV+BOvwG652Fvgy5pM3H+xJ21BMWBaMwk52UJi5OHYLY7Ttu58QZH7jLAFqbMsbE+5TcjxZQJ
8ztbS98H3VUQbdzdxXTYYn0yg47KuUUvrYjkmsScWiqXyBCyzbXB8DRACCqOpqBqWSsIOrTDWPfW
aiqISM23QmZtJrtbhANHQ4w+kZ7qcacrZw1dNZgpipVjSBPbcWOOOYIyipLraJZUVpcHWZDugpGW
ASZjlGwVZso9m+y7KbF9pwcrBxXIPFnva9ymNfArn326H0CBnSS6ggYCUudrAfsDXzGUdm6Nq7ik
sesJdrbuHiedGVe4jrSCx7QYasDlKWE6TvLcIw+Ao8AFkoc4mUNt+EDk8IuLwMC0lOl1779TE/s9
nIOEFqi4CUruQpF/OCS5PLnpaDPBLvPwRBSVqQ2lY8TOwABXkeA1aZLTC4hw0WW0UU2Le7ERLvDA
y5zNPwhNSlLz6IDMxxk6ITJzfxE+/d9p3j3mdtNhD/GPrzgHccfSTNA9VXHZ/W5merc6yDjKtI4V
TpNLag1tEGOQFFLwzRkcE9bt9MTobwHRyNV9iOqXrAscAEL/2VrDTW/9E120eKMixbW74Mhxleet
HILbd74c2Btst3YRg4SMRq8b+EGTgfeafNDUKALid69gyS63UjoJyQg3+N2DD/8F8RtMNOnVpULU
/y2f+aR3SCxQsUp14XWDDUK26XylDQuH4GVHHW5CHwhYI4MTvEkYZ9qvjkVJZsBPY6Fz3mwyS//G
IiLfpDxNhEXer1543OXcjQlaYA2CehQh2aSk9+UCsFtkXQz26dulujjnhylF0coJcbJKSRF0OfNP
X1SacyGCnLxspYGUDgdOEfuW98KEILWP/n4gWt8inxyKhLa13vpQLO+Ujgos783owp4ASrRx1UO2
GXtWceWFzCavdgreUJU9SBKVN4ksyI1/fmuRz7gI8fTkMYabHxqzuDZOMXAXQVFEwrzEbcCxlDl1
GkVHw/TncdRRLJfUKty6qMPgoR0YvMocaS0sY46y0DPFX2BCPbledGnLQtPcD+hIvqEkc0tL1FyT
RYraHL6v2lNk9Lc+7xdG7OkNkwmY0sKgk+zSMyg2eIMV7hKHCkDXt9yQ/K0w6u/Yv0W662gvTTk8
jwFacvoEoBgCZRIUValcx8kFWd4rydI+80fXwrrDIbax/y3+UWytIotrrNcsj3KobJmk3XNEIlx6
yTXjgeGr80QM+EqEV8vtKr20UUVKAB7XFmIZVQNnH0Fk4ZhFC03tbl9QhOcyJVayxYKAYFMFJYrE
bUHuODEmMKtzGeJogkjnEltpuJIjRjQvKN0BqLQEGE/sJ/q6x0Ra3213cveKYkDGKHvWP6IPLSig
Bn4qt2KsZ9nAqN+1NvKzVPgjWGG94cqifZdRHZgp/X1FR80KU6xcjNixbD8cI3Qs7Iqmj1klffEP
VFDNh/iGTpbYkRJKP9tBR2yKfXfXuvm2s5J9C/cBwWbNpjAerP+Wq8a7+hGrIBBItMxU+mUPNlrd
IDk3ohIRApuM9l7SSclVE3S9rioYj2smeqVDJLvs6a/Hdj06EIOYZlZaby6dd8qsA9Sgqs0A42BA
U8W54sWS7Mkh6B4ETzXXIPOoy5+mvSSns+vGxptf9/TfPW5dxmeyMFckQdtdvw9UXn/uGKYot9hq
5Ri9fQH1gEvlWn6Ol5ITI7dZN6KnZ005jLgFK98bdxxze+bX7Ru2dy27ISI5bjbuxEyd5Vzjy6L5
2XVjMa5rDyHlJ9H+TwKMGYMLylY9QN7XfTqryCxyN3YpZfWJU4plg9OOvAgS1vaJVN1fmBeAKVuW
At8BJRYaa6+N9b6/VpyVmvmPCMeOqMRRX6MiPz3yTiFcHHnAkl6EENKACBgj5ou00au1JB1wqtxM
2/QHNotv5x8uR3mAzHMpWcA89JjyEfX+qb65GKuzPjxk68hB/N9YJ2zXx/f0WfyiY4vhwdi3agQp
Tq+pxTD6KJx3RKuZlexco3UXn33w0m2jsuHqCow/9HMD91BqGmCn9moWeLZOBlF7X4U6DuUd5HQB
0Pmq57OmfjZSRzHD+WXfq/KsuncqRl4BfSQgwtUsJUcFCuqcBrR5CfYRx2xqQAXI1mEAiNZaz1/o
iEsdxe1wRfpiLW/gfwItxn2/KlJvPvKRbo8Hpier6PztZW8wsUwmq9ngoItOWpNgjpCbEbmZbFXo
1qsgBxr4t0q1Q427c2n5cgV+iu0aG3avvCLpx7FUdwJX1RGdJX+OBxicQ2Stm/iLYOO7V6HIDjL/
lOA8jUIiQqjUQyf1VEybrKPq6Na1+YC6noCSPUMkfxAyaTf/K1AqVhl9+ir4baB46aszCeTb8rAk
mEbg34uwSn+Xb2u8gSinB/iL3sQVMJvMPc+FJkujrkm7CFryYwMvB+OWnM2aST7t+XvV8MgY2LbZ
iW6T59UZaqCRN09fvjAL2lzBNCxRv4VRqiq31m9C13ORXpTac7He4YWEzkodP19vBZiNOU2fa7Cs
Zml6halaXqDHnrnYrlRADeRLwfph3OnWHuxMKEz7vdyyVOv30UWlF4QAPTsXA9T9S8a2XLNLNeoF
jR1ThJ3fRwpIqaZmV/+QefRQjlIJJES+taQ36Wjm5rMMBPCmnt/2xKIz8RrDw6HHkt1GZxMv5XVg
WgKNtr0nVs5kL2jvoFHSnX8Bf+wcVaU0mPSIUinE8+2PV8kx681WBeHhA94/Lcne/mDK8k2Hy27Y
0QWe8ioMS7VmRBELiwi/cidjeDn+IMPVb8tFJUuNXp6S1BoxOhe0ktw/7EXYZ9g/ZTSR2DGlmUfI
l5Rcg9QfP84CIulzRfLBADPdejro3xOuIqZjWxyIBewZOzOrBmjfuW652tELUyLtSgAi1Co3S0Sc
YlfjU00pWFU1fqMJCh3W8Em4qNoIQ7y4/O0kpkdYYSN7ugvyVy4TOaQk4OB9Bhxo1g59t894hN4T
A/Wj55vnRnvM6BNXEJDJkl3ehtuzru7P0LumKhhOqbbFD+dDWXmjghtwAmfpnmMbZngYalxF2dE2
IeiaGHqiv/3CtnlVd37/CcTRW7Zd+fZYFlW/R/q+9BD07dEBNxoCznaCGmSRe310vZQ7FxHFh1Sh
c/C848Ap5Ob2xdMFnhmlOmWcCU1qBumw1SJWRdmi/c6kKUvrmTPUrdIZke2JMCwEZp84gbEk7y5P
hmx7b6Z94WFtBZvMuUHb3fjp0ESXiwQvyDtmr6Xxw6HtgPlSPUtSPz0R9VWfZ30Cm3f7z9NIGgoa
wLZtQrtEgHYswAjthD+2PELFjgcq6wcHEmNHkSoCdlHk7/JCHecPNXa8p9of2JctseXmpc1QnYt2
7UV2H2J0cBwGDhqKMGYmkf0dZ9lt0XQcCXUsYytpNY0DUD6k1QBD1+4PQmceN6dq+IlNWLQbyheA
IE0ZuOK+J0sttsVCsNO9uRq5rhhlMV23PjEr0YGWf7Doxw0oi0MwD1D4danP/gynGm86Ro1TqeWP
Kg9Hjyy6Z06J4kty6PhVWnfCtwt90PUY2hiz8x6qbi6P+RZHy6f81Y7bB4APOma74xyWVMTS8fuV
hcHFs7lw+vDHTEPHtDWrN00VM32CMydUBWWYJ9MMYwz1A2mJsBiAcDIYoyRe8gtM5VlKxgKQObFP
ofzW9Zx+eANlFLuyYfo6xiFzF8QP6DshQP5F3CHqxUaAVorlp3tJhp7PhTfynxMUV5OVwAWXmVH+
9cnFfi0CmUhl4bzmFQW2BxOdpIbziGcU0UYttmJnGVh6Ogx4ZE20FF4hAUDBS/Anl3x/ldiF6Fu5
KfRrNX5C9J9J6nOFIQbMqFshxeckdFNzCwqXn09iL0auOT1V4/lcwyKqtWTKD+6SfHEJ/eyOZYx+
pmZ5MpmJIhEW9tMhfyfof9g7m8Kb2cwz7GUXYsLmb9XdTc8QZ824RVbwjE0Z9lZf7IiGCzrYMe9e
Y6d4e+D5osYP4Y30vXHHITyPmaUZF0P5WC1FcAxMFCVksybmX3v6IenxmRNkByoU6Gt0tPs0d7qf
GPwvvzckF4TsG8LxeHrHN6MUDBWw5dHXzqiKbf3J/Q+5/c/4rWI05YCWb/ooGfiFB0NRbq+hf5aM
JLqe6nt52LD/Jk/7sP1BD2tGE9Or6PiqxeXTAscNPUR6BSMfocK/1f+3S3d7+yG+CroecK6y0pef
ms+vgsua50E70xYzVp3Fx7MkE9Ww9zvS/QWdr4p9Gm4zP0rbe4ivCrhwrq+0AjuSUuQuGK6x4+EC
Pca99h1N7I+xzsAwkluCttPxRaL31UyCXajQHtdptM1J7OP+Y/TrWMkT2c1hfayzI+Clat/9faVF
NH/Tkk+RKoGq7/d+Uj0/Y9newfW8Qlfbk1BBVGiQDybPyTVWhcjFP25x2dVLLGpUT/trFO19JmSQ
+5cMNWu4KlG2AYPleN7BGShUTEg6gM07APX8XkF2Mz0E4CLi4agLKjoiMS15ooTaBPJuvH4iGjQA
LODORj3M4qH9NcwxU/b2N3q8dwqNWi5KDCUdNOc2BA0H8495uQjzpeeL6skbtEb8284OxZUUxfT8
pLMr7eUBQoO+1xRVlSq4Z3ZwdmfmTzwTCtZi5PUzYMLzi6nAINUun+V1TGk9MTcWzMdz2CQ/5jkj
KfZfhvNXeHq/Q10EQE6N2vfPD7C/tdePQA/jbgM39dd7gvkvzcZ/9bTjDnZD9fivZPxD8VvP5AX5
hQwx8egfOmaptlvrcCJZ2eOaeCFcsGDlmtERLEOoOKD4nHfoNjABPRo7s3lmOH7k3B01MSUmXsjd
wOG4S7KP1W2O2t6ZNiGo4EAqnC9Jwss/pBdLzUjhT6kAhLmXu1JM8djvqH7WcI1E2JcVJo43pqWp
RvqTY5sBU/P8RfpxJutBcJa+r8GMZoU/LOxtZBhkyqc/oRfA1mvfW6eeYUDZLLbh42qY05BNz3PK
exORgrkXCGqkbWgfiMYcMI8ch0tiknoMgVfo6hp6uq/sjrfHxHUEkgw2RNEecwlE6HhkC/gcNoXs
5WyQjyXuzWx6gpv6CrWmipN/Hjba2PpkY0uSCFzVrers51XqAWelBNnhvB6U2VNaeJ3Lw3ho1NIv
tKmGPgc9YZGb/Kl6ps1VLLahghh5Ed0sUuF8kQyqtGkiTSc1IhHJwbxba3I3G47jbyjLKSKg1hJ9
/ov7Bg2uRoNeRWuMOhgt40Fqdle7aPuZP5DXtLVKGU6gB8xqD+itAWYKr2AshmHGdFRLdggIW2V4
XrO8t/HcZeX02UnUX07hXDFYEIiYCM4F1CtFZr4N1O1E+72wYeb4nnsf78kzk52V6Rh1ztn21/na
APHgFh68NMPvEyM/LvRB9s5fwnGamjHpRGBi/iCJtZ0b2fxZloGee8bu5eEvttxE3ByHKdPCLus2
IAFGdK2ZRIZFAbhU7NBRSSoFeTk+YCBs8EIUTAmDMfZWf1/jCYR1wcazVKuGAlk9snxp61BisyXf
/4M+gTeVxBZqiKBKn0OzC0/6RVdxClN7L4Fq4ld9v1WRHWNn57bGYoPwC3ARjRyXYdk1ictZt921
hxkLLlT8yDrJJJrjozOQBD/ZqAQuCPT/rAXN2TdQNKn2lWksJm72d3zLh347v2l7aBOFrV6hhqeC
VcchIoGzGT7BkQXNk2PcpiKm+j3eJPoKK2OEP8BlPx4tGqBcppt1pI/GrqCUV0fcVIo156UGHn0U
RGvq+uKfBtXXd9GtWct5ZAxGsLEiWJDFPqBIlP2P+0dI5jJNRYsWgyqYM0NFE70Xxi57tlDBOyUH
qwMx4DTLwErY2/ARRTzBnLX3QtBvdRf+3Lu3tDWsic18QqD+NbmWKs2n3P55QrvXrdyfTsVTngJB
XOzHsEqpP66ODWzwagEQxMSZ8CuRnlOqjzOGKK5emnp/QwuKMd0bO+gHXfH4NZF/CUB+DHN2ooaR
CuhbEwyZdNmO3yuEDlhLXXFLG+/TKNW5LRwAfZHgLGZWbzgKC2JJxEeRd5G1ImlMvNLaK0yZ+2xZ
i9kGQ7W3noDnw0jzUyOrK+SJGt3gw70a1BDdqtdUcPJtm1bd+5m3Wl+1ED4mGbq8jIGJlEVOp/mg
0iyXVcCeqm/NDVUgpYmhTUNNcORb+IRoL4+fZSILAUJaQCbJaeHARMnSkuIip/9Xvss6sywtm7+s
ufJDJsSf+AhzpIWj1qzpa30Q//1rt4N39+ffcDY5J3PDvFcWk5skwhSw5yHgcoBVeHHDX49Rhk4J
yX/GkNNhMsIrdKquMEzB4ypEBmk2uCjl4O6KihqHFjEkvbtYditeAbQR77JMYW0VW1gzFrcjinIa
025AidSUTLjIbyarS+Mv8xQP/yNjgd3eySG6MyumI3kQNJKhl6rB8HXTFo9Z/GNLbcyOED0V7g9a
ZN0xBtVfMWvMGRAGSi05EMa0S861MCBvK8AEjId2xsHyDx0OtZzxzIHtv54msah7+jJhp5sBTy1p
WDCZoqUWZxFQLFO9TgIPywS1GIf+w7bcxYGX5ePLiDy3ax/XWwkLBwkBmiZJ/agpkOGqXNfxt5s4
QSG9xePhJ2HR1mbN0QoTGAYYtvpjkpzDunxV/fnZXGwfBPM2flUXR0mZmQnqm97eTQwsNj1bRzR3
JwDQZdYjfRMasvJZl567/4ClZCuB4UyyCcHmLlrH2bYa9B86jQnCfGCzQz4ffiNifEhD/G1E4Bdu
hJMtZ/y3ZFcYSXyCWVONtwYoBlpRoEG7vo8y02bGPieQAIIWS2hnK0GHL0jL4P6apE9yKKBJKDPE
DchbVHG/+pQfGpaJgjpg8rowl/8eiybRuxtHY0j69RD+eFBlZzi1QFZjn5Nm6iPw5hZZoP793sPH
zI8/bG2cJaaUFu4u3cWEO0v0o95jDNIGr1sxdpRSNvWARwU+0W4D4N/bP4HcS7p2gyM71Tv/BKAb
kYU0/215zd65WcvOB5DA+STrUMGLVzfOLAchUGskjWP44bIY9MFyK12M2nwNeak1rmqUvzGVv3XX
UTrgEMrBkbynq++rxPv9tSlpprLT2XpuB03Ok9Pp6JS08Be5f5uzY48SfrywxWypzr8kz+IlF6LU
wC3vahkjw2ptZyv6iWllr2VInECLd5t8E3jytjOeHgLdPeZXSxzB5la4DR4vRNcrLouqgjqp6ktM
D0kYdfG+H5/6LqPW74v2NNzkSnP2EJFS2tdslrl+u+arRmSTec8ypAH+ZFjBDyAf5nUwh5NV519r
hHsgb2Zj0kA7XI6xcJeEFiFnqIRaZzJ7zj/jqLhc3wpP5JxRqvqRCKLgRaxovy8SHixACbuMEuoR
E1lKZLzu9rlJO1Uz/rOVHkNIOyE1yn34qI7TOYT5ertQzbJY9T55eEq5/ykX9nKTaUqs6k+lfblU
WNutCKkjVN+JJDDBbVR/P6CzrV7sebSfesULW1awbwiG+2YHrr3ndTjyR54ShQ+wIRIKIEowzOR7
k743rq91wm3WigF7zfhQeZBQdCanWFj5/lknJmeFoe6sAY0/cFEyxq8RmkfblB7kayS+wMlSpA2+
WrOrCguG0KVT7DPOQQEkTmcXZzV3BdewHSPHUuAJ58NcbBsSFCkIKoNT9w3xBbdT4uJvijxCgAsx
V7wfKyDvuHyIquc+wZXSmq04rJzIxdhlu+gDVdoJmPssGKzERqEFKV7osnuLDqgkClmBSGpmwDcq
q92mcBPfFaobqbDxcR2WhrlCu46Jrci59l0c4dzugMYgB6SmRoRl1KFRpVxyr3PiLGIRtG1n6woJ
uyeckJoIaRO2dXg93xYc27SgXXqPf5lzAeLf1AA7Cfskqq0AcEw8OX96rSieO6ImPnbRLOg2eh+l
VhGec0DfGTqyhGuuZXqzsarLdvcJ6tryrBsRKU66UprgkfA89tOlmR6xZlf6/NQLUjtkRKLIUy6d
w6r3U7PrfwOZ26W/R7lrMYuSENStuuzGeteMponGYNrbq7kAv9SCDADi/6Wz56484Y12LDG29aPn
xBSksUuIL0XGNnME7pcAW046PrAt2PIFdmu1BkewoIz9tjdCXk7U/Yb0TXwsoMcWL6ZdtRcJcpy5
RpnrqnAQmk7A/r7c+6AyMTV1NQ9yDBzpvYNvQWsVd0ItsO1BC701mGXwY49wURW8xfGgygdGQCOk
fVdctBHEEWiSa9YZnUCtJQxo7373wsxZe0QjHobYlQ4Y2WOzrQV1LPAKQivXRKVl4JDsDkZwYnl6
xw0Nexgfu64VcpAB+D9PX1oA8hNHxZm5gRRrlQjoFCoiBmXp0NeR5gbDi3bSqlYZcrrqB/CUEO68
FDkijDtVKyJ+0S2vjOKVGmlFhXkkq8+IRTmveoAtmfDtkrhwfwpjisin//PPtRqBtU5ZdYdSshJV
s7qLlH7wLppVS4n5S5KIQzFaKQlCnDJ2e5x7WNjMfC8QCtAOOqoRa6hLVXxqEDhZSiYIYe3xixkp
3rtsYUb44KyfclHpxBQFuH5mYa1vB/PHGvwwC4J0T99CZxtHx1RLsXnDRMhi2A3joXMWVOIRRq0D
w/9GLIvAcv17bie61fwj2hvTCMlryaO3AqelUT5vJt79QBpS+uG5mNegjp3OPjynzOHHuvp6+pmf
3Zr8Mz5zJDBlFgFKlr//DV6dd8ZYxMKdPaaDy9SeAyMLvuKfZ7Mojt16N+5RSth/uhn39LawiUAb
LtduVU/vfuoeLf3oo8UIZfgcDD7eti45em66lUTqsxvdypTosV2ocJwPkALeHn8Uny1qnF6Ngq2X
O35Ykfj9Vw+VsoyXfUdtBenf2CqCKDTPIwyT6X2/gE53XJJ2A2uWUhHDTt4McJisJtwbhCxc3mFF
wNoKUi3/U08n/JnoCxcu0xH2hA9RX8Vbenx9NznCPST8IVi49P8pYTnDxIjnJhpmTZvNkewtflR7
CBfvRM+ezkjtIZ52O7Gl5H8O2PHH6ODS1LWoGyK/bkZakqUrCbcpf9jX/+AaxzLGrszH7KYuwlHW
jwPtWNNg2uswCP2Aq3YkQ2Q1O0dCwos01JLEBWTsjHH/HKYfbR4N901gLGDb13gG3kJA5QUobcpL
RvG9Tc7lHzdOgxsgeNWigpL+Iz+9441hEmMysYhN0i897wLbxtklyTSz+6E7/pZ4LF1iEr74kF92
5JxLkEk1W5EocVpXD7zWp0HcyPz/NVQXPHHrSwlWrELxMdM30cLv03U8+BOVNMy45Xvyb1Gg5txO
J2YpaCylxdYivqLh1CnvOzZGk9s3I+w3xyLh19fA042Wmbcf8hqn/OP58Hnk05BwsnZeyafKZsEE
zYiHv35N5yrr5oQ1RyYvvZyoJFhAnbzh/3fo6ZKu7KwOEnosdJ0DQROLZou3Yv0si2oxjfMUl1iM
iGhwZuDCFaaTNekfQqRg0AOM/fOMPXhBGBOiuo1Noh60vOczb75+qi0BJPsuOXWmntry0Bv6zcyA
S0SisUvTX+p5zDWkm4yUdEszvJmaUxze7tx0QRh661w2QcUF9TXVaAE69YUNFRc12zbao07gSe+m
9CUZWExToqw+3j2w6SsVgqCxaNgtBD7ROv/VikrTyZryof+da+nROZYZkXVYC1AsyHtkM4+34i5d
pLhzxv+CYk7hgog0d3pGsbV6HnCtKkzjJpOQs6l3GfjQxHHMe4N6guw3BQQJ6+PXEeE2gw0hfJ2Z
PeqYuyAHNgam5gAdgPXJmKi5JyVeTf3rXC0YxQ655XToz+iEOoQTEVqEWyy3V9CCEgCvyLuwrV+E
GylM5apb5dIUsehgTzVpTwJRSj6aEvA5ZV555wHjtTW6bR38vk9jt4FgW5DDzjV/ROIdSPW+0Xyf
3IjWtvKPAfVl7IiX+ae/pLlK8rux9mpVfPuqTse7W2PUOsd9PBe00YgH/2IiLx2iUJL/argTKtv2
JpjsVhwN8SgdkzhYiGRtMfmYwRUU5lnYRMZxKRH0sWUai25ibrSrAFeghzuuZZh7MlagUfFzFvX6
3M6gODIghS4lqLV62bypqmS0mqERc/aMtyb51VvxU2ffUtsJPI6hQHXjL7u1jQTQ6aL84hkEJ2QY
oL/V6iVfp00sXIq0/haw8Fx+1DcPLpua8k9jTGebFd8ppnABmYZEu2VpiJdIKzvsXrHIcuVTpx2I
OXx2slx8AJ3zJAM9bbFBPWCbZIss836/PYHPUUg+6a/6MXrJacXeUooWOUy/6lrY4jXU82ZlMhze
4pByEQ84tsS+gle1/ouhP0lOkNQUL3nMp7Hbo1N/v05nJLwZAz3EuUru4OU806NiEpTcja4hf/ag
bqONJoKm5hif+TE7lp56tUDAXx/3NLU0uXb36214Kt/btAjckfYz4bMfG6J/vKE2tFqcrl4V3rs7
KYAsBNQP/eAkl4vA/fg834+clW5sYhJKh1UZzJAt5HEpwh5QpGavkfqEhgADu/mzPeopv0ZH6LRQ
qKSJa0buv3Uy4iOku0kiopYxBPf4whl4UgjZBmfkdSk4YCrkvJSA/0ov/gn+xd1CTKI1Z5SN0Qiy
NERU3TgPMtvWM0VfHm58ZUGrsLq0EBoWuLGf9hpxQYVzgaU5L4MyTNA5XlSgEoiecxFpEzW+ExRJ
tzyKVoL3JhJhqORrrR16wsF4cqjHuBB7YEc03wfXlpkOsFXTiBkBguAFySXXn+f/WeZORUVpJUGB
5Qg/mj5nqUG06j2pCIOYfutdPFfN6emPPkRYszde8XHhy4lVXQ1gpXDAODcO89V+f4e9+hdsH6Bp
H84+6tNLp/u94VQEFrBBvtfzn2TTOvaUEPsnZyQH5u4sg84vFmEpcl71swdOVduhnbRjW064pHxX
xp4mMMKBNL59X4uI+NGYQDpG34NruaOXaUs3VlnOJGynGlPZHlZM0SMNvQpqqkLITJsy6bIHljAU
hTLNDxLzfb0+5nTenuzxJy47gmdQudgXArRAsc4/cuDex4hcHdMAuVu0Ckg9Rnm1dZV04z2hb0D1
zUWvnt7XBmMoLbnW1p3PL/uByWzb1gDSnkNsbE93u78R0Qo+Rh1A11h7K1+fc+WHDpq3Gr4IFoFu
5Rn5fD/IT8R2fV7HMt7w/OrqsUKaoR5/i/MEYwUf2TiBEz6JZdUySvvL9y7ACsPbhFIyhChoiw8s
dJH4NJxlYIhDc0DBkwyIkV4CScJOR0FBc1irLSlqlxPMiq0b7Ad5b1vH3xeawVLQ0Kn6PGgYtuYB
1mgQF7Huqsb5DutmbGjlm5A50wsqpfPdre4g1xIoYRMCMGdyxFsM0/OBBHYOLt5Wvy3CVP6T8Jh+
lXKVXe1BZUZoyfsATQlkS241Zwl45b6Sa2fXlbk6OrbHDxK8hRf9bh98yMPuo6nXKXlmkwEDKmVn
zT8Aouc793U3Kcy5qeMI2ZgGpmhpNUBb/nFVc3M4J8/VQsnRRebO2nBnNo0IWKmK8oWCXjF4pAu6
cI2MsOm5/nVQQyzafAW9jeRswllvmjLyag2S/DN8lLE4ltsJv3//JUwYhm2R0+SqL01D/B2ngnKF
rZhps0JlFTM8dDwM+ZcMpDhWNWc6ByWSGMM6a2Tsbt/wwmsTp8ldM22GZhsxNnJsHmY7U4oubIZN
Hkcoyzx3KVn9Qeut/BzUChjG/1MAEaJ9oKFDi7hJKh+QP560DrDqnaOY6+p4CA5f4cL5aGtN4wbM
V0Zllq7m2GKeJ5xNfwSMErwjEHy5PHVXtPgahO0qa5tjktOOfT56fTPPhYkHRPs8hYhV8Z7GBhAf
UGx0+G6NSKviQ2ZGIX7QTNhJWAqPTJDBgWZ/FoxuWjcMaPYcrYeUvcWbqqWpokUUBQv1m+HX+fz7
mOHFER+n8n3/ba5iDo91JXFy5NH2GDw+/67XJ+0QZQNKF+oSS+50XVyzR0d6u1DdNpz2CgiCBWO2
7KDxsv0v1bJRPb73y628n05UqiQ3ueY7zV6HMxJ4TqQVyYlZLg5dj6Wqc/iPNptyg5APyru5ab6/
QfMy561+KiVfwqlYnwYwVwCXPaZVmu9TmsIUwVieBgk0v8RejY+qoJYAxW+p7nC83qgU8bXnl5V2
hUa4VAr2Yas9l0ImtRnQLhaI3F2Gh6SI8CsO+ntbERCBYBBUAlXE42Fs10oTxbpYNQebqS6ZaN+I
SNgYQICXj0GdXNvRdPsUcRMpLlV+ptA9OzBUDa1h/GK518AVEJLlHASZR+hlBYjR9KJwO1x2+Xax
fokeYiUAGVkv/zaS8WJ4z6bATeDf3spXdtXwFq/+15iOuv95o+aptzAefXoQ1EOMBUnIvVo+H79e
Q2XNNRTIsZdNG2x/vBOxpgedbU829e5awwKTdGTVxlyKPnUF/SlnwuTbpGn9IEclbdGEeES7NZHU
jMp7rezRhpIVe6CcLKX1BvumIcN9PhUXNnGpsv9z7+I3zsp0ZyuFphGm2+powz46ZHOSSgxgaZZX
E+ngBRGV6QdBWWah6pc40a/A6tm78gXfR9YWN/XNqAofBXCNpqq6kHp8p2ilJmH+B8eyOK8S/xA+
EptBE/Hdd2i7We7o8IdjSDWXgwmxCebwEtVZucA77Plfofc92Y3UHkyQKqgJ6InUW4if3FVguyUa
Y7+q9Csws/0mIbr0vTS+nTe+EzTg5AwwDQGNNOQolBCyLd1zUTZ6Azc0dnSqlMJcleaLspAc/wCz
mw7E/G+SBTO2fjqzh4k4p556F6fGYfkah0hr/hSEJow/zYYdUyblxAekhuRC4JBDqnZMGH5cZXE3
AnNJW1tFAvesUJ/bW1u+gU1CseY+leMSgS+9/borRgTVWTJz3zrbdDzsVtEh41r70rGvI47DMx4z
sNtQadhugaO0LIir+/FWONQyIxr29ZxHcx0KniNrGr88d2kv0Dx4SuqRIGffG2iWiEaUDxLHO/7r
qNq0XjZjcDHJ4x0VGjWGodlkLTlya9PM+DU2LGQpadKW7DeDA8npAiVXdC3FHClgKuOfAlbqb2Qj
eh/O+5cITYNQ9r4LGw4oLoXWbfmXTfyjz31Fvo4u8r2XYUDsIbOb+UEhAPMNKlvB1Q+o1TNp1TAB
WiO+ICS8UEyhtX4YGFSOWC4TnHfGrFemkrM+NL96rvjRRNvdbPGYAGggU6vKpF6IE6jQux0EAEHY
mYnnV58opj9qNbSlt/6WffnLn3Y4PFymK4NUCzzlNWIhOVvvh0OMueP+JOx6KHK9TmyN7mLekkmd
DnCQhRIg84ZZ2gaH8SnCfTD2Tj/QekN99KY9eVDl5sWf0NwWFjmMS517Oi/PxB/HRb6DOgoGsQiq
mvho5s+zjrIyl9v9GrfnBrk7I6pmISEueweS5ESIqaWKxsyzCgXADWNPpOBVcsL87ssGfwUn6fL3
gG/5Wf4kuCtHgLWVNJOjxl3FEgF28u+c+AVzSusH4plnigc1H6sJEnSKYXmy5IlBMKipnVWiTrKx
nR5837Q4+faywfzNf+iwaK81DAdBrTgs28eHjgE04HvjrZbeNwvYuIBvp2oVnutMsNFD8FSN0sWU
V2/Yf+7S3Ty7AwD3EQRf17bgAwYmXCxRnRKVjRvD7/FNTx3rJoNc8eXUXiZXzf0vOp/HpFloitTN
Chtkhrrijlh8F4nejMfBw043zc4tUypTb+6V11finsod06vXQEfHOu9qt4zXZS4irqMBoLmAxlwb
FOZ6Zya+mSwy/pPKRyoQeacKLeO7QqoJzuKPROy504YqCE4GjXIHbrtmjA1JXHn1ZELtatJV4YzT
FAiev3m+/7Cy9TQHzaJW6O/sd4TzkHpRmtzBsoTB/EPubbIbmjsktuviOc0A8kwCHb7nxqKiuhgY
ygw9IieaqeqO3wnUPkeoRx1uCBAkHqXP1v/Q8iE+a90da2hDJKdDRRgTrUoLiHdlXci3+LToOsh1
CAzrHKbfVxP/Rq6lk7H0/LQE8NZa7iCz241arYPTLTz0NVBDtpMxFdD+yfPtGROYzHijOaU4dLUn
K29LEr7LgvwxtDNjuFHemxjGKuCw6jLZvunJrug/iZKK//H3b8dCoTGKKn2mEgzCY4XGKS3nztN7
cJMr6IG67IdxmJH+YoXd7P2bM+QxxXSDPcXf4gbhZpt1I0oDmcnKC4XNPIaypjpAWxuV6iDaDfHF
RNOTnb6HqhBUfgBawmlPZU/F65nTKYMRbWjpIvryEc92QGWC/t0vPyfeTYR9S4wq7TbA6TDSlWiq
gTV/8p/i7c5VIMt8dDg154Aj/u6Hbt/DszNsGqxRZO7Z+ykQUiiIt209XZ0XhAtI85cPdqVo4NMg
irfxzfOtmFHbZjOy+9WKs9ZAcpCocjCHu6vXaI5aPq/oys52GnckhpueMOICeeKrWuNqCUrzoEfx
FkO485P51i1lA4o9WXm37l5FRceGHTD4OViKYCdA7yyCTqgDgcGLRvRV7fBQ/YhFrzYeKlOMlW1w
acyyVr+N+PSrYkU53YRIP35qLZEHFjIRHAWirOtKmqZER4xhEGcyFDDYQOEGG+6/avUwMnbqXGaB
jLfZAWipPWpZdZWWWPsI73cQv8CUuI7lTEn7TaHHqx115mJur4FFwX22begdnXRtRzvbe8H2/k8I
gSYwKrWc7VKAeIuDrvx5Mbl1OC6Q+2lIyABpyrLH5YNVTYnxkwiGzcgrYJJ9k28YR4120AszxGc3
bFBbEQcv5y3lX6jdFjx4syz4TXaL+ur5AFKxVRzxk9Jxzdo/HC13Rg52apEzBSHMfZuTuANrcaJ4
Bft+T2Mh5Jg4Fd8V/7OvFZLTGkEqr787Ae+Gg7BryTmvhdTi0Pwpg7PZS0mn5j90Vvm2BYTHlHTk
zXd9u8n1SxhdA5037g4gr78xMM2BwkUf/UQjSspGPm1p7COZqlfbBtCvDCnIHmrldljFP+DQq0S3
TLhxHdT68u+9BzzUTHL4kM0KoUicbtekeIGTcg4M9L9IsAyT90bQmAahPLB18aYphm+fZCdMMm/R
Vgt+xovIrs0bcwRyWsQRBKxJuNJ3jdq1NlN4KDqrt2u9HH+iDfD2ptQV6gOLacSsHmKYIbxyeV0w
4QngpPEaFI0LLvSDTbaimqhUrGx1S1QnPa8SqB+uVxyMmXkB/tyToDbDwOAwg1YV30RCBAvjZW/6
ZRZBe+11+Pjf21hw9B0ucuEnwmILjlo/B+6nF6HNh8fpO8Zn7UBNwFac95v9fXA2GWkIHY4a3aU8
NbIgfW433dxRqHZFjonNNboJ4fE+MnSTEVlI5u9BhmssJ8OMjSTo6np8pQ5Quhv/52qN1lam/qXb
TWs0g/71iqt/pS17Agj/cZkKNLVo9vMHQlTO2e0mAA2g1l+fphDSG9YoNow4WXZYVKzsUgzQlBeo
fnX0dxuzobCweYsf50W+hc8lPOkQczGA8ypWrxz/Bj7hQNaN9cZr3BB1sT2NKVchXYaB3nVi+uYT
xjzcsSQcKLqU2UEewjG5iNk3tvhaYY4O6tD4wBHLoQ/FtIYsXLjVW01yoF7FDL4R2FcifPl4qIQ0
iidhNB6z+Qa4kho3fIiU+NxgSxgjWqcZkOccO0m0QtJ6YxM0xsW5OkiEobL6pJDgoD9IKg4I2Pg7
UCm9RdQmMSt404jO0dUZFTxAJgmoeCaDDiHSvQzq05HSXAv8GbwoGb4RTP7epJMusTNrbP5BDUlq
BNR/smPjGE/45aLP9KbijSHg/oQ3gKO8DiqRhJFloFfG1aMh+QY/gvIFFUHhtoBXzD8KxsWZXXcj
I3dQhsxt8bNaXees92qxsw0eWsnKQCTMUMPxykOkCsSs6RLQ3MCNb5KBuB7kAgFANv7NF7DAb0iY
Ygwg4WWwZbB+8O8lMQbu+LqA6UZd2dHj7C9cMIO9ke5ng4R7Oy6ZouCHFgHSAcEM7ZzHFiXwmgUx
mab3OuhR2/LjLZ4WqUK3BGa9G2TfjhQvHSFphXzpqUd5VtyZSMbGBt3lWNspziBr1Q+WrCvNGrll
OGNcmPzgUaYNMB472LzYq93JeK7s1UhSWlVLt2oV49EN1ylVAl2guEprvz7dubnBUQ7ZzjkhVYyC
YKPP5gSexJ6ZzKDknEKvMzS/zzQdkODXDeno26d70lA3X1sTYqf+48fIFacoXd9tVF7JsCSDkmCJ
JNAiyw//SB5tiINVg3lPiekPARCvUftos+nlyZr/rJ1WWnCbj6K4QECHOGOP8IptxpEBssLydR5i
OmP4t81aD16gwzvKPO9aR8TOHi2G1JT1tTEimfJzpNQTfATvjpsc4lOSmguDZaKVHOJg+f9mFs1g
OQfy488Zk1gECWoxselmrm59JjgMGigu0Z4TYcaqrhCM6esm4knq2lThfcQfLk8t+bavRyV4nDAk
kgkHJ9sEEVdytUlD6KLf1nzooOBxggJk61stY25WEpbK39feMeAfXj6ZYIcF4A2M7PcEBHni/H8k
1tX+2ml+ejYOvz3pyNQUBN+J5uKJdUD2t9F4X6Dh+n96/iN+G9y/est/GyPYUsmujjnLOh7TjfFJ
RQMCeW6m2XRYSyPRpr29BM3t63178nLTPRl0v6MbFFcwOgH4U73ivmmWJly9e4z5feoiHKa9BCaB
Id8IVQ6T7gZ4JAL8W/CA6ldmxz/uYi2SocFJmbNQhnfgzNOTameUQtZi4Sw3wZGCInh2N9Sxs6d/
ufVLy1hULMiJsJZuQ377lg0lOfL0LgY37me0/d1ru9SsKVpnS5TjIWEIfgD2iQAwkAKheNwKq2Dy
hf0sfRsjAbT0M+fMxlmgJU/3jBMyzFQOr6UKOsov2rBWC3IUr+9CYYM5ure8toxF9sunxctlhf9c
XScY2Or6MKbUbr6uu05RZn92drTVoKWGLvb7GPreIZXgTlDZKMbPUQTih1HFKRZbSmZI+rbMyA3b
rv8OMshneSzWIutnmp4fFE8ZhOx5LmDS7xhxsEA2fNxJX04q8Fenyq042GJQ7jjuI838b/C+PQCM
O7aU/atlsXEn2pcRxKDiZAofEQql129t+vMkDAQhRViTXzscj2vRusbwEiCV/uxPtLpY96GjxEeL
uyPC7wAnsm1oGEmx2uatz6gMexQRcaZhtiaCwjL6mT4K+wfy/4c6Ao4R5p6XYEM9YGP3QeUf5Ebp
Ka2No/QDgN2uaOWoXJC8AD0f1CsDjr7iNSZAcX9EpzBzDJ2F/udhs1FHa6G64d+dpUoDIiZuech1
TJKE53DwSs3VTTLqUkHtqhXULJJT50qGKztHUJd4PVsMYNei+VUPHO/cAREiqQOLz5dULMkln1aP
YsK/wDp7guHFw3J/Lxsqz9Q/WKkkDa9pk090o8ecDfdmoMUg6QGuO4xogqGzixe4ZpcJ6XCjEfuq
Jg2RA+bYk/+Z9eYoXbvvvyrZw8zEfq5tNM6kXuRqupJfYFGSKHyiojlSgWZeQX5Lphlyjvgn9Qn7
T9/xlrbmzcP7feq+BfRP3ANX7rUDrKbTgF+t4x0EECfJrzPQJz+AFzt2M62QobgnTTvlTGQK2G8l
6K4JKy2sbn9iO63QE8FtWR4g+QbGqrX9WDZ/CyKKQ1WUhD6ay22bsmEwY00kObcRzWf1C8WVDyW2
OAvY7W/ZOnd+BzhLNVQslyBgYMDKxe7y2KAiBA6gofds4i4HeYOyWT3D8cjlgHdnCsUNJ48lfbQQ
YCcN/w/39oNaNZeHx27wZzGjuiz/0LKY1kBuG+kCM5G9db5pg9PfpJs7DDJcA3WpEpXXFXZ0/lPE
gWhWDh0hnmV/r3BayidGyYf6fGI1NR9aSaSLGfdMa9In2/rhQHE2MRVAZvS/qPas/RwuArw3Cru1
wxyHy8GpAu2MS8oJ4sC4p8du6zBMNesppVf0zHTI7NWUNY0Iz7+ELltef59TakIKxbLD5laoUYT6
VuuL7Ry7aDeNxPIL0cUkRS29gCgpoJu8J9lmepREiHGKYKK58BRHnXF+aF+ZLtqzWrPMAT5CgGgB
Fll9+rC8A2vmT+gSKzr3gbpzmrj+GIUILpAXjhK318Cu0ul1AIuqG3wzaUi8CNYUEdLnpFXZn3T3
DeakGNfjJz9sUaJ8WewPRIUYPXrE5IPqQSffqe7I1dJcGHRAyikJOJyVXuwxQgAVjIVMVTxPZmSU
2ZCVSc8wXf5Wi+/KG3ZtJoow20pw/xpOiKafRtLR3wQ572w9hQw9/oLwYhdicp3+qIdziQZ05aww
UBJFbV4S6JVHNWk44h9O4sEs5bpUEUX6fiHDZiVx/aYsL0coNEfUzsxQ8h0E87D+qLh9DrHBHivz
2LWHMY1N+AijXomAB+7XbbAWzHnCWLV/5pisS4H5DBtKpyfNCM8lI6DEg2uMnT0yeVic13Zzcwgq
EmicY2o3MBrZoGrmbov2QL26NVvq4fI1FGG+4B3BF8//te1XBi0nyzyMUlexTBXxP+WC6yWF8hoa
+hsEfiR2G8o8PhcAQS7TooZ8mGcoaybHfynld1lqrjSn8K0u7kczR6/pd1fApOK7j1VJEo0p0rv8
d6Q7GPq1gCcbSDqzTFNpG+TYmlbQyDPsEyGtLNY7xcbMCrvU+Q2+h9Og9fK1p3Qn7qZJlplyW5vh
WgCyavies57PxNAfKZglxf9peW77NrFo22CEePbs3NOiryUD8k0BetxghiWUfQCl9GZyOZDcFCER
6QqKtrJuwlXyBFn8x6zSgqPRr/qmd+Cxv9L6Zy0ME98oX023i4S5Wiwct3wqgW2RIWr9j2gs/QgO
1oWBRcNKyhIKrIyvKOc7IjYUZnd6p5S/4OytqiiChaj6Crif3DckC5agF2iLGuBW4qGM4BRahc2q
pXmbiF6D0qbEPqQBsK6VfzaHOgkgd+MIail2l6XygAgQeQzmey26dPix3SiWpRL2JUaRyIGXIBV+
CvjisbTMwIhH3DSDSkSlK+gVRQRpVZYq+1g8fokYirpREdU4MIS7DrnVkSMcdPJz+voghAxFofkz
yQeb4BByv2cWkRF2bs4AxVHqaudkTbtSWbwpVWipATpGMrxxbYY0p0JBPEXQ6OWED/Ggyit/Thjt
FKAx54YDWZAYVVBtkXVv8N9LR8Y7McrMLX6D23pe96LdHY+o+odo7ovkQoUPCZQURKV2Mc5jUOwU
dD28+sCsNmzAqCICt5u8JEbOO7FrqZS2dqoCuBvcJcTQltn1t4W0c2iDuWM2DQOWKLFJnnjuH9h2
QIrZ/iKW1FeCxRmhZ1FkEwWp32q/sjXskq5jjDdUbXMDgY92ARoHN063oNxFnD8inhf8PM3ycSh8
fyNhKs87OY4eBXXlKUMqAVenYWGt+q6/2WSVrJLwDYbltFtRvR5nVbeLsvAqyJSJALuxguE3Afq4
SJ42lTj/F7fUF6qWDX9vKhZxfdblgcYrva4IkJ2ckE4uv5uRZkBEruyeKjRfAnYV69A/5PqVfT/g
BLc9DcJqGT2bSDPEAuO5AzvxqP6UO5C17HdWqhy/pfDhjqpfwcT70VgwL8ZMR8mD/Gihnn5ZAMCM
28HJqrpET/5CA4H+yHq/h0VRDinkgQweB86DZhje0UgNcZA6KH2TGj6yIiTaxI4kN+QtncA1vKd3
oLJ5vH5lDIsq5StWC+5/csPPx4VnUkRj2X75TWay/OsS3eEVeiMU7QB8w9m6RGPkV55bNQCvJJuO
56UI2PbjP6Sgxhk1eGCqwoPXd5LhDwF3qA2I4PqTTyz6TkooMSpv7/j5pHMQPcL3SKRrquL6aeS3
1p0V6A5tANdlUz02RgjsoNeNLfHOJ2JdRNr+voGsoYiMD8DNOkKy/iL2t4GRwrkWprn9m0+eFiNA
1RIx1L7S5IvQD13uaL21wBAp2/BdMTX90OYgu4APXWPU+m1ItrqG5/dSgp8YfjANGQvYCMSfazoB
KfrMPVkCilfObpD3xLnUf7sFmiYQWI+PknlmmuDkWGYh+BjSVa47FxH8i3RPmOiccKYYNfxYXIeE
4qzLUbVkIH+1OKIDJ9aApLpS7G6LgyUTtBKcy9k9Bna4VgIY9QOOnWutHVYaM6qFxZHSGdLd4j6z
HoAAyKha/gKrt0rhmXKbtZ7KspJgOPlUgWQZukY3G6MlAxoJjfVfO7jySjHuXamlyBPKGWR21l5G
Olk9XGQsCCUjcW7KvoaLGrCYdvOZj2QU9T3Fvtxv5Qt/22hgdQOvKmvUIjOaIEdkAukPLLoQPwC+
MNXI4pRyJjQhvmZVxhoRMwudsh+wXhTGj8c9sVfJ7GTIKasm3BDjgTM0kJoDZOn8SZWFhrJTknVW
jRFut9VKSao3OVIIuZxg7KN9Om5tUJudP+GlBT8xhJmvNoxunqz0DdsFg0C+pxBuxeSfcbYWesO4
3qHD9Ffl/bAh0vtj0Sh7Zt5lZbytc9oSEMXFLOI9SRfL4iJuQI5h8J8T9BEXt6M9LbO/i85DrSFe
wBZFKiVZMPAmMjwMoLfhDJPiCBrCh3ek8xdZvEix9OZBe6y+vunuosxA8Rdx1NuSC4tn+mJhE/gn
3D5Gs1HbAufB4xglYdK4Uk1MK2iRChRPEFihs606iYGTHlZDIeElCYak9N6meqj7L1+9gHGT2Qr1
r/LuxJqUHL25FvUxb8XcI8q5dM0yDzF/CL5Jvk3FhtieT+MduFSMBpc8HTSWmwbOcvw70+WJRKFZ
dq1r4+/IACy1B2UX2a/Qb/iQj+4EYA9x9GxuTjQs7taej5iohtePPCxr7ykIiztP0XHzfgOCyvzv
GbW+vHYR6XDgPgwCEt0RR6c4TLbMqLHT0IYUfCykzVn3q6i2d4hieyY2dZXe+BRTCfzu5DWOlyMQ
Ahh5P0+mH92esxBbs300WIeNAac1CisGTNrJqrrqJpkEiwI/UY+L4c8Xks/PSc7wJmKwAjsULe/t
J4as7A3gCEQ1bex54TFqAJxCR+hQj1OX7P17O/sOOdKKOPeL/MI2jg2IvimFw7aM3vmUHg65eCOt
QHMloogLXIDYChc5qEYDvuloivpMDJ8yVxvbgPSp77H1ZUFKsYswLDqHtS0mhAjxvjdYLYsqinhh
1qJNx7Wvgg7RU0nOYKB9R/bdjAADxKMKIm75NStdB3jGUiqEznNiBh8++YCquWfbOZuwhCMnUPW2
SFTwtU1zErDrTRoGkKsObiiDIUhRmUcwST/A/97cGWlT9bUacs/tDFqF/5iNBHRXlGLyBmMVwH+N
SCE5ATd7Smb8TtXC2EnVAHSHuLjKTbquqCGq51qsQQrlJt6kIoiYmeA8hWS0Ox7r6KorJsozHDiB
lxWgo5BvhYR0OgphDdXUAsvkf/pEbCXJoi4sGk/gz4bONCXpP4VuJVAsHuyBYStuhubIeuDG8i4W
rqIetXlhivS2yMNKKptYr3+pDQcefiQG9X0PrRl9iMwRkQF4uZFIlk27ccNUZ/0kdWzD4krtced5
TxIPr3DV3QGCcgjpTDgDE4Hd5ygslOWS10SFCyn7Xj10Jaa+zlHIJkqgo/zHEcrjRupr2U2Jb4Ww
PwsT6mqAukzv+qMy57EYS/zixw8wH5o0Odr30um/Hr383RRDmLxAFu/SPxQ0/Ih9ONUjj5SiKoqK
4bE+kgquAvYXlynuqgrrh65EhfNWp2vGapFDrW8zN7aLRXNs3byXZHCpgfc+AjQevFzYXNuxnUJM
COBo05R/jkyWsR2ydr+cJzqfp5wLtRbgB4Iz+6UQFhOtpLecTzYblRH0xHxacJf4QNv4C9MwuHpf
Mon7/gW5Ba1ykUvxSVP2pjGxeQCAA0thuuJdctAs8CfeFRNUNx9z3TSfh/PZ6qpSDQi3ssHMSCGK
ObB6gjm6h7ru2qfQFozBUxdfsKLC3PcO353wVwoxTAtP37unN4/15dmNkbSQdIxC8XSAC3C8PLc7
sBJEKaooLxVx62acw87pC4zrs7iRxab4DryPOMhPObxQnYuXqyov4mQxc7tNhN4AHvRnnub3xRwM
3erYvBJVJm2Vg4VcGGPeyPiFtkFmgr7OyXbNs7DEOWP7DukdHMvfPcP2V3/W0TaHXT1KXSepSbKt
OdocdFFB1pAKoQykbdtCqzyctpIw1yk9j3qgjQ1ZNY0T0dYxc4EWDCUxfM6PX6fp/At65+rl/5AV
TFkvtR12f0fYom+DjBZi2n5ketQJave9Ql7ObRb9VFJJmEAXcdOxtmwf19YU6y8b/Y2+xln+mWSd
CYVtvIWLV4ABksdXK0yRmqsR3Oar9a3bZPUAZQwyUU+IHJb5FMfGSQtEJqdFdI6OZaUiVREijewu
fFpBXPeOom/7E3evmk3kim88KN1pTgFsHOWONn4sj/Aqluh9wTXYtLOLMT5fe8FY0/cdEc2HZmm+
ojuQw/AvVC8lWC5sphoGHlbrrJlBZXE5LDmKATS4NC9IsRCrvoe4bzvRWF3uqMWmD617Wrlx5iDN
OKtxqnC/JLX1bvWOL9vfBese4H7OLywTQjs+y7D7yaUzfBLonSmSnBrXkhTF5bst/xWCwPefc34P
KYg+TP9eQPf5bRC45e0lRq9zVCmINq9P/Rs1yK6ps1UcHWGS4yb/CEJ3Qd/yTu9pZ2ab4rR1se8W
57ySZtl2S0fa/xBxkFck3GVXCknAHj2FuO8foPioRW5rerpA+QDNqUGaNRxzXF88M7ABLeLm0c3O
7mr8VAh0Ur8+eaLnSuz3C4oe9eTv9tdeLCu7p4hmVaYLUvMZ10N6CqdceG790CKPbqpZU+syVqdp
e7AWMIvYgLJxOGjL/A2GjprFyd1wlZx2N3+FuDD+m+7VnTZqKWdRbaDQzOFtRiIaZwSIsCfDfNxR
MG8q2ZSVNgBXdF7YN/jYSEQK3hyFCXbLGqw50bHlXK62kUcXXcgTrXpcbpfL/gFaCM08D+pZA+yd
rxT5/63xBpaHAXuk5p8LytUBchUQgx8goothV/FTdtwPEhk3zBPRYFUvrkmSteJ6okZA3YwnEktW
MY1OX9sNLxTsT9Do08hPRqhDxPbQfM08d5WMIcngz83LOehTf+RTJKUxwJKcgrKvXQ6ZP/v90KG3
+aWg8hnoT+c4YyztwVYimA6OnvJrHMpyaCa/Qr5eAtbnGdvCnmhDUQVEpHwetK28xMpl98yjhi05
JucaBNN8E2XjW4LchgCcgBYmWTb/4nNaENx7X2v7HV/uJQaLMKg7FZWT5dsQORd2aEk13Gr9hw/o
mh8eMV9t29/D1Xa+dEy15Q9FUvA9wfn/cE7LKHrMJkpgjp9E8BOnuh+arIj+dQ9DV4izjRs9eEOR
BLub11ZVy45iDOtrQk7ZxWz+8yhJDj7Oy5wduXomfDBrTzIfDjhMaVGKEKJYSDboc6o0t1uckqqJ
njJfpnl8nqwjEcWW4Tbc0i2bF70Vyn0+LVqTSwNH+OQummq1gSbAdT2J/eiPjS+i0yaImRlmajKd
uY10CoRlaQsex/FMgDdj45/BbOyyXvY4bFM2vbbj2puCO2uxAedq/qWX5H7QPxJrjQUzGpDUHbZP
qsRmI2miJ2ILR5p//fvxUoFLucLOXvf4PFRIB97/XQGdC9aL+skVVnAJfz38Z33DYt8VqbNFlHij
96CBmpbyLrry2YHXyWRqZZDgudp0GqtEmRYbhLCVivLJtxEJStaOZNYRddSIp2meXBe3V56uK7XB
77mmkrzcFZIUBslBaGPX51vd9vwH10b+T46ttJvIq8ddWs6I36NnulU7qjiwkT66Wk9OCITr8wuQ
wYNbLFl96YHLABFYUKqRonl+J0vqPRdytiZQB/dbmsvbDDMMnrj9lXf33ET2SJxQtLIQUmUEhdcz
rsGn6jWpUhKejHOKFD/yF1p5WD8iMlL6z5loi+qKAriZH7SR+TxBObx9IG9qRt0/3Uq4B08DApKn
7qCkXSXYP+rcjavwcv5tRBtSWvva3n5Ru+xVbYwMB+nUrtv7BtqXctyEGipJjAOTqMo9nzL9FzVg
S/mTR4x5OWY0snya2jbY9ZUvef3si5HC4AZtHoTMukiBLZvBnqzxyXiirj2V5lTTPownIVK3c/yl
KMVLC7wiiBxkyoAnp7cJB86KZzlaBqVXLlHhytwlPQm+lfyI/G4ldT7g0EYzBmNP5+kVW7wSM4md
O6AxZ7oPSEsbbrONjXCpvpf2FF9GtBiTcP6x78+HhHojKCQwDJ36lcbX05442ZcS2yJumggkOZoc
exM0I/A6VoT6C8eC8l6eja0hXZ26kiMaK1K8X3GLbgAQfylo79fGPPsFJOMSEtUW4+mRHKe84aG3
TE4eGY6HKf6OsdPoS5XYB88XTZ3eqS84E4kmcV0p7bf+Eu2k/VZ8O6YddLf13GHqjr9fTg04Vfkq
0ajIr0IIZlmmMUbjZZ6NVUx+JuaI+FE2lhuLykBaISDauAZmXrK3+SVSfr3uq8v9HB0Kog3rQLjY
C2mDgQg0iN8Lk5jlnFZCxrVxFd3UysZxKc/rMgp7Xwb5MZWszitCGDt0uBlteX0BFWA8LKuw0bZ+
0z0eyhOpVtwGtXs/Ojse5vNFnimH2MOdC8sNMT50oGIYK9DdWCtPWxWCArD098TIxtn25Lh55PwD
ro0k22u1vD4sjMylYie5Iq/C66dDvzBQI9Oht+e2oQjI7QQcKr+FlPqwrTwgJWNRTm0w58AFwX1r
a/VbeHCPPsfJ+uuR3hiAnUqH7MzgRWsSHj2xQMnBzMCt1aCNStjFKim+W/GuKP6+g9Bf+kELd7ee
bEUDQXfUJsiuNzK5O+DjS69ZI4QaprzhqU0d1FDTcK+h0F+w0vCR4ZFiyv9sLVVB2AJWeSgDrKBR
dPNdfv0OagK59TZVIye7f9Gzp2RL3SwfjneWEwIITnDlwlxp0yZtP3pE39GP1YfqYipr8exJjmpx
7O665NzAI2I6VVhluHBrkh5zLDfkjN39tvqPBZR5ocVWT0dkEU0bl9+vLg/3d4zjwkFKg5quEOky
oPsLGnCiwHaZLZM4xVQ8KkQq+r2wTqcfJIc8NwRcxkFT2GZzRel2dejJGLY0rNA7AtA+XUkeaUj1
f5lOUfk4t4N6vfJw6FuSuUShvejrVAdWxOdwqFWe/MJLRbxoPRLgdf7gIxNctjRC2s9SERlDVZbp
iWE0jZBKpubJo1GtBzyDXoySuT0LC5kKhLhSM0dg/D3RlrzE/ToqEKqmnviWkTYzFmSi/nseZhoq
ByvYkpagPI+25NtszktHCx4zyzQmhLcK36GCavYH5vXHtGD4E3MQuM1EivX859CZh7g1qtqIu9oA
j3LMPJuLT8SAu3miS0uY2BHzSrcOC9au7KFM3Ot+JpRwDynQd6eOScoYOlL95ZOXRRdh2fM78OfJ
gHA3EWp+QFtZamlZBx80ivgzByZRFUntHE8a+6MoOCzrsO4xHOy2RAAh92wosrectWQ9+77ZROdv
zRXCWbWFoTTD5AnABnb0sSswuD5ZARmyik+5JFUzd6SisRHG7pdLsv9aXD+zR89t31wiJV5KizRN
XH0o7Q6r7zUt8rJnHDJW3kE8fe6m648wgsCEtM43BYdIY3lZAhozD5fT/JqKfqz57gcI3yzx2hXl
uDQ12ZejVHRLmddwQJg0wf/n0S4xfDCJOJER3buKjOBW7EUe36EnQQtTi6gslMA7oA5BJozwJxIW
qMi0VMU8hDrK7vCxWso4D+qZWWcpKNjAyP57A+VqM3EqC9KIDqv9/E/VwPXJtXBdrzCBWcsrMSkN
KH3ypOT9tSk/liODmdSl3Vaeu9Txk4DC7SbT8IHhJHLlSY+ZI1jrcPI6OtFv1cdrkyeZ+Mw5fM6q
/HRJcFW5TX0ofsLnCNAkldAsYdp0TZSl3J8ufVfXIY25je0V2py+/NzaGSwpX5XPll+8Bx/ZqdMO
OBEnkWPltIQHCAawWPEyzYNv8y22vIilbfQ/cYZVaOwg47XcPOxO32COtbABRBpROBqKKLSAUQJU
uAeIlvyGZMghBPpu6HdQCf0UYxnOEW1Z6eNKYhuz6WV6Ix7fjhLLoSnPHA56qjuwADL0EdW7yQJW
YVaPUjMwI8fafgS4r4rS1FxUXh0XK5oiMYkm8S/4NU5E5v2i+Gonql+W0S9Vrji5QNuSeJoAsF1T
+Mnkrfz7vO5XHeZljr51i/ZriCc0N1fklUde3mvwOKfGn1THM7qn3eFbnt2HkH6maYoOg1SNV4lr
/1xTnqJtrh7vXZ9wZuJ+5kdsnNQLHokGwDo69zwL70VPerVLTqhyBM2b5NB7DqTD5hcY3pAOfSOq
W7UhZSSZ0mcm/p1WVWa+Mh4JatmybLUTExw9/VfJPfKgJ7KP1GPEqQnMeeGYA3xZIk9N4Sepfl1I
aKan9WKv0Q6A0i62qBCW7fbhm488B8qFxccOJQ1WCyMHUCOecT5+NEdC1eYJPaJxjbNCPx26x8T+
qxWA+tib3KlAKnSARbxjZ+mKU6OGSHZmDHJUoa9RzIO0YEs277Hzy2NWMsDN0EwEG6HcWTd7xIET
jTkAyPCDKX2uSRYTnKecsUXbF9YRj4MlfhW6ShyzfIyQLRfkzlO6l7ceik1vAwepQm+N7TRUmGwe
9RVJndbml/e+6hMTOSmQWy1QjSX4gMtQOqI9F7+pYhf0fSU58eAYPGO8RKoRXzrLmKrnUIffNs2V
rBhhmaI8T4RpUpSdeUdb8k3ARBf3zwJM/qS7jpTzFZTBC5/NVx0AaRJhc32Q3Budj1QEZK+ExZkv
61uZS/OBmFeJQ+s5jXPPnw41AEIwiK056K29BtwvNu8BdYW55Aj3xkM/nI1LKmAex4dZeijML59b
oEb0Gf4gc1mUxZQDQpuAje/HrHoiqgw3qEOBu05tQdXoKYxtve81GEb6PYBo9MVhgWs5CrhnAWYs
qUciqi9iyUtRytodxRYsug132hYVRQztqJ+i0pKwV5/+jqfzh1dj5ZwGHqLnqbC12Kj1ibU2DCU8
AJpGZyyHA+f10A5wEWa42GqgJpEbHjT9aVycywmWbB90cpMocqrcRfNi+32Scprk7IlBT9PkEdn5
HCqGx02ZNHsOubzUnJccTqxuJBOFyK4ekJ9Nqgotl1yu0GxiEUEhkZtO7MgCKFWiczSeHcIoVHEh
ePezDQn3LqILLBNmfNmQdwtg/+ITxBX9HE3iRKX3WiOyMIBeh2SBl64TjwKlpzF4BBlx5VCt2SVc
0v4ts1Ut2eh9rxT9DzBZQ3Qcu90uqhYmDp9f3p/esPF9070Asywrwt5FzmB1afigZFcZNU+o8Onz
2FpETi7hQsYhaikPCTCZLeRNUZnVWdZ/smzEpATvnoOsmAWDEezyTF90R0kyjZgeQwHC9m+YR2Ys
kY+ffbIhZ2qwpHi5EHBh1DG1YOf88VUeeKypjeQ8wjBvvVns1cdDYmzzx08ddrZLxwsQ95hGHlLL
92VFcJaX8t5u0H5S9uMIw71VanlzYYhru9s6f2s+LWqRTdj6STroaHkrt3IPaeIvw+Znv8ITukpH
QpJLbSnoSx4Z+f641jCrpY2u6BpW2X4HvhvtR6C/uz//JZvD4FYDbsXyY6talbjqKjpYnwSWC8/Z
G7x8lFlMSiPfPzQSw+jAbQRwRpqZlamugmiETkC6DhW0FuA1PK/0V1VSZ3GWdVG1HddtOCFE34tA
i2ECtm97UVbC10Y8oiHQD2KIuJ5kI0qHPKw5CnEJmvaJLIS8BSrlY1arYpjMKUzGFjMMzEjhg5tB
RG//LZPHhVPv6XxBcjD9WCRRoocd0R118cpzWCcyNK5LlklZi0Au6+KjU4MMl35BGlZmr5wWS2j1
Ng9H1p3OF2ysGT5llQd4Dz+9z7Td9vvYrb3vZ+5kqw+OGkKCqB2886DBudgOeiuVz1r1liRCJQvg
pPP80aoSEi3OyP+JdU/zCKWxowF5kg7Ei1vNQzIT5Xjb+k2T0FUavUTKtl6RozlqjdcwLqu3IOQI
6wxc+4zCWCj+lYJmo2tQVPyVvdD7M3vcA70x5zY0P45gmnZxmGSgjFEEgzknrxSQSyP73CqYBMFB
CAY9DstorXRr/0AvYYCOD61dyYjhECySui+TYjEsL594hA2iwENZjawJNHRfnrZeyqDMNrcKFnwo
q2NYCF64KkX+TcD6nXymSB3K7KfI6EX0PHHG9I7TZDuIsBXQe+CZPWYxQSH9oTZZ0M7F7+a17XRY
ZSPnOTRHcAumh2qJeRSD8cd2ITQfS3z+2viRu+JY+J5v30TmTVaXxd/ghLgVELm82MU/Xbj4RMqT
vZ7hXtLn+SGKN7kkGQNm+IusVTHkk+hPlgKOrkSwc3tqC1WDWmr0s6DkNFl1sIFw7nZ1wDmn5zcI
XTbHgRWZIn40GLTMCXZCC2xNYIbm3vaZ2rT8bmR4hnvEzYJdceLuRKryBRa+5rTQ3SMuHUcElk78
Ke++lI/m8gMr0ih4DMkpR2n2sOe/AzoRE+qCwXBVgMAGBEenDIcugS4NHX6i29uuY2eJdauaLglB
uYDMI0vS+9+CiDb2OO6U5DlnXcSsTbJZKjbn1dE7fYUa1tBPe8A/iqI64rOJn1ftWHr2xvQVPC4q
oFY009LDxX1701aY3sTBPFi18T4UKD93iwF1lc1QCEzjxtc1PNq1E59M3slU2zRt6Vs2tQ3CiT6Z
e4ABKBaV36Gc6yl4evistCLctQIiJF3afU1thN614i1PqxCJWOxB6lgpK0qSCW/z40cDKXaq+KHB
pNIWYArYodtbkzY/Vx4wIx4q8eGZFXCcfznXM07YtKkZwjh4Pxdd6VF+IGwFftjeuEtULx5S0Zz8
SqUCm3V70sI7EwYNLhnyLMCPZZDKkKaaO6oNq9jxbvMcaOQ2icwM4Hk0wa+7dQzi4ZY43SVqkZ/e
BobYvyf7JkIJs+Zv66TudYIXkTsWAyYxQz//7MJYMPUrOdqGis0sa5bib5gs2sK/1sEhcuVHkfkK
qb+xdEnJ1Iuw0ODUC/zMIesYV3kA9vj8QIA9iqNNpl1oJZKMheyExDIl/EvHVWvoTMXrrUKeMjUm
6xm+v1ZRRcYq3L2bFrR2M/ZLGzpP0LY2wYZlmb2WOJD7EjefpkM1pgJ87M3RTroulblv8k3Rsn+9
oG9VpMraRh5zkJg8s/e+ljiyqOj5ul1+XGWYSro63Q8Uoj08tL4k7KrKfozm2eoLJ03IECMV+3OZ
eJe+5NEZD7YzNTXKveiHRkbUpRmTKQpr2MG0LJ3CIc+Y65YUtqa3jOwo+jVGLwIPPFyEGklnOFbI
eJc3r/igyfr8RsZXq7wW83NhiwSHN52z4aI8xEkSXMRph214uqSmGU1Be1ru7xHysuZP7+u6Mr3K
ifkbWuOd4OfPeOR43m1i23XyVzNjbj66lZjqzTKdSb+dHMFVpIDTZVP+5I2w60Ui4hSiJB3bXcbx
qTYb7P4f1j2IMeyOmRFuD+3UveX1mPfwcegjpbqmhJTVc3tEzn3ERpvu0SGT/WBSEZ/z4dKnoDm8
sKsld0YhBkSlq7LYUHBh/7u0xOHK2pBmnmi6bLE6SfX8hmex66v2zXBoJSvrf5wboMMRB/rv6eaO
HJzodYjw1EnuC1K41gCFKPog2IGXaafJKOodXAEvQdqeaW1DFVb4Rjy2pxX6eHkkD+0c1f9DC0cS
3Ano+0ZWnKAdglT8hG7id6UETecir+gjM3wIuXznmALnfue8TiwZ97r1pes44DvGaPyjTTjOSIYr
OCYBE/7inn/Ej+eDYFpE2/pRlE2DtXW4eOFaFI/ucVgVcCilowfGCm+d+NRFREiG965ODEwRRLJw
4C5QWrQnD80YkCiaooBuVwkOdlZ6ow4aoon24mWuWapE+ZDfKwrhZPcy38t4JQvZX/AuAUksn//v
a2Bb6YwF/EOaW3f80OVV1mWURwL8lK5kqaA6kM5NrsLxeSgx7ChRrZigNm4iyH0wzsxqg8IgH50u
pfHfTeWp1qp1dZtbaTVv+7NGwLJqxmKhPrYZWWdoYR86ZjgPiGlyRKPG+K3HrLJhOl1AWriLd9N7
bq/p73ei94UsqriRPTFwJfRmdOaVqmhp1bsXcW98OPYwXYf4Gyv8LqEs6XWZ+qdh70iphO4SdJ+A
gehyN6/Alo9ri3+/kWRTK+CT/vkuDQnrSO7aYNK8vxgmhYP5HB65vz3p8yUJQc1f+GmZNmkeZ9ys
xJjSDLHZG6YI8d7BDdY6o+A3pfoFNodK7YTMZyIls8W+N3bNzOQpomlEX2OofsNaknSv5TZJku4m
1bX8GBa9Xe8kMW6rIN1eFdBht8dRrDsv/8W1173obY6IUJhHbWFLEJxqHk28A6C7y7PUz9IeOElJ
iJD2krUjLWwI61liEOq8cfuMNiKLBRqsKUkGauQ4+zfoG3LoC2e4nPKregTzPMWt/Ax+7D83pcwG
5lhtVIqyGJkk6Oexvo1tkdXIaOI5WJycAkvLamZNAULd056x1sC6SCJxBPo9tZThVWfLgOetGdyV
k9wft6YqQr7WaFFO4ykIXzcNbDvQUxM2qITskOVRaudE0IzVNCFVMFjxrOcPtvsOrrbSM7q4nMQx
+JlSCuEffeQkESH7oF5nrj1QTviedODNabzh4N9nioxM1r37baB56VsMn0ZkdHDbU1E+wZyj/apl
Vz/JABEN0n6x+BXEUbb5Ts81gL94x7q5QkjRpI6GFHvOYJitdrjBcdUpVT6C8AMbnvUgB7BQfFBK
HdYfT4gEah61nsqKUgokrlNHygRhbxKewVqAmZsgM2lcD9m/P+w3JeORl+fjkfULqQ0ftMwlgIsV
22ooGuKCWz222UvwkEkUiSlG7UVX2OmvycQ2dJBV92n16h7z2GAIXLozPg56LRY3IQf1hDx96RSF
SKI4oVHi5ehsg7hUdXGJQsgRV7v2ypWecAm9C2tdsfG9aW/jL+1WdbMt2ew0dpKVDy9oRDhNivDc
tiHqEeC6dOwVc2WNeeHHwtVqU0E/nBThL5qtyx5ou4c7uzbVOuzAEpRo4knPsrBc29/H42ljkHmp
uQQEBmN0/8XE71qiLQ7PUIvNEH5K+KWcuN6/DfxInesD217FTVYzAahUivFDXGNgLEqb7g/7+1O2
MGIOZX6DuIkCrOKA44Dop5gNOF6a2uUU3hUlKkNgxRkVT1tDcf0qCsSOaH8kyU07dCrIth92TVGC
FSnBjVQp1NWz99SHGhY5bFBLyBI/AbgKzGR1FpOWT47K72u4xfJDpsa1LSxr7zwERg0Ckjsa/c7D
q6neEVZv4SH0TVKjsQ1QmXKMZ4EADu6GVSu1KR8WNkxSHNc1Q1Nz2gbZAXTJ9m6uR4FFDZOyfLJi
3sjqqetHDIICXBSiyhFEKjirDX0u5WR92HndSIqgEGGe8CXcwQ6PfkvEk6vgi7vGcYW61ubs/dXf
Sb8YiOOa4K/zZ3HCfRhsNtWZalpQ507lxpkErMKJpPHPggvbTXJ1FAPfk/8Zfw+KS1E0GKSOJFDl
8KPeA/r3EB5mKk4UKW07ZA0whZWW5hyxeqS9Ql77QQWhdi+cuEKwuX474alDmzRmdcKrkzKFJuQg
0TbZjeHv+JnoRJlD44ZVG0sgh3K7oSjveSczLG0sy+gDWUnVvAwSB/Qvh6wxWKFCExpOggXErw6g
VidHO4s7r1Cg/haM5FsAg0tjM/Ins+utPm//cbd8gAl5f7AEAQHrxOnuFlLpcNHALSbSgaUe6EZj
51BIwXD+CphldAhEKY3SER8qiVoxN3SDznjJRU5T+lOldKVCJ0EQty6jxQvtScd9d0lsqwJl+Z9n
OQ9xPP+9AxrpfOVCoSvodKAVF6RTBRhbkEwsQ7cHtPBGOH9xbq34t++Ql4mfWnr/StGxMZthZowM
MeuEj+wwk379UWMO4Y/63Mf7Mb4zmR7MToukgXxoVjEgIV1MYQrxzgmofVbBW8MDQ1t2EhEyHOhr
ve2qanxen6qmg+mRKKRlx3d7zmxflpe7+st+7H48hiYZlXe9fj4DMQqbL9eJsHO4Z70E4+1ZMbWe
J4e+sz07cYBbDjewK4gjoi6zQKoe7NBKDgoEZ3YlJotUZc+QN97PyLUzWgDB7WVPkf5dHPfMx2xm
9njYRXu3aDiSxeKNHeUrcv7kN992wkj8oDocKl0yDemIoLYJP308ufan+C3dpgOY0ztL/ccykFVO
+KdTyPkIkfpRixaOu/nDlqJDLg5h7RjStj8Cf1+jtajJXI8rSIe2VZ8HoNLsRvD5u1keFpVbDAYl
VVByum4seSYG897ef+tlm+Sha6Wi8sR1/lJghLSf1RkQpd8u5qI2bOJ252oJH4N9olbSGgIy/dlv
9qEROTR7uTRZxPs6KguVUT3eGGDUbklKFebzSKDz9na0GeJ+ehtYF3BTX53tkPD3fYWW5ToIifG+
4DC8O0hcFMFj9BLOLSHZpaxJxZuEveuT/YU9GXKMEj/F26Q/2WMbLM0ifV3Eyy1uH6cEQtdyVm/6
3dFlV6jc6atbnvQ1gjuN5fJ86bxCVq/H1Qoa//roVNjtIajJ345lvNm5CdhvtJxfbeBkn9/jgP/0
tOXintFAIZz+osJ3jTZGsaHkBC8xOhPiYuhT/tNrS0vJh3OJPuYii14XowoiEB0SzNxDDXOEaOFt
oW63c5UBWlkjc3LkB15aezY8PqA3/BfsNdE6EP8QF4p/krKcND6b6Qn9NzcUeoXRo8BTo1vhfs88
clal7Uu2ZhcTuJJNUnLqjL1WzFFWBJYJxBMo3BLdRJ0kZRgtvh4LgvD4sxjtqjNGLtemPM1RiJKt
LTJdLNQCksSg9F7LXgC1QORrQqCLjpMK2Uh800IFmW00giZ4A8Swf9gNjmYM5BJ/a61PvFiaTivM
hosHi6p+4R/1Q4SyKr87HKGyr4K4+AmG7ixHgznvmbk+SLfSE6/GeAg1KuavGhjmARjUVMQo21rr
ZsymNfpxUtcbVoo1IGgV7SC6y9FuKXOHUBweVM9Bk0fxqVXTvEw/LZrVVI/8IQfERmaELd7h+FPi
4M4hiqyZtlxYfbeh5c3QBNStIKycVEi6jzTx7fEeDzn/otimXVfLGVZzTaZTXIUZxIaQpC6tvpUJ
G/fDAW7NpqDyXpQyoJzJrBOBCKvoHezZmAHcQu4QRJHd+sr5lEux8nRBNwpNWwhA/O5atTZ7+Sjf
7mYYKRh7QfHz1vBUyNE0S5YgHvim6Tt3dsk6OtEm5f+5GpBDHs0rA4kKl8jIcRroEuFFKxPlwH0j
ToqGgwVJpC5YJnaoOzl/INADMCIU1E0nSu/OXFjYjNUhf043ygxgI0/3gs7SwSdxSVZelFfG0Zes
1niJUtQyXa1apKmItMzLDpUrLI8jaQ++sGWT6VaLftUa+sI1yqse6ZN4lyFc8+IagvTrVddHJilG
nGBClZ/piZU9TEGp8a9Pi2yX5BsA1kaboXYvnarK5DMzLSaNRJNLoAZT0Jb4kCAojrrScXnR8ey+
PMuqQ4m5TLKpodOqE45FSIcn52PKtcKGBtLN0Y09vWHlOhMrGVuxVhMpkCJQ4yJlelJT9/qGXUO8
+D1RYjxxtPAxz7g5CAIuwUPSzsFAW4SYanECZbnAyuQoaequnbwV95MjG7qNWCdzRkoOnZNt6v5/
5Ter6IX3gIWCw5HQ4URf5d4/rxQb2tX2oLzOYzHd3JmQ3igKDCsFmwJTx9+BxJ0WN8/PiBowitUU
K3FtN2yPOz/pxVjBwFhWuMdb8VCBGG7sBQ6QQZutcVakwzczf3xjtgruEKeCxBV+DODoyZEmdaz5
+Jj/5hYX3Ohv6h5CuXY1mSOqLG0Jeg7ZPfz/pjaMcq3nVuidywgpE+//H4UO+17Zg3JyFk/h2Kdi
AarsA5VPzClSLLUaljsfnnxmqrImCsU8tNo6l0TTlXjlS1AE8TFcNp5koBF4AqWhOyH1NEJIHGTJ
4AB4RYKMupHn8+e1GbL3+soOQWckxomw6b61tkVlLRZsQHi2pxeidCuKx186Ms5iYWG9gGEoMRS2
wSdeuM7nrmTxF91HRlBqLFkUbjpiKT5RhkTWPP5LPLMd+Gx2ms09kli1bs9rjnfjjlg3+qA68Ytu
pA7YoM7ueaF7zQdUX4GZJbruQLSvjxDCatBAC0gpoy+CzGNEfvpaK7TxM27OT0MA2D05rhaPEMWN
gTtM4/d7fXeCncZQ8rdPhSHsDPjPJ4AyPyz57+NC9PQBlE1amr+GOYn3Y+ll7PZ/AsWvVXLcsIAQ
OclBZYBHRx8slhGo5xvOgbh8MucZ03O27Q0y1lURfywrtvVutoZAYd+IfAwP+V9djqFi2ZmIJsPh
/D83wuSNTgnH2vM77M32gHPrOJeOfbteQduJ+3qjFzpJgXdrFPQxuy80QBGv5YrJQ6f9oX2V514M
sEIyDJm26kS011aKGMUq/ueJjfy++elw0rfxGVJKEsjJMQrc24yQ0VhZNiJzdZRQVjVmRk4x5g65
py8Rv9uV4XMmJF5I9iJUIRBPJDdKRaEcly/7Xf3fDOWH7DTlQNFfDv+ZrWH6W4AGX6xEG2JMGtJY
rehQuJc1k95eO+sd2oYxgei8iNLJ+l2R4IzrHwQVpWK3KjyxMO/kC2xovLf7OTJ1nkAasbNgoi3N
ih5JMeFLNx4CgZtR44YGEoIl+ZxKFAgJFUH4jGuZJfvm+dULWm+wA3aPYzXb2ICftlujiwg59qdI
8S/Qow8yEq86KjTmQwn+/Km4IvCR5wX78eyVzwlkaLxg0fJ+htzb+VxNChdA4YlIoTYeVZvTzQB4
3F0KVnghyRxvnZXbqurR4LO18cARWLeVptb2+MFyYyL0XenX3rru0teAG8QbYkWHwkDoxXs/eMvG
KxSCZBugSjF3ceLLQq+r5ttaFEXO/daVD6D31fXXTge0vl+JNCGqplJkj2nc/cHlMQKC/zpT0DWu
aP8oWqiiKPBlPpT2ihY1igRIuUnscPVdnCjzHS1W0KoAUYvfBzQEa5ckT3sMYxay9lovRCfzESsL
0njgVxi4lt4pjHIPlCFKTBnPYeC1RECtQNJeEG3dWDcq+zicyh6RF5iokTQBKNuRj5VbK+bUZJ65
e2vdOpokI97cZcqBKZxnIv1+/aK4CTsVKnK9M7W/+2r1GTaEQhBwiCv2FrxfDjSpVT+o1rAA5KqI
xMwRiRPfWGTCEXInex0ERea1ZdJZH34LzSIMM7wwQ52LHhB7dlv+h1c2ob1B0VEdHK/0OFI95wd8
tTlG0zIbTqkGVpL/xcGFvCsXrYp4IYslr1PmV9574o8OmQxgARImw+rSvsNnmmHnQY8H1xmb9v/L
6ZRgRTvOV7/YA6BHWBUy+q2DTxriuI5p5NG6zpH2otzn3/Bbag6egUU2207UKJpkU9te9OaY9OkF
yLy5S+QeTgOzf0oJVQF/ITvSLV9D5/hoTOvWVixm+3LJnHYf0slRDv/cHtk1pE9pt9rYRUidd26S
sOolky2Em5ejjTllefH+KOpmvw9WjQ/AYzLFfVVcM9curjzp+t5AGc7DAVLRgLAdcQTBGHkt2rfn
W3+o5zN2D/mmRtumQlV8z/YBKRkwBdlWAPsMLrAcKEMmkW3e8EDU2eF5GuYmckaxas1H3VugoSCX
41kYbiEY/VJ1KLfJKap2NSC0y+mxRaoJrC16elNW+t6PxDrU6pLPg/lk0XGyua+bY+JguUJdM+uh
NoeqL59zjRucqxjmsY1uefcovjlKun7yvDcaFRwfM2nbQLWwlM0IK9GMPg38cumcKy0HuXfaszUg
fRcNS3E10rvjmDkWTe3nfeNCNoBsL2Dx4IC5xyLXWPiW6Lz1vOfRZ7xQw5dPe3JLi+FNgFQXM0mp
lv/IQZMsd2hJ5s1rMi4fHowYV3Qx17Yl0J/0B1Ky58janyH+qunPwPdLZtmSLUFZX/YilmDGj2IN
bQ+0tapecqvhWiqllWXLxJrEbjooGLSqrhq4OLzSEpCLQrbcMxbttHEG5p8wkNxQB1eB/L1duUhm
enG3uFDYP5vjPx4gPBjykpp/wr+aNlBB87mq2hQxKZpcvDRTtaXgu6p1i09G+P1AA36Sh8J9ZRlw
r7OsBY2mfR9jxFC+r9hFFcV+EKJPQL2ONVmbOlQJsK7sVcHdH5iwPo8TLKlyv3PiQ61Czx5xCKHI
MEt/S5+KuyDSXWmzU5VDpjLwnY9OcYOMQCFGAEOchYMPAwd1u/g8L5Lqvd2Xaiz31jcEE4990GpA
lh7WWnpKypB2WHa9dQKmr8yUNF9zFE0f0jc7se2ilu/RrA6tH8hEXgn+PPi90QZ+LtvhuPOJrk9+
De2am7cnaiaHzkmL/Of5pF4YRA0C5ydsuiA9KXTQzkraVJkAWM2X2cun3Fe4slG/4SNEp3uTiJzg
bDTC+/UDfP0buuu1Xu/nNvP8ax6F0mMhkdrzxCNc22EAo1GmkcyCaLTO1eGFC6uiBRe1wBDtFbRU
q6Ske6DddVSOoCR2QWfp0ihZ7b6PMsKnXKalG/v3swP3hLYI3gBcz5wyfaAWcUM8wp2Fx5/gxyvQ
Dom+Fx0ZJjxoHLSZJ9ocPyIs2L4DfCzwGDEC6gi9/tL8xSVkSlHXX/OevN2AGER5DvTCjmhjOdgG
6S4KZPveK/2bCVsLZgsIVNp+u1DL4Aq8U2QsvN6yOoHnRSTSk8RuJDCUm2eFKwELVqiUbjhbQ/JZ
dckCNNygZjXAQAs2QTLm2DwF1a3lO633hyCWvjJA8RbWVocVyQW08AbyIANHkdVzYNAHg7j1qnfI
HaF5N+3sXYk3veSTGrRjsd1eeOjEW+0GRqojDuOvbBMQgq0fQcPVclfphh+ANS5iCMZN8C9nOdwb
ydDnQvQEuEtedU22aIV+heLPlXNJX/M4ykK+PqroYFrcJ7CewpGIPSZrkcCGhbCl4ThIkmfrkoCs
EALWV/9Aa7j2P5TyUGAoiBdeAXlSjpchJzZozCNvEaw8jnuPSFio0+/yL7wOXJPUTPifktDHvN0O
lQVx51N2q82W9EYUtiBrUYplSLEur5JKQ3sqPnFpM83nAKWxYCz27ewUEzcBmvC8TDJBUfN4uLBf
mqxhAKIRN5wobScpWQH9o9yXDATHOBA6s0gZhXhMLUUdQXztrbnZLZpo8Adp3ZG9XkSmftBr6RZC
LbdRmi31IC/Q3FCoYldeJe48DElzIJ5A4wc1te/ROMuPtjlnRkiRPbV1HqMf6f++Vg0Q6l1Z7Gvz
Yu40/oxrSTzn3LTVX+ySfQelvSPgP/J5RhYxMB1M73cHkx1Ox+eqva8cBrhqkUPUPekPmc9Iv0q0
3F930AbswyjJGu3x94kjW1nDZ0oO4fRsv7TqumStIJLIM0y5UC42OVrLhaoM/ETMNz2tzH/V0h5o
bRQQKrPoliYv2c+VZdFgySKPea9Ojt5qHG4fUNaWkY4mEcIGclwbWUHEXqbyMIc5290EChHpwyoj
vwCznHkWod1lvgaLvhO+u6hb4rhwF1G+WqA+nDmBhUqBLvbtIwtHex5ELK3Q3rwJqMZTO/MXXUoj
dJbdTJ/w46gkzrV0tEG13MNFtTMBfn/n1LBP8WMi3NvxVvVHYLmuN6j9H3VX4odPniVNnrMJyGYf
WZIqVuOLZJKZYftOUSg+uJTjdRK+MLXrKDsQM//rs9tKUaEgZ/tGLVykOWUkgtMZNz94C3EjxVov
VURBXh6u/71RB0qS31wEFNzBI3sH/pX8rGGZlia9pb0HrQWmGilD/rxEsIYYrANEM8VQitbf4cmI
h9fi0yAhox7kq6avGFDO9gWNMWm2MjTJeNSsiS3rvSdtVXNvzAZqwyXWebsRSvxsJLsBOUj2tL5I
MutQB0Azee5qmMLDh9sf997xgpH96qVxOXiPQbV+p6kOl+Nsy3zWCmS9hPXYnVf1WCthmkO9bLM5
sUftNmtRKorDkayzGAW2nNzIiLQISZhceVXCninw1fk6c0j/1yMI9plCOr4lPKnk9nNEIxhlG8Ot
ITWRBRPdQbgLLAiYA7MsFZLeLHZzOxMaq8qEe1AmoLXHt8i86IylPKBfEUg7AgdZRuEMzs3UoYts
cwZrqFjqn9bpXZFd6prbxCOOOYP/HYVcHakXMDGDJUorBt0v6OyXjmxImWbTgTW36tbVS5gt/Ggp
h5gCNc82rdIICWIdQnbObLc61Ah1qXGN/gZOjkc/aUDXxD6KlklWKkGW0I+t5CnzxGoJFf1TBLH/
cgxZaEOCOj858GExwCs5K3xaXCar8fsjAzjOp6ZeLecNrJJq6ypajHnkLtZjz+evVLLmE3DDdTl+
y233HYwSF2ruZ79EI9c6Wl5AygBlN3lhL2K5E8ev8dXApQenFQJIDgvNyEJ6JPhpTviuhxYJV6S/
qnP8lTHuHX8VrKuz72ff3fxUIy1xwkVp94Swks63Vsq96WHNsTysCCaynOg+8/bNF+nua78WH8yf
jRe/qF8Li2oRWdTqBNNTIOt+mwydOVcBc9cgNT/wVj84hanrxdvCtULpUblbXSidDqO6KJyiNmge
GXsbkFiEKbqoMAm5txPNU7Caz+TNzqc4X8ueEczgoFTc2pvcTcPOZRmli32Pk245DNdsMkXmhEPs
EkwlQ40ZEbpRl9Yw2322SVbp43xuRIKMlmxRr3hjWI1liXQq/dOawERta7XsjgSzcphIO5qaltJq
apYxVPOvjlNS8w9RNXRAJHgrP4MRqDMpDtPe3VHZ9JBrPSMXvfl5tkY+0cVlFrJ0paeGMaPoGSmC
EYn/oxh17JlYIsLKqpjpJn0Jw9fMLLy/c1M5mhLmjTjJMD3emxS4xwmWs9MsiJ/CS+y/zF8otOC+
gZg/T0S0bF1dPMFsGy3sToimfabBk2tAXF/6t2loAiJBHdboQKReE8galJ8k3GXkpAVAs5E2Bq7r
3dTq9eJFK5L9DjVsZFmIQh/2HJv5NW5loS5iZ/bDsS3ZFbLRhp76fRhMcU6TyZU94ghjDAl/hJBU
reWaHy8Gxy3TgH9z3uXq5Z/Km2yaJZNQfIrv5CSc1/f8v811Dc3nO8PMAFx0o9Aw9pv9CfsRWzT8
7P9KJ6Jv8uUFZM0vAlUu9TV9X+fYcV0M8kzDBd2dLeDb/5IXeZqoJFylTGQY0ZMXKcy4GwRSjZZx
txT7BQmsI0FMIBi3xXJNjS5KH2rArnG/WIGVg/0TZGSG6B3qnf3Z7juNapATGKKFm5LZrazKdeQx
5bzRxvPbShod8DfI7IKXA6pc0tN068uGNWuJ8mjqJEnQBPGF7TyDpvAkVpnA3YOGGTaVuNRZIHsz
KvjVpwqVfOOl+uofTxT5gi1HJhyEic0NGI39+CEA/731jjaCy+eV9CmzFxYfOiCNV1Q5nBhsaEUG
s7CzEuD1ry+BjoKkY+dVEduCEUH9NWFsn6gkkWB3DogRj3cwqJVVCboYIKaJ6rIE6rqPruOLoq6o
97slZNPPUySjGJYvdsiWaBsdsGYtTDhCCDxhq8tOAL9wUSp++uhNSy8g+z/v8g1Cgn3DqcXjlq/c
TsWUPEOIvDQXgQl4EJZKk512/df5OJWq44AehKpPLq0zoeU1PQ2M21M22v6XSuS7UyUoq6RG6dBq
0YJDI1aMinsjvAsw4siuIJ0BplDkH2rXSJdyh3VcJRXkPRSywEs5JxeYcoMMNXo7DCN3fOKF3rE4
uIfMOJLx/4vbIkHvS5yNpVN3TC9JpuhaRfhDKNgEuVlOfPeEzKrnroIyknZS3O1OmlkdamM2sxrt
PnS3CNJ12DAyBIszsrfGlbXosIkLgOWl9gD6E/HE7U4St0rSoqJUb042yPKHu6/K5yMf9bdfQJ+a
Y+4xPKvoqza2ofLn/RE0JwFtULx5j1srQOWLw1TIRWt58e2xRwkrwg9SbQt/N4CigUCcCDznTE2z
0yGoPqcIDQ1Z7xVDGSZ/uU7SJGKmEqonDMLglPlWbYSVACR0OePdgoYct92oFLEB7EdpIBFIHLgk
DgZyZejYvxg66MdQMzMGZ6hXynX5GU+1qkkTEHUF2KYo2BFKdNVNICSNzTxeBf7HRlPGF1183Sam
abdpagoo6otYHDIaD9RbebtiHMw9gzns1qZ7m0TPexKh4UFBduy2iyrsTZXxD2Iaeqzq4KUmsbzV
j8jtQ5ASurrE/nyG8d2NSWgMMvs3D3BZrwhtij7sdzvoKGjGdq331lTkG4uwGhS/a1LFONNNc6OD
POo69SDdkD5hhrv5vWo5mfJG1xow4O+2rS8qOECC+hWqR8NNasg/3BFat0sWFlL8RL1uJ605IFZA
z/UlwDPlXr5ED0aOEBuYRFrAPtRsZSywBEbT3zAKJ1QOqaSWmnWlpu9VScGoiIKHy9cJhxqxr3f1
TuNJi74IyeD0aFkxVgy4dyTrnlx1l6Be2gv9+JyPQkhcBaiI2aUh+SIEmYfWcgQ+9MnHbFlh4dfr
W6XqMZ+tUlOB2ueACos/cBR8mdzsWUQxSIlehKG6+YvlydPCjBBWck4/RWEi5+qRboHD7zNcIDLt
OQw/HjK1G037YLXxS71kBBpAoXn+YhEQo8BxzOKBjLCZKPPobQEmLAxc2nHFLF3HjiW6XUCxG2Vy
+FVf/9iFj8tOtqRaDHBZ4ClF32E5r2qbulaCPHzJyy+z0o22F4iGecSPAAUBJEPhhnhDJ9sCaDUR
7QPzqWucER1XChL7FrVxxbyeWaVru66+9iCIshGQkl50rBUHSbZ8pgsPUmjYW2X7aiho8mrOmQ+9
EwkeUZFqAuzALUJb8Ziv4PFY+Q9yUsyHRN0PLL/N+rZXqFsftbnRcD24z1GBu3xB+XX9GGpsMpxF
UP3087iA+EzlUzkiqdmO6fg7NKQWvZ0nQVf9sW8n8Kz81NaQf1xlIsFVttQ6Oy1PEbPA9lb6kZPR
3GsBQ5cNSLzCru09d04kYrgSo3Yak2yQo8Qzz8OriDOECA+dHiDJver9OUisrHjF/vF2PN2X2Yde
ULxpfwkzKegCC8h5RiyQjq0lFnNZEAzAl9ra+Z52Z1Z7m4DaHIqVXegokOYw3X6l72G0hvL8xNfL
XEjKM/Jgfd6jDTIvsRf/hXREZJqoT8W2GdA3nzt/U10RswL/+EyOcTtZEh6Ap6ji13Qu8VzhiEsZ
jE/C0Q1kITPqYm9xKAaomJgFFP3DkSQ/nToKugsGSc0iMkUpdcca7tPBBdScabUi7/k9EWcEhGmB
uH3lYpStIXNP6akKbfbhk839C9kalm2bRvJvmuy9BuBGLi1IP5vo7/VBdNaOyOX+VcG8lOVBsl5a
9UXZB80GYS8p33Cvgi4vT04HlcbHQBGbOZpdQbxUoW6bwoe/Ow0BLEa2moUtoEInlehryBH7wdQ4
HiCSHVvkC411Ar2L3OEjW2rV7eOoCxAYKWg2Ao/Nt+ZGTa8XNd75nh6aQFZ75uMyclJQAGAkMM6i
63MyvCm3ixNdBBJg+eWdVP+RUmO6v9CTYdct0VeD7R5hDrKHOMXY6CiNdIJq0DCa2zXGvfLi6Pd+
VdY11/jU5v6CBGUR8tbBtp8ZCeeK0JHeutEC/Fv+oX53Hp5OR7mO3D6nGsF8S28RXSmGUFeaZWV/
i9Tlr74WDDmp3WKlmOZU/2rd8pLTJunopZ890YokNUHBnT6z0xkjX8kZfo/OyLCnBWIe/WjL+cqF
5i2E9gazTjBZUplVXoGNB7CufBGZxD0J34Nm0kPSLRwr0cIsEu9LLwbFqWGDRT+p09BnVWm/Nvgl
20VJiWHTTkzo7M4ML8GwttZ2gotlIXQhSNHNqLB7/eYv3ghcittS0phR0hqSRtehuBhB0QsFA59d
Yl71O9whM+1Drq8TZj99K6nLmOlWSskyldCJVhDQG+n/vyKeD7B6130P+WhbC/sPHhpCmKc/sj4b
CBbAUVY/nRXskwca3Hj77HE91912HzamKSoAxyo6rYPdk007AoXcLEmRCezdipN7ZtVZYor/zbrB
U65JKBMcWqEe3kJieD97b0wVTFwIUHFx8VTRTjfOzSKbqfa53qOd5SIhRl5h2hjmbJ0KYeIkwpoP
DZRs7pII6TcRCUwJD8d9azVOGw/+xk2Ft3/5iRWhRkGNSJCVDdRhblASmyl55+AY7Jb8N74xVP6Y
MjBKNoqcmTVdcwo5GeuXQjgpbkcGsiuUQI+B2eHHW1lsXFSNKz08bZuF2LWmBWGRBVyIu+KhATuN
hU/wLx02SIlO0uM5yAPqOIwmKXY3mvL8cdd/goGK7H0REwH9KK+LPMKTnzo6CNcBv+H8uPOgO25u
W0D/E9/AmMx9wI93SOmfnmiJe1SMgrvJ6gp8hXxfw/sWfE9FQDYLNJLFZ6M9jIJQVLPMjspYlB4i
zxsiogdfZA4tS3XzSBDvVc4gBNOBZbm6PJIv7vm8fUTDpeFVDkM+oQzDdu1A+qFWU15X6MCSSJAI
jgY2AsaZTzqxspt/nfswQRi5GKYGfBdAOO2CKBxvHQdB0HCurKK7Sc4gvFXYsna1o/BSZB5TMuV7
pEv1z0V37GkXr3EaR/7dHbqWHqQVTLDyM794Ggx2NlXtJZdCl+UCZEXBe5wYLqeoNgIXzhazxvzk
8nOyBzhiFK4xaluvZ2JzrshoZnRzpUQ8mQiiEdbhmF5WpkEEFmU5LSaUmRYs6z9fJJkWmt6zfRIj
Cd3rYgaucud92PHAbtNULNiKdg0sJPxUWCB5wYwul/4mU9/drjPXEbfg74H5QBd9sL/+dPcGj0A/
ELffH9BxPTgFuc83wYCoXX2PlptmK+i5aLf9jWJTzFoXp5CUOsvRkN9CjGz/doR7syJSHSjZYlGD
/Lb7UV7AwFG3KeFH6Rklwuca3xnQK27mgiKEb7fnc9K+UVXB/vltufVZB2qYYjE8yHFPEGMFz5Ns
0WeIYFRQeuKOryj3l4JNMODNHhkRRUfgsF8wX6ZOmP+hPwhOT1hzYhd3mynymc1+HjWPcwo3oT7U
FzfW0iwZd2iNazwHn/MDLkQdP1MYVmDGYAloY40ETu51tM1BC6x/vlS/K/q2dfr2JbppA/D+/qTQ
MZ/wV+E+liA8jw4Vo0NLy5fs6v3CJ6wJoobFwTX/Q9Dh/PZIuILwT8B//xQQNiAochKDb7HAGdJG
sLS3adWDDBa5IvUAghg3SqjYct/H6PjRhfGNsJcm7NdEOrkL2oUOaz2EOQ3AfWR5oz+iSs84fbBX
tC7DshhuuqxLiXm5PZ+TUbu3zasHCDW0rzqQMVkYFlbRRIZdsfqpDkzVNVVHyXK2lb4JZFjKemKe
0UP0Jp3j01Fb5/EZH4027tnQqrrYVMAFgBqe5CweMsd9RNK86jWT7UZhOijbEEv+j7tZrTvCqfWN
iSoTFfUXlqKWh6QoFMf1ww82vDVHFylu+Rq1KpiOagz5+54IKKyvyLN9hrZtggjkArkWJoAxjann
STCufYb7XhWJtJLAYC3RMW4mXHj5YQU0VV9gAvVAPYKUdl1z+W7M6pTiRjpeR8N9yTMPX03ZFpIW
MKTM7guEPBaMLrVNsv1LHF83Pzfui4WabPv/79wwRUq+LMoi2p6y0ykeAvb4ioa2nZPY0jOHRn0V
LNarLZqA/66InUdVMzzCSywepC55mD+EtfllL9xnvhroi+wKlqkLOK2I53n+LrSrVQjru3qxsVhF
WETajEsyIii+9K8CBIpTocwk5v7B2N6wQhSsjJFK7l2s9nnWhiGcA6edn57Msd7VfJACf769w6yU
w/LwVgYa3FYa8PsJuGlkrsV9/rSuvgwPQ6zXvccpsn2FoPn9OKXveoAtMHf01EiQA+eDbSdKe5Lz
r24zg9/XuoOPwmgvYgJsFlef6UK0EGr/+Mo4OdmpCr7EdNYgD3e5mZpRjXJHCaXtQ96Dn4mXGovM
ugNbBHE1620H3yKAGxsBhC4ozrfbAHKrdWY/p/biiI8ej92zpfWAOxfspI7y81hznCFEp3StQytt
044SrB55U/NXICgWRYv/bYr3dxNQY3pHc/iNCuak9faPcFPP68vlv24losVP7jMlDIQEcRXby91W
zECikIU+DW7QD2AHZHnKrnyNE3O8N63FdyvYnpvae9LdKs+laVRMp+tePJUWf9J0qdPT8Wko/CkO
8VnXAJDBKTfofQXpnMFb555M+K0ufYI3Gm7DLvrOR+M8Y/nykma02NUIlcyIkF/SB3xQxZU1Tc+6
1XhtxhWm8MaSAqAd901QSHtSLVLZWjEUsfE5KfeOwpGUkXbdmzZ38oJrM/6zEcfvpYb7ouQZY+uz
/ilh4x19kCNWdDZjyXy3Na2j36+CeR5HYUBMBE5WcSY5I6SYecSOMrvRUy6FuhGtzSzklHV7REWX
c7V9DlWAgW7cIZoXuSB3DoaNLKsKm9gvHZWMaMvu7eKAR4CuRE4WMQEZryvAGMy1VFCsqIqnCoB+
vt2fmW5SiSLO+zi0rZZHu9haM1IsPGf7izTUnsX0fIBMd6ZtLdBwjosVxQh+66ZEi4ZNPHg3tjcQ
GVzoj/YpR5nnRQzzAZGdEHBGhhMHUVQ/864dRqzwtp3MP9XqaXEcIIdQ7+eurq4ZMiKwYmgPpGYq
ndxXpEPPB0xk5v/r4aFfQe67Epdm8PjODjuXVOyB9r7aFY0XkE1XTt9JwOONu33dKSTSOLqRkDGH
dCTRG5ErFoAVOW77bvGmiDzIfmBq5n3blSD2syp59WUEy/Aox6V3FS2uaq6LLqrrLp5nixz23wky
O9s5HpTszRr76Kuu9meX3hb2RgM1uEBNQSa+LmnITrPNsdGYGJSU0+t5EtA7EwbzkKyOpDIXvbqh
dlHGaDZ0k1B0syX38PnaG56y3H/0vP+hB8iOR/JIWpQfilbMZVLEUzDpr8hW7q7NeQtqsRc0dRFx
ENiMjepJn/5+xti4pcy7pX1fJ3hsqBX0orxuY6taSQDK3PvUkTnbTkXsnSYvSye9iUd459PGjfAO
tVKJEWISDaRunl5lKC0HhYBPoS1UF84mlKA4wO/UK5O+dQXiwDcRpnTNTe9pKfoedNsCoT8Yxnfa
co2vcAwjtRWeYTq5+WsH3BYwIy3y4URoyqYHd1xoY+x/louOHMhyWrYqvfwpADD54skMk3dHKKYL
Hfd75HrfSq/1XlAogKPIDExFVba0c+pF/eg+tajlBZF3WR/HrIrrEyqYQQdJJX3JKbZYCB+Y4pBx
kY23iDc+18ElvXA/egA0jonYpevH0M4rcz+MoYv0LEsWDwmV203809yqLDa8m+2PWqUxOg/3U4Cd
qO/xO5fuJ81hdH6BXRhQLTt3g0m0COXNwWJXT9zHRjQLKsULZ0f6SF2o19CYFZVLGCMDymwFpWfO
YrPM6sIYzRyYV3os2eL49wusS2zt6kx35+QrHgcDKuQDw9N6sZY0lpBTl43pcBAyIjcUGafQ99bT
KTMwxw/2OrotAHfLA8qehHVmCruxAwU/krmM1/rN7YEAOUkp/5H4SREp6OxSZIy/ksna5pZZq62i
9xtcGloVvC/wPGCZUoFNj89n5o+APThl4fCs4EyeKC+4xEibZjRTSG/54GmfbaY4XsCxIAgqZi1r
kjRVt9Nld3sEnHNc4KuYgU/H52WG99uhXPOCXgkOOFnBOWG9tSXt5Aqfaw+y6E3/fWYUH81ZFcw5
h2etJH8Bi6S8Y/C6aMFGXtnBWxc98F88zz+zCl70n9yYg9eyGa7HXreza55hiwU22x3ixvieT7lr
jjSYZWKNBDz9lJDz5hYTgQju/5r12KW0LtO9dz0ClCelj3LSvN8i71ekMGy3HRRi/o2yqLprUyoa
A6Z7G2fSu4JC79PTxC+zjc6rDqeomwCzJi7CkDLcyxxv+Gi9mfkAdcxGunyHNtvboK02PPmHEpc8
UcTBBx40P3YUPxLztLoOleEBzV6gDx5UyP7OViRzV3XYVbKXMoPYfAtw1khca9bxJhhmYVQF3Nfm
qzdkOJjR+80vot7CgpoE8gFIHyIDebM9ftmy3Zbg9o9mUxQqs97hvw5rdK7WDBsw3m3p2IkNs9C8
0rO64mc61wEuRcv1k8aQYpplk+8kt+7v02UOP3zkIiSBuyEHtxMe6+NdD6UNjyxWOH0ZvuPmMEfe
8AFSdbCplutKgWdFwYmj9khNbiRhcIjzObZtAnnW/dzBz1UlmdWlXIhakE3y4E1dZYaMNIP0ePf3
w8x+WEmmBXWl833AEkavDBKqMfOb7TY1tIkCNt3BzE3B7UBvC0/GItht+9rgNpqpUCd9ip6XB/+L
ccH8ZK3/yEa3qYtq1QjvqyhuLwXKUhOfjZ2NNvUZGWFyv6vmsM1LwWCyulz9x+kBF7h0Z6I+tYti
wKGOHSbqvGhpnmLYYy6TUrKMNSxvs3dO4VJiQPS4bxtmAyye7GFaUM+WylbnNczOf7LGyutGz4uc
WlQlvF6Wv43NipNCktLxFx0vHWwtGYpM0Q4DcKIaonDyj7T2Jdhp+sQXn/DJR1MtcFpshAk9QRwL
E/j0xdDl2Ewg0ozKdAFvbQyTmEVLoDS1zmEMJGjLAGhtGHcb/DSJTcPWP4twlkd7bYgvWlT50qFE
vdpIOz+NQxf+9PWPph8ZAnWRGvnvcA9ZlkZJvxZLGuZeN5xdirIUETZ22ocC4P6TqUkdMYwkqtmv
gvxMtIHN8+EKbLD3CTLttkvuue5VoWnoHroyhEEGedy+fBqYq02ucpK1vv0mFC/PSrOSZEN2tdpy
myexc6MZ8N6Ra11/xeb5wb2jhPO9Gnr+hv20kd69PPCq9apRDGO+W8h2/R3pBoE192jSwGPRvh6H
/hIgSx0cmiQ6SPknHm9K8FMJpYOaJChaMZY/09dOlCUltIplcB4dWyome/fr9q9rimkQuC17xc1k
AnvvbRE0JdVKtff0c7Ocr5OdGxztojDMyne0qiW3evtsyRwP+Jn81JW++Eb5TGqCetFRLVA3vLhQ
8GCrAPB41+KxNNWqAIlu8HHy4yhIqQ7WNGg3rpZcPt69Ca0z4HXc0TfxdpUKzMjnrcd3XVmbO/80
xPWJdDhCc2arPEsJz6OMT8j70S6jlO9r9enFToLI98xHGUylBNpFGiDhNsIK5ogXlUUI6DQsoVuC
LaRkNloxMG1DutI72F7wk6ntdgeWGlnRvMlWW7oAc6AzV/bHUrYeEgg07f0zUFHRqE3HWbwMVltp
rPVRIL7KSRRgg2Lz2tsUUf2w8Y/jU9+JaZVVVID2B8O1lRiSbllrgKlKaYW9PZTyb8FtgiMP7Q5K
th/Y2HroeaQw4QyQ3JZn3HxjUIv5VcVPXqGF/sWdzbXccyEM5Q9QmU59maKtQl3gI8H0nhwOUfZB
Olbtk+mDfHerCjbtcs4AILcNry0hmeQ8abeSIQpTffRLzm8HKW48ZvIHBaMHsuj9+SiyBILkiusw
B7DQDP67Kuyfs+X8D1RSk3TVikLnLJFX8sF2ra/ib2aZQ90JrmGPu7DGusutQ0M70iCJMrNzsfMl
DNF+bO5YTyaZqioJrtQOc6f/yFnrFGWwsF08XJ43HErtxW2UkCc+f+WVPYohocnFtVvyYri4R0Pp
lRdxXa43LBjw1iT6UDi8vQ4Zwmb5V2JYdwJMLA+wbVsxdJSEAuaMW/+zRhJ+rlKbzM2bhNiI4Vpc
IzC0eWSfMHVSItD//VFy/gXaq2BUPexlIVWXrS2sBFd1gKvpv+yU7z4u6m+yhu8tOUFbceebunsO
/rRuZdcIkiYZelBSE+up0nHUAu62UaCPpIt3kdf9t7uP0hX6KvZf483RXVwC4OqgtTEm5QpP0fhy
TtKu/s1vcUCI/Z3SGzL0ndZlFTS8oGLpcUq835h2Jgyq/5rB2JpQxowcNrgQDzcRLJOf6ja2j25Y
AOql/wiLUHTUg0SQUGkg4W7Uh1TT6k8roqR8mVj78sul3HW/sieDtPfTYrg5PpS7/rJYTb9viTgE
WyCNreozZE1Bop6SyXEJzZ7iidcLNeROuGct6qmFEIrUTbVx45q2CPoasFnHZcLINnBcyuPakjU+
BL4LIXlx/bBMIRk14zTIwHxs2mSuIxFly9rGF3FHMG0oxEH+LLdVWaF4zu87Pxoa22ugs8jFfs8w
sMPwwiZrQOxlFNH+qcnZd7QJLfh52bHRhNgvZyYY0u/kiYk5wnsbttwRlRtjDz9bMxcRak2akei8
EVFvYbnx51ryp3Np1EQW9M7HkTO7lya/yOB0qAMlrX+JeM0qLEXz+wUrOIDbN9f/t/MJgypgK2J9
OkWGrPy/OXX2HjHumQqDkp0wDPeMx1GZyEayx8I2+jQ+PfPmbt0WiwKxeZiTFJolyK5Hac/WLsDp
wt1+eGjC6dR3+T7J3BG/f1mZIYLYahHmYEGvCWzYXMAdl03cQ/ANVgJKJDW5LP72Gon5sNIE3WtL
0M3ksHPOin3ufPqaD7Z2pAPJai4IoPUgraaCVXPKzNS+b49KouAWx9UGye5JTs0yhN+lGzuOPeVy
uwM4YClDw2opvwV9Pt7s00P4ppxy7WI+dP4IpvjihFZ1CZjXER7b6dYJ6gxuMkAhDpRbyLz27ET6
DoKkwNtxbRmVsMCAXPIgdYYX9AnEAgrtGKYJaj29aSg1GwsKOw5+jrRpodT9bCceadxUDHLf+0/S
44/HkqqE4X5rOOd2Fc4+5EmtRBDAVO/qUH3Ca12q08+hguXE4jF7wHiRQ5drMXPvumx8G4QDp8OR
NbqtElXizNlpilcUH4DHsX6V6X39PzdEpGxx4tOYY0P6u+pjpF9YcN801ubk02jePihsfZFjjz+n
otYmqgpoQ0SOSTQmeOYA7qM0NLwCwRDOnYf1UMDDXn8i+FCIZtwYgyMI6kvdK3byhwmGmaSHWML6
/Tc8zizJqgt5J2/PWLDrpJeEMqgK9xDeAz3Sh9MDejhm76Zb2hAs4uX4OQgHtFMHhE5gCSkk5CZA
0AR42OEDBvtmcv11cK1vNW8YN8GN4k6s0sveGITLBXC1b8hw4WCtXwb2TT0fH4/HVJJHIY4/tgvF
hX2Gt6FB4nhum8GL9Y8k+lmS/G0q4w1ueAw2DSHIeuE/7eaGfpZR3cMR5zA2cK5QtWRz9TF/9Tnl
58PqF9hPdIRDJqHJDZ7h6AD28VEWf46iECYb/lNlPtofhCr52F3bNb6JALl9PVDKCN9lsCu1zpYQ
g3xns+yTW2w1BpTYX4eI0I/lOWMmDVxxcWswc3oUncO1JPVL59eS7X63UYOh2zRAIz8WsliOx2MD
zDA3FTc+f+LVVv8EWP9i+jNlhph8L47YGKzL0xLRaNbly8i4mbPgvRIrfA+94jniQlBwrAChThod
zEnoBx8FoFps3XgsOn3CXViZFw+jqCeD0fOO9UGcGzNh9AMGgpfLG1oAFiPmAJ31ZI+iO5a0xQDP
aMQEituurLSABoWWhmf1pvCwTax3/JvcOWmgNHjnlKg+UWFmU6Webs4GNYZsl8cxFq+xW/x+7H1M
tAl8zqDLxfZrwKhM+RQqMjtUq1I7BQYNLxXUGHTfOOw8AolxU3gOcNjBZp0yvDRHQpDVTDJxa8GW
UaYFqTnk2fAUjj/lY4kIoW4trjvwYlKQIFdk1DdOv62S0vAL+DR8ADNR46sMXTM93MP3iFnI2lfX
Cc5QeCwSGPlKEJuwPhz+94o0+u5KKFLctHwR4tnJaiaCR668iO6u0+Ty/Anq5rc1CDYMEJE6fzes
4hxagk0BQGrpsNofOa/DBNk2c6rTsxAQ/mGpH7ZEts7TQ16ujfcvsnyK1gUI2IEtgsxgJn6SkbNv
p1MTRYuP1Z13aWDmwTHsywKL2NXb4Et6OFx3i1zWZxbTivSYmPzyCpd4Ns+shkBGR8Ig6kLNRYE9
Mj+nRxcg/BlgXPXd/zrwSTr8LeM9CvyAJdahrnxfDb0KV/JhNje8J8Dr1JU7n0DPwXgvubQf/ers
FmiyTudcgJ71L0WtmvVsftINtvU6XBoB8iQp1vwhiLj7vRgAQIsg2RZCedZidF2e1AXg2RcLOVHj
3NKaY6r+G3nHckkcDWfYIR/P8J1Bu4wIWI3zWJMposq/KlcfQ0HGMH77auxlEyWTv7nWdMGgGDYU
2oRmRl8jvRDroKY/AbSrkYbBqf6R6MWFdY4WSazEuocCXb2xf0NY62sEG/WS6cxY0DVwX4SzLSQb
pVT6ArIJrcw3lEmb0OKME+oxLZ7osw0IVgu21BTU9Q0X6puvq6qrLdEUMRSa/oFvP080/zy1c767
mF0YTmvHOVyjywf9PVCLrvda090fL5EUe/8iCuRY0bDWPXOt15d4w0hz+eUuZfJyBnHaIDBbBkMy
p2JRIHSLvW4J5oqYgeOCl+uN3UiQ3Z/S70oTS3wNSvNq6+Bo3JtekbcDzTxGOoL7J1PvP4eHC7Im
yNy4O9XjgN4ykK81SMyPS8r8bxt8VtEC3cTyMr4RxdM68Fwvwq37vaPDwlFrz3O+igaUXETtPzY3
7ERSrLaK0U4dKa2HjmmlTv7595rim6lqKVgkkFjp3/HdX1OBIZF4+qZdaoyuswulKTnZ0MfnKgtI
oAt3ggECXOFXdm8hgJTcc9NPKB6ZuycdsJsMEUduCXyDRlH9J7HO3xStBlIrYKSAXSVQRqd1ePJb
Ry0pkMjhCTNoHiCgQEhlZu8cep8dExCdGnlQeV7w/JTWawlaGzRSwMQlujS3JPK36DmLoBjJs6hp
ETHSUIPQadX1nJrtsQDHv6G4a56joF7g9Wvk/R2ylNdtt0TghG+9+qixutV9b/xZy5+1Az5bY9lq
QBuoKwboDhTYZD98mAYJ8014GfXEcxGG9xti40aDtN5+RBpuNHh8X8NIOpRWeNGSM8Hi/s85AYsa
pfRq3yJbT2OG2DQg3j/EDx6nJjRM6g3fxG5Li4wdb87tjiiN3V8gWRir2ijQyeEaLaMs1yaVDjbO
gU4liKrO9JCzLzfzvrnEp7JZbD6BK6n+473FN0B4B/GkkENB39Riia27XO7UdoWIWEAlUE6ONCSl
wxGX+tBgKDjQmB0o6NmeJ6DF0m/TcbBcz50loV8P7U57TNfb7dotScbBkVx54b6uoGlyjLvj70g7
BHy7Et2l5+tHYo6DJcEWPn+GrFEfU1wuk/HQiAkXK+LatJqc8139repu4sbIzxqgIjVZF9/edJpU
yzpe4+FUslq/hbLhdjFmz5Fx9CUo/lZtfm5JPOoInOKvWDdoVdSVWgRohT3k4QWNDBucgcRG7/M1
zwdd2Kr3qrcUjIRE4tXmWjI7eTb2+xp9FWvMLjOxMp0gi/Nh3QhnvYllyEt0WtMkFd/7oCZMITcF
aQ5ONoefX1Ihg/bCWXlWHiVmLmfbdQYAS5BK4i2gsj1W7bNskyCdeipfbXeM/7/fII3mt76E/rhh
IxAv+/K+PFsizBkp2Onht9o82efNk/LgbnH5aR9Rwht3qRatUd92rRnjRj3buoyg6dYf/BpQ73At
juJ+RESkxcW5iVdHEU1PocgJl1i/CocTZKhopivGmoOiGFfF8cmQVuu571rB6hTxnhHoMq5Zjoie
vm2i2CIbVXgAOi3wFrsjdHB7cZiI/4z1gMTo77aLEyGDkElAYBMseFEoSXDLR55pigIATiMIwRaa
RKwSTMbUIhdp3ES5W7Md2N5dtWGZ7jCewaMzpIiMiVOQNQ7ns7Pm1+PukuhC7xuisdIo5A15qukI
uD/YghRJM8QBqdIR6qDcKpTjXKoDAeBKaWO0QHOeSewFOzj1bNfxnxKsLFgtnuUl41zq5mYI+WK2
yYeOUHwFthLSSp6nKtu1fH3h3S0bvkLZQcpx8wYcIDguJ0F+505wwIniQ35L4fQy5vAZdg03WySH
oo/bpDP64lrTKjLmaOo372zXSEKnwIMmG0t9kHsQ6wI6QuaMFhgYf1gOJABj3uiDm923mmNhL4eY
xKTse5UKkT/utDD3nCdgT5+80gFwiWAKyQR+b6QJttTjtupFXGMnk0j7NbRD/uhwIsHOvj7m2lNj
t2tktCLsdNfeNKlgyhtRZwSSdK0Bj9GNLlzrsgQqLFJloYGIKzzPrM1UtbLxELCB+jHM7YAagn2I
O3Vd9kGRztiPBn129Lj1dmqqzyOQDbK3Jv8aU3f9bwBruNTAMqYOlbrhLVBorc2WUFwpOdUjFEzd
LcPvWWFgVtIEulpwLNLTN5fVMzqOmXsjmRplYogLMga7UJXZM5FIfYiRCMtxOrIiroauXfDWwF4r
mDLgamsFBuJD99Cua3G1oRj6iyLqHRi7HYdYw/5kvP/6rCifrEmKQEKVNvD8f2WzXPnMXul/Ur/J
MbxWVbJVcNSsBnayzblADHsyDCG8tQN0m/5Bt+oCDMbg//QCuhPwEahUzVxjnVxuXBBinoUy530Z
ZYCHxOp5xrNWGyDK5aW0nN0A58KONP1SYnbxJ/P281cQb7cm11WuokZSiPx/96fFmaQEeDSuvL//
WtudVn8sXHwLRGpqDVOKh90VX7VelIvhm2sW3L+/bVa3Ayo/7sjNfRTPRQPtjKI8NyNMkCwIqNAe
mmT4880bX2PugJOoDB0Vgr6lQFqj9PR7jK/blO2nqGQECxvHkGF7l7mqrz6u4YO9KE4f0Fa6jsWE
Pmzhde2X/QMZcj7ErpASI4STsT6FVmUx//8KDg45QS29NjChe0wamEnDHY9y4uu0zlonT+0xnK7X
qOowLvSp55nvXy6CHLEYRaICa0mwpNB6+MrAGxydJqtmni8x6ZnysDVN2tUvNN+3AlpkVfyWj7/R
uWgFXbU9fZ9aM4wTyp09pn6EJ2Gda+N1cBaIYnmJIscAfGkvky3QjqZUvLqmFviwoVgG58A07YAX
c51Not4e7DJ8MiWROHyD5a6BC12L8yAq1ip+1p6KNNvYoeZ+q1I7IyVrDjz4uIGR3nqKAvdNJI/X
CaXy+u5oZQo6MBzhhafjUNFsM1l3HV9MlvVzzxWPsNJfJP5czEg5qWkwvu1/s7o+YX1eKcYQjjFv
WJcoTx4N26c8v3NPSmXNUlX148rg4VOZ6sjros0JsVp8Y21OMBJ/I22THPzJg4efA4nWbPSYP6IS
I+L6kMYqf6bPww+B/7u70j5w7rCuVc4hAq28uaOoQ+gQNNFO7HMHCNp9s9aK0kfnmvZi11en1ke2
zEbtp6AS/22yMxdvbcT7A2KX1QyqOMv5XhonlLvQeU+ID1w5AFWH4Xv+/Id+AehGXF3BKckJmSrB
E+YeZMsfkcXXO61xXgEFsi+e4AGzhj5zROFMJdsbcRFPRAMAl3tqG6t9zy/grsbv8bAKfOcfO4PN
9tungH1m/m771j/NkOCr0VtAQRhxfYMNlEoIiwZPb3L4mzBwisny+pGvbAY26Ey6r2XmslXpaw2F
iUCqNtwb1VuFFjLeIvaVsaq/gT3gODe0pMwY2KSfatmHU2MRhTiS0hpc0Mo5LczEPIzA7f/I/AF4
sM0YS6MngNBnoGENqNktQ6IPzzBNdLUv0uAokxu60pqxWH1HYMiY8dPWGhKllKXPpKmXWknRm8Hi
Ccud4cO+R7e6dF4XVCHfjP+04JtgZzzlcxEPAyw+pjrkYmBuCAq/ISHv+RG2JCPwY/0vAPcMQulm
4/1A0uRmfPhLiVUjiyv9ZZcFRZqz8wQ9Q4VNFVaGCiCKaeeV0pcbiUFV2o2N7KMjiZnQpSYMiOXq
yaeqNOAPGoalUIjlYBJljVLiXLUo4TeBp4hCagYemY9Fuop+mVUfoe1RhmRxqF/MFCjHEgSiM5jS
by3M1Vfe2mhICSiQTjG1dczYOUdEuR8HVilGsdTms1vTJJGx9Z1d6Qy8PziZEIrgRGtLfMvXbQmg
t2/w5Gg4h+TjOpGZoKq810QH/pZzVokVjEDun+wNhGlISr6Jx4REoxsVdc3iiaJSzjYZDUk38EKT
jDFF0IhL2UqOk/Tr55L/JEBIBfFyI8fLqriVVmoo5+Ny0vJwpg3db6FnjwRlnW9fV47dTB8Z1IEL
abrXXhodZyBT133CPxQxBScl/PRvFk8c2TBpwjLDd8pV29hGRKNLcQliwViRjkivAei9vBc3edIQ
vLFc/jZuZs/95+pWIjkmZEiGkF2D4wKUdpBjgcRaPoklZCbw8xdd0jadq3CTcGjJrzR3OQHQ5b8F
usJYv8Tk5dXI+aLg9TDdL5QA+rAYlcrCce7rOxgRLueju5oeGBQbaDoOUWGAuNnf/wFbyuV6EHgc
mGd6DIcKe6DM8mapluWSCtz8e0xklG2BDmLG2ydD7yC17zRwveYXSKE3lSUuPlKpvDiWWNVoQsfx
qALaAFV8l6wg6wpO8vVDj7S+BhbfNp4Cqp5Wh1GuflUIYJqR7zj+c9j/CqNa9Mde+kWeG5eX6CNz
x0wB1erDN4vv7RyLDAPcVsXjUJAUlsaXYlABxjnPeUMqlr60xj30r7D3zunspj9s+xh/nA62gtT1
8VJ0OubKv/dt2xl+xi95RRDZX2uzlsVnvNeY2L/wO9PgySqQ0zfDxJVc+gXiHRWT3O57FMlE+UQM
y+sSkaJIQUsEuZm//yqi0zhjGQXgpONmoVwdZo0Ugj89ASbdp6sWNwizypM3Q/LWERwpS8V8nqFf
0AaW9EQkJQ+gjSqVPeyHBXHT4w5Eyv4k0MxeM+SnSb75QLPKosJoSlFUTuOAMZpwL3mOitKf9c5a
P4uwFcC/DRZpDhkOOSDCUA0U4pJU7mzI9sN03f3i3Y3jO/BKu0PbLRzKnEOuZ39HLlDuWSno7fFn
SUjisBVW70DuBN/6tuCdJ+SHZCXH1Q3E04FZknncDki84cOufF83F86xq9wsInc7u0aioZRdOdCQ
CNvDe1wRcdmE9qRpOtBrtK92vpxqW9WeeAmQw5Hq93nb91wZjjehpxxDYG+/u109Bwia7DjKCBN8
FqKEe4qpvNRdv8LrwlRMRjms7nlv7pFyLA4zMUIdOpglkGMRHowrqFIkyPQXCr3eerRxOPM8sLeI
aSzO5S7J05JIiXkM4OR2122z7EI5pSGbml5xl+lmIxCTEQWdvAndKSKx3Ty5mfL97NFY56OsTvnl
6kLctvPEoScnQk7joDIiplflNLQbGvHofY4vbUr+yuNqmS2Tk7OC3DMdBcI0yV7exdG8C65rY4nw
t3jmOLa1g+tk0nNFUeXnHAJeb2k7bWWGRyHqGV00vjk5oFEbXETff54HdU5ewwjWXAhqR1J06CXB
M9Hn5UZxFWBU7pAMhq/wFTyWybJI9pkzlbPOnivIx+sZ3KXOhaxuf131UWi6Bfl+TY37otch6zCF
YLChvYFQavvewDpbZit6fI4HbQuXLr3CJimedaxuf8CIQ2/ULG0F+KPIWcv7g22flXKhRChBCCTT
fw9xd3Dvka7rEjJmpYooxXKMAlgrh6aemwsVYnw75XyIWK3VNfDA5ZSbB4qgXkpLu0fqnAK8MrAH
tTD2qxr/LeFTKp4uyGjLSJUDufId0cFW5jl7cpWfV5n89y6KKIpW75FnAfj3Kt7I3o3MnPUgD4S8
Mo/glUSCzL84mh3tkM0cRbXmwn7XrFJZ7IBXahEPh6ABlBoJRPS8/3K2HGlWd0J/aPR/jUjPF3B/
n/gAPI7Bpk2y5n1esAo7FDtslHU1dOr68MyzWIOQNTW9aypE7iGIZQeoSGDKCulg+4Wmn+Wmx4A8
nLh16u+/nQX72IeTXcIUojeebJeFzXZgIdsKYUAAh/xDcRyOnJyDM61e77AMMV1D+Jun1Y/G08q0
STvPjrgQvsUxfoXNdALgwfpza3alsR634XgMHKKtA4eyoHXJMb6oY2RdIs/0Fe0iy295laATBBsm
VnY2/RMdSDl97SrcwSN2yENqFkOme8f7ywCDg7xDWtlFlz79z/fkpA7O8yaFyWZ/wWadxxxQ2645
OgR+abg45u6rRtiUwouG+B5K3giTKvHY/O+WO/T3PIz6sAX3BBLsdRPfRfe07xbvQKC7X8pfSmn0
7LeNi5PJkmlFmxA//AKzlp/47kAtL6OUzkiCryeML3N9Pp/bF/N/694R2zzWpzDWvilcz5ysawIW
AApd5pl698hXYgiQ6sIxB3lmniSSVBxdJ7SL3AXOtpzNQT+w8UWiQf8YtVthiwjfa/GEKgWgbm9Y
ENdlXAC/iTWbfM1x5ez2bCYubnoQV9nSj08InIzPms3yS7zsJyUg64G4NowOXypUrxR9/n7jAw4V
H7ipeKUG+a/hIlPm6o4TwQWgT/sfdA8huRWWtEAPbX2Wo/4VvQR4/SQTht6mDs4NHGSkmibe3v//
jiNivn2Pig03TqWRFjCqlIfxmQPyjOfVN7tAjrixJ1MyP+Gdt/061b0hqc/0jkOA5zK1zlfciUaK
bvKJvRVh6YHxEHak30N7MtU2rImnZxyCW0LYjYYF02uIX6qfCX8Dqca7smXKYol0GEPX5nTAiYS9
rdRPTbG2pSnfqF/hvw2ZlBy7BsOdi6uvUFGQeisbFQGBfdAZzsVrl6OARciq4S/ddkQt2F17cLTI
KjJkL3tFqmxcBvdDdlWh1ZnkJUGMuFjQ9X2mwZSPhXB3WMKPPb6MSYb4WNFm6syOS27idByFToUU
IrDyIPQAELfdrxly4HUjslxrXGnAT3F8EDa7jzrv0foGfbWUTzBNv0Vpr5zLuZcbFfIMrhlOqHbo
4SecrbEAHl25YGB6dGMMPkDPtlf9hd+LKU0dNTNYQcs9zdh/wxHfljHKZlzSCk7qVj62yTS1ULcW
l8FGYrh6zAteKl0Xpv1W4wMgKIwQQ+BkgVQbM4cGwmsFFWTOZs7qouwRmB445izM6lDwdi//CsLS
oqvuRwLz7zQT6hUfhJIIcMsDsnlzxFoVCu2ulrUxR49GwS+wkVB12ax3zKnRnOF0JsCa6DEubzuH
7KyHm5SwDrG9AAueVmIvuXNexbyyoT6Cyji0uechltV4rlB08eQYxGQmm2zgj6/I1Rcht7MkJC/1
W1O8EIjspQ3lNYpC3S+lcV7GCFCoJRdPdL5U9OKFU6EMTpYarZfI2eaPEVG/47lF/ZVnysc9R+zN
v/Ipxi1d3Bb+ZtstHGDEuYh74kme5dGuMQiRA65pK03wn/r5d97YlRa/aFVKag+DbjkQC3IrOfql
jGz4bZkdNV4wb06AZwjxSxcxrHcSR43dS+iuVMn/rGxl1yoiqgq6ABHBB0S2kU8jL5qOCSQqBIdE
/mj0XIdo/IPkDjmTqf0CgCbfW2Cd05oCx1Gnxq0ba2TZfefP7LroNH45WlhMbxofazwtAD0umdt2
TWSxXMWCT6H2T3p4gLmsSvSVis8UJq+ZGwhczUEC75gqElbEcc+/FrKHFFItwds9KUgxWXShUutK
5GjWN8iUb21CEsb40Y89khIi86DfyzTnGbnBehpzSoOqmhxoJ8Knnrh7FHO5NCFbwnVrZuXpjiO2
oGbcrpIf5FJllN4ahfOIA5WuDwTDeKla/ZJb3v47vGf25fZRd0srv0K6N2AwO8y/EwXcjp2/Q3DT
O8lNGoxxysLCoo0+L2eidUZfC362+1giScqsi17BM4CQaZJda+0/gxG5ydkVFshP/gMAsS7MHQgp
OeI/8b8ZD1ej1C41/sQw5BgsD/tNBt+8Q2DDtJtjVPd+F3JtmM+rX2Pqd9ll/Xsb9NDD/BWLhmRV
OOhKaWR79Dp2gqLgz6ChGQTxZGy4gVQl9VLsbKrc3Vs4u7JGbILaVyaNV0u7M0jQwB6fcP30YgcX
du9kkurDLWj7zfH4VdCY28BR4zqminUZXHcPq95F4qOZunP/1WHmBeKF9T07h6lZ+mdj3+qw584G
ZzqTqf5DdMkxsMclmyTZZtYB2xE//B6BgPR2niYBlVoHAbwmFsr3vc8z4wddjzhyOzXPYY9uLJ87
D6z7agiVO1tsLTydHcFnRdZO9oFH+PgXL+QtPk7IebZ01+nh2knvy55M+AgKuOr7fjPUVkW485fW
qbsXR5mq/t2WZDw4e3Xzin32/tRG3kPVqidRUmpgHfBOXkxLDh9Tw/9rHsdDJ9GzKAPfwaX5xnDK
Y1ncJ4YIjTIEI1HfhOhAjjlhDLndg8jQL8kxExRsF1T2t/p9Kx2rXPfekkWO+ILGIJ5WkRygQnTr
u43myTcXxcc34Wpdw/8Zrg5sRapUCVayqYPc1AhWB23H2hTqgHVBJuDTDJZSF7T0D9uF40BDQo2s
mZlIG9HspEXfpNreUsELu9UfyKVjj4QvocF2DthrI0bK2wxBLTVHGoJzh0dk3tDuyA6SMLVObB2M
AvmiHjDGh3d2akZjEg30VCBz+43IiT2pggk1GeK/k69UUXsYb/M+TX9gnzEUxkPq46mU+VNJvVKH
t3sLGurk1LXoGKdr0DXejmhVHtbw7pOHECIq8ZoCC3dtk61LwnZ7gc56j39pHrEti06LnKNMqD7j
jfECi2R9STaMXZNWellzsqueZu4ompQM6JUynpNwaLc+QEcKLpOPZ5+WaMh1rcX8VBU++bKzLYbF
vH+hQL2xS4QHMLtQ8OTsi6Oyi7BRd2avDwgHe8jeW/k1oqZydUHRkllJtSyAF4azWaJXH8hwKWF2
QykV/nYUTYObLXacbRj9anBL5UDnkjjPDmqnQ7ip4QesXEKohhvKNH8Xav+CA1PSBnEcCru+OTSq
/WTgAdLv4CT4UTtbPotJwAyDMhRvLEfcJ+AL977bwOckmgZM/EWa291xBSkwNnKwLrm63EotPq97
DVXX0MKw7Nb3aYl9+CzY124eD/EErRyaAeccEz+7joKH6iJUEy4te51Mpu+W53JwxXSqPvtErOTO
ulCaR/YV/eoN1JBLcjmCcqGdIjs8mKiGtpYQxJA+FtxB6yOVp1wsEemA7lot+FGSHZjC0LbCO9nc
g4hbQt5h0QhrTL4oDtDYNTe6f8dzWZZAWSwkWcthuX/izwqWRW3B63t530YK47LZLbcEiA0qMt7C
NQ/HFHa6OUzjIcqYa1gAfRcklJ93xMcn9yy1WFHaTEhA9JRYsbwXstKmPsUk36c4upC5YIxYquDW
8oaTltAzoWuTa7Vj+r9OTa6ZWoeSMV3kl+gs/+D50kGF/fAUAPcrr9bHQpWiCB+s0JbZSAza8H84
ADw0oLzcyXBlds0q745EHjynFnIqxkikOix8qKH/Jlr8gOBEuGXh4SeKFOMJoIrzjVIS9IanIgZH
LZWIxJ0gmL/iaF/PAU0Fb8foyHq6deuscRyWnSkciMfkVsbTAVvNR81hrF8Z9p1qX2CtkFf4Jdal
aeHJWhXJg28L+8zegeEPYlkLozTafAzKDbnQI1RP2w5hkSJXkbIznKGY+4d8Z4Sb9ggO1mfHnw1L
SUUNI6QjfN46VxZjukqHd+vr8A6TXa6+YUNjjkkCWYzTS4Rx3UeSRhzNFaw97wdNT0nI3sh6icLj
PRxCidM+Ntgoi6yL34HgbTVfmCmze7EtLQf1b357uLQVyuM24ww8l4AGCDgH9cTThxBIfstH7WVa
OzBxaPfKXs9sKliEplFWsHC7rgoHBSbpTv/me+acc26c+yCd/C6eWUBsP61NJ+CQa4tQxpJIwfUv
k804q0hoOOaWdAMOq4bKS/7qN8OeQg0MMQGdV1X6N8d3qKvXiDuRDfKUtqXWaXFtqhK0cGr6iO0f
g7M9SGhDYp/AruJVHpYOE+kdaxGLgnaSv2Sju6udyO0nBJCqeWAb14KjCN3RR58Oi+xn7IEOZaQA
llGabOid00gUzkfvjl0868ZlFVldVpiIXjRihq7GszMhu0qe4HEWiaHQ1liiN/1/AE5FbvTBPdOI
WFnLX4ozzqrsnTWlLhG9t2zpDDLfzxzzpntSpndW35Ks/wXxk5qPLsldcSSlgHRhNPc/HpAzVT1t
C4LP8RJRJxbhCsdx2545OUhIRC3ERdZapnqVJc4RE7gDugGYBiL3+4DEgKAjJgycYsCctYyFe8X7
dpLg91Hx2/IUtKBdUacgpnptxVeEfkAtfF3OIPuOwnkzkU/p4+r5RHghvtxNWFpBZXrTjDSUVp0U
LifTqduIDMu2XNaUM7soGE7sSSSxsC0lVKW14KGJUTmEb7aYjFE3lAQn35+DBzuD38KWU+BiFhlc
SMhx48vKQ3cKCQCT/5gfLuBZZrNb5zR+YuFsDiTCLJVgbsMIN5Ky6XMr/9YRwntEkHiva11o0mRA
QgX/ZMUqyDZ4+4yiojtNs4pbOpGUj0jqgDaG5fR10hqsKiVOBxCEFK+Kqd6IQIKy50G/xu1ACnfw
nTXXrMerFhoYif/IVJ4whyEU2QnXsJEJ4qz9XLxsBtqyAjGJXcZV80aBroDQ2DyPnWouldpq6DzG
q99rGRBiUeoQMRLHTQ4wMlaO5iT7D+AyqYYo5qeVM1uyrvFGKPBH7tdFqwNLDrHdnTbOr63it7ts
+la+AXYQP2ZvT+y8TnBwCHi2vVqxdUBAvakIAq4hZ7/djAKChUZlantXjED+zX2nc2RQkMCC4sa5
7ep9gtEyxmwDD+EffbFQ5Xikrd2MrkeJ8AO+O1cBsR4oY+oJrfCG7p2+77lzL4NcG5/Hhj7Yb9/i
ZPXVxV5WSUabR2Yhkl9DuHkBryMo00Tv+lApQiKy4o6xCZtabgo6YctIRSacP5y9sCcq6trIplZe
FSNW54qMT58HcVFd1FxUTN7YdEZmRysADtib7TA1T7mMmk+7HCKmfOHOEtZ6fGUDb5jBwWZTn11o
EcNkb8NNXHDNmQr4Jh5/LmgQr2p0CpQ5dbOHAsrjCNMYWJmeAg9oW64GVyUZ7uM/KU8LmqWFAkBt
hocpSw9RR8HDzQIGVzvwTTieJoLRkK4SA9DeH6w2ccGFWX4E2//xxdoMJWwIEPa9Z6KD/lfhPcP/
ItKzB4oZnXJ+qcas+vJCpwmWt8OC7l71aUu6C3P+EK/r8x2rL1AlzlbPg8oZHt9NEk4yHG9gBMJQ
vFMNxAlEFC7zJEAgt7Kij006L6HkRqAkFVGwWgcR+0kqrmKgQnRpv+EbIwfNGKdCLuFGYyIq6aaD
/bCZCH36VGAc0I4Agxxjo0J2haZveZTKJK4ylZzQjSRMWvlsrZBfK639k6uCF3vZyEV/06rMuEWG
JcgJj+IUNLVCWdjQoXuEOmGSRu6XSvUHy3cU5xJlIspw7wf1a/YIVq3zusrD6zOW3X7VFmQy9YCB
qSceX2t4usdBowHZQhkt+iM8unX7k+Ic79q4KGnrLKpxlC9i7fWqVN+Th85Pz1qHREfUYCmlsKUa
DK8OK0Bn+ATzeU7yNuHUxzM2Lf0m+Gad06Ekb935JlGtq/iHjBjuZLYxnK9O6pxUM0EMAfZQt7ML
lJoBLBaxeJLaTCxJrIBElYsJW0e+cHS/ucy5aTZpON3CELc7H+VmUf3ZCoqz/Ezfxb4WEVcCzx8n
tVt6A8/bkr8B9tYrjH/TviQMlRStDjJiQz4V+pUSq+EHjRPhg+Td67I4BiCTX08MWOLelHYRoujI
3WNHnditQQ9QJaoStESlAVl6U9GYP5mZq/i2TuA+s+l2m8u9MXN6imTTNzS7nksTv0YLDFmz4j6D
0LKqEsaSuR3nLns/QunU/P7DtUaj+LVC4vh8YIOAi51yICjhS9qA3t6pYNt0itgARJNcoWswh1yQ
fcdjvfI1xDia1b95crH11N4/qVZuVl+f/iMshNs0SXWRN93mRsoPn9MFcpSGeanj/H4IY/WEsYha
9ataF9NDh8e2l/WvvKnvdEqH5qVGFkkDA7LnKZ8hSY0sTNoM3K5MQPge5Z2zKAs4ckCEV6AA82Px
YMZlkyFHF6u9B+0W3KHOhsHGZSiK5TOIPWmJaDgUtgGPqwOMMkXa6jEwyDBvgGYi6CQYsuxwuH8V
oK18HPrEV+rWHJsMV37ZZgg6FRCPBHBCFHt5CybcC4krIF7fd0eqi4Cv3uN+z0en1lH6Rw/z5w5R
/+05qeiF1A/casBPCXu89bmTTB4O3f5/BRkhpQ60KKpYaLTJOJ0yE9hNda4sevtwACKug8b9SQ18
xvkXMMHIMUAr2xpdNYPbVGLRSbIyCk3xcVn5UBfsuYcyqW0OW4yTVIddJvgPi/Fi+RmdmjIrgO9f
KjpsM+tHRmCP+f/ULiHPAITvTnAsYGax9jpSQZQXGeD+Um8I/zsDkPkgzVwEq1QaH0rkqA4CXCMv
EQPXsbJuvX24EvV1KotQ4SGi0Ew9rlZ9FaXOgDn9LERneqp8bvZsegTsEpkWfM4/bxOGYElrqrgO
Q+aBqyfBe6wSzrYPmXT6WM1htcPhbACLtK6cpp2z9wnRO1t36j1pttTXOLnFz3S1rDSzltYY30Cb
ksL+vJHVmAWvbLhdZbGbSdT4np0s4CY/fRThKzDsEMasYZ4Tuo7wicykSqU5m1rUjAvIRIeprvb7
48OPweUJrZReaJbBK5W0wR0osCvuiDPct3DUpVvzqqRCwEA3GYZhZ2CcwuXBM47iqmC/mWRoXHtI
MUlU0X/v3AwgqFg3xQCoCpgIa4n1Zk0dHdcye7wKL/tWTP+UPFHDKtATQtieUMoa6Cc8xcbPorAp
fWqytxie7HAzXxKyZKesdbUG56WZufr70TI6NMv2HTP52/ScoTbuIk3bIPMKzPgQ8x75s4fcXs4r
XZj56m9kqicgxeD6gzkvBsknNuf0fqGKiBcbjczPRad+yMxykN79fJYRfVHpWkPbfMIL8i/TdOK9
0w5vDVluJsJ9sjGN9Fw56lEVt24Kr7rAq7+Uj9VD6VVNIQ9PoufRnTHQKSC46iJ2Oq9VnBxjtz52
CCf7I+sKK8bLiQw4s/C9qR2jKYD2j+kNtAG+V0xgk8J4eCCwRZHPASeUDMmPiQZHAegTENUM/vO2
/kagtx01SpLo5eskBBSyKp0VvjRtLSiE/ns0QaUurvzntmXsJVQvgJvzggr5EmAQTn/tW55N+EnQ
+Q3h/eQ+KcK6846+vdsFc8Rg1biPc2BqbLUZy+7AxN6GnGhSw+PxVWqrg5pjWl5hUUP+8r043kfS
Lvd+7vMV+9VfpR9GtT41hUyfdbXVmAeB89QrHqCcynyF89Zj8QxSlLv7xRp+COPKY/VXyWQALxoP
sssylXlTmd2NMcGzFx1Uhcxb2cNFqWt56WG7QkAR4jNTydgTe0T8U+E0AlRoVEyAQ02+u69N7yzl
4HHAWDPVkEGE06MppbiwIJIVjWXvgZ8fvt2Q7zlVVtGnTMFdWYWfUWsDGyrejKsvTzjtR7CLjJJ8
iNihgZKUPjIYlxU4akYHyOGTKTylotRm5o5amb09se7Pw5JO0LhL2S1Ow+7xnJSL/gv1gA+cIhcr
UdX3EnkRuqbwdJqSA1wBXaq6UkCOQBr+cjCguozgnFAsAJ4Rmr7eiX/+Tkjxr36fXRmwAyxNSMY0
rs4KRKZYsbFEfI2BqR2UauNvd4IP/nDincpO4LxsEDdACPWtMnSZ7v3mRNYRfAnOn2jFkqP5pKy8
GsaMtEAzzPecK9vamQGZHTx/Th/7kkYmB275xoLsGXTgfncOLnCSrG7Q591kfRU1vvgF/hk2K39H
MyTTwWJJlQV8BEFq08gouqhJalH9ObQuaGnG5XwgDWCvt9nl7eecPKDFGPSyjAGUBNja7kTHNamN
EEscd9Sqpj+mZAMY0UbsPEWnj+tiBhKOt+yBJfoxUu+j8R7E1hOOJhuuWePbwCnyXU1CxRRbhf4s
+wACjHcvS1VnHRm4WX5ZcpSBLOwW++0Z8GDUNOln56cvnVII2MqvBo5V48fIBb+m6Pdq90Gmxccv
a6vWT9AjJUK0aFTY3v+4eYIL+P/OOvQ/yCx9J7wDPljMNj7jvPkOZHtuZqxe2MJYYqEdg2SO47MF
38f4bLgkx6LCjCPwfMayjXWm/DDzv1N+5o1B82Jw2bqLAmVNYL7bDdEaCnAs4gNyic8JC1kKujz3
t39lM8LEcqMjibn7Rzvqx7OrbdZZM/MaXEb3evuJSfzeCAFDm+iEK+xAvQmyVNR9CicWytkJXBZG
qnvAbngpcKTM6QHeshKDDxuM/d0PI2giaKeZEGe/Is79oleE6u8VqOTwxg8uBbf9BEu9K1SzSYxa
SlYD1bp9d0G2CtJS4mQX9q8DpeyEKYPHBwvVjKoPCiwMrOZKg8kjMzZyg2vpdFFz9v/vSS0fNLsx
9apVU3ZPL0KbH8rFaGrJ0Jw2bcby1nQbrwWsexzJVX8ZpobJGHjQ3eDPM056tyx0eWt6nPIOlLMR
OK1msec8v9zVlhD8FhSkwoeCc/wkGgH1RzVD0O0cpsBpc0ZMdGeMiO5asvZPpGmYOcIepNTVZiR2
D8COW1jVoiIR9mOoSAD+7dTwMg/8IqCW1O/+m0bEQBIY/wU4rcqC+aiLVGnieZZChCiJxeo4vNqI
AWn5QNWlzF15CuPjEIFY/YML52gACcZAn91lBNnpxW43t6AqshPJovBgjXbOsxncqiZAWN7zVTKM
rdy1EWLLBfSUVuEYDTe1ewbeDjmoUF1ECUnEIfDi2fsnV8vE82iTfPrEBby4xu7eAwnA28faaGXv
UZeqcuauAZH7zMboZveJ+Mn4Kw6rBfzKPo/rT9Anpn8cRxOVckpQFvK+uGhzl5nQnerD/zSHrIrK
AyJWYzT8voc8WWHgz2d4A5bNa4+YPqHE6f+Su3b7BmLUgV4GRUQOkP4hYUb2Jav7w3liTHtcx+hg
3E8iRQK5veWHE6RhRdg6dvxWhaRUxSRsywz8EACUoZbyko5ZQsI5tRJIxlNdCiAWurxSEOm1YjBL
+viC6rnmXXQ9EeJEmsvNa+fLULNGu/1vEBK/fa4n/BQ6JzN9vsiRe2geb3GoK5BAwWulzAmdroyF
CMEdOW4fYsEj5CS1DjgiXhs/QaXZBcXSkSfe9NnXR8dHORg2YLDKjb5u0dvv2S8rH3QbJHQVyzLP
KCY4yRBQ6fJiv3X6Xgvy/HeHmY3S0KCGJspXGplEzWWXHAR+BtNYwsBfOOlPPG1oxW9hsSn58D9l
M8K1xzNUP4dWJdEmh5Wa+Fv9M58aQkbvPhBRlSx+yqaGTqyVaOBK+m8CiRO41LNKyycAeVrhQUdx
PeCvcRtU76RI9tHtFJ5TpbbLbjXo2YHtMfadjKOLO/B5OGzWAO5awvliYRqiZaotiEMSYBYVE1DH
uX59SC53fbeH2pHCHdBhlfkWrsF+FgbF+ogat+kFr5DJCyDhu4oCqLYcY+LDHfzqsQME2TCqi9VK
UpuCJ76cIlXPBJa5qn3olC0o1rXCwaB+rxhCPL8UmwL+fhAhr/232oXFEJxmj+KmH8i8HfiJOpAC
Zj9fIrm+A84JS4OCGzHJkDFZKa5Nkq70OlrCijVVb3Xrg2DcDJd1DV1mbzlP72dVE0Xb2WObKEUC
jXHVaI6HrOONyNzRPC3m5iSWcobyoNMkfuJ2GSsl0IFxUKt/k1E2dL9fo+WX5iqTH4FBpr4b39FV
8UNuuPZCgOEcgnQzznqZbgwCEtaeZxUhT+dAFYOr9Q0oMKlwZkHY4Fekf0RQOe3Zggi5qAwgT6xI
1/FSh/7o+t7aKD1YszRCQUBnoVXxDZjfPKktFpymbNyGpWoFtdIBSFcGjuzN1HRcNk52i7ATkQdN
VoN3Qr7ykxrO/veyx/om46KVe3F9P+2Q3XiEvccZ69hBa0VY+FyoI/PIbOYCmxvkcP85C8uXt5pS
XghThZIaGoz0r2Zno0oYmv7D9giPSexIOtF3mcG0S8A7haYZIoIk62x6b+QvUHxzXc3E8N6kcrur
d5dtgBPZ3ZGmKBWS2swTc53v4vrlXXSUAQCDPpF8FC6kiaqreiT1/E4qWDPLe/C9EjzYiFIRqCQq
c0VK+S9c7Zw35XMAveh0dewIlbS8uY8T6ExbElckcu4mRYRAzE58kFH0cWgxgZCdFjT0c1gO1AtI
aq4UaJeKSfwBkoVmw4paVLdnxb65cPprknG+gwKAOYO79010j1c9UaCdWzILTIMRsqANRGnF83bB
Fy+cJlu2cevfMghFgOkvoUZ6c8evcwd/2YTuQWWwDF9aoO+XPsVYmzQ8HuRvN5USnYbv4m5Fm4kV
3LBSiltuDMI1lcBTz8qskVAViUMFWexTatNnEMCYpTnYbXu8POmtDUMPqzzNazZVBReQ98AtAJuX
Z2a7xtT9lUhEm1ADOD9PM7+E1TXCis9Ig1U67NkZQ827d8oJ/MJDGQrcuESy1PWn9ifnWQj+52AX
AgNa/25Ar7L7QTDHAWPwrE1thNXLbHcuMzhH3aUP74tf9qtonzY9TvtoXivSxSdeRpp9zgSycGF5
RAdYOlR8iBnWkutAJXHRWpdJ8hiA6ccqF7kmcs3DD45m4HJO2OSKfal07sm66a1FiyboyK98qRI2
SaJcUGCcsO50omwylJimjQBukifhVGvLEnHhv1DSmWWR/MjzefUpbwZhatPt8mlUOpNSqaUN/6h6
DojG8/AM2cAhn+S7FnCSihS1gtsBYP6zsOGhApU04+eWhTtA93W/YJGkncifoIwC1nlddLSkTLT6
PKFTav8ai5YXkYOzZe5G/q5UdxqIeU0mVy1Gbq247h2qxN0EUyRCHCW6NL5D7YaZQZ9wdT3BCAmT
cxpAuDMkU9unb1VLGN8C0BakXSoz2nF7Sqf3XMrlbbqoJhU+FTGGaoxV9uuaEw8qplCeJest8CCv
MLJKAJNXXD61DabEe1uZgpF4JJii8Hw+nglcUn9qHHpAOJgQtM2CkwyjJJVH7kh4Rj09bjaasAWy
4YS+gvMkssAj97W5XRGgYCnKJ5CDxrfxjj6HR/atTVqJUQT4Pj4aL8zs+mzGHywp7dSpWbvwI178
Lu90XU4RNN40dEsk9T+qU7VFysEsZsNyoqzJTNBlJ5FAqP6kKvyzqkrDYUfPsZFAmRRvA7CPSXBX
OcwevFGjNc47hMDEv+FRRsa7OB2X+P75a/cHpOL/TB06IYXBUnme0DwBgie5+9MAMPuUDjRECpQf
McCc3Xmcd9ffCMMmWBzb2kY8ptLXrK2UF4UZ6V9NFX+Uki2Vs/58HXdNNnUgRhjaAo4GpMVFkauJ
8PlWnl+81N7JZZWRQBxH3gDbtJGJjTo//0fHxWQXYRPnDQACocVDa7k25ef4rVoQj82fr1d779Jj
wkYmOjOQ2uH17+E12Wp0eyziJgN6Tf3Fw+mYh8txZXJQUTqWerFKmnPezrIoaw5HuthUtFu9/K5r
gxm1kTvMfe47y1pgyyxbbqAKuIONNzj4ml7ETxHIXrYUBxZl8h2/CMfd6FzHo/0lQSoj4TNcCV2j
Gt01GDRpoI7RW+7GxG7McCpGzgWHtfv1ctoxQ08wJV6qOf5RBq/3jtXne4DX1ONGNt1QXXnXMmLO
hSYSATiSBq48gedFIfgrdr4nWslE/JlJO628g+GQ6PCAAwkragvY88eSSk4kneJq2ydE0ftV8KtL
+RvadUzO/ordgQOfpWXQZfRGHqCM0fg8M+t9rUnWEtjnM/XW/MY2sSROVsxNaC16WjlHcmdJTk9E
uj0cGsdCBlHgl++E6KLYtT1Hx6HzgZYZlau4zK5RQKdKRlKmOllu0RDbyb2H09x358t1mZkYaErH
GnUxH1qcq1lqOUc/Doo7ZhwlOAF/0rP1V6Fv49HBfc2FrJq4fhHauqtS1fWFp7nJDt6163ObQIzr
tbw/YSEviFyZyA4uu+NGxk8MSWmizEXUhlfZHEqteh0tD8RQk0onB22dOTqLsqz2m5fpMIOyrdRr
Ksuo04L1ExFs7l6LtPPgVJEJe6WG2ecDB1m+aRvE5zKVXmN9bRnRr3aUhtvGeEfEJtpbg5gWiY4f
jcANryc2Ga55kPqFar0qlS6BbViDtlZLv3e7Z91d2syzdyL/C21ePXJ+Vdq5/8VEHcqu8xRYZswr
1IL6naZfCLkVP6mtWkn5+MgmrP4RI7T3XfvBplB9wNklYQANXLkOow9ZRFRVc6yG0DMCjOAb1d/B
7msGUlSqNMH77bJWpYn4mjqAMgVMOy9ifN/CfkRRnbWIfHR+XtGT4ivMx8tavMRta1AVX+e7yJ7B
93Pjfrld1mxjMA5Q33klMDEdFLD8w8OX/5frWvn6xbM9w7Ysyhobww+ECk0tbiWAVBf83AZRhCwR
W/UfCKw8rMdQN6uQDsZNkLzqWw4DhhMmT/K8w0RaryP8juuwGJDLaqEER8sR6mNagIG9b0/Y38jV
PzVg1xtJ3ZBYhYAdB9+BP8WUF3BbzDU+QNIqG8vDkk+hMCQ4GPlSaZ2n01EtMvqGLsNCArtYgl1s
Gs/YjSe7W/W9FxAalj/MzRicQRRGiswgs61oGnPIfOvcwLjw44gSdUh6+grNHaojb54O0j5tc/E2
+qoSFIG4/fjmmfv1J50fVceV/NMNEW4857teJKiKm8sFcRvkuCnv26fHFiu/7d5PbI6dEsGhb3MT
Yv01o8oNNoXORlbXhAbqShamAifAlSUgA67dEkWsyNu8y3vjsjnfF9ou3B2HPC15jLgGVihId46Q
8YeQSbl+NDa383MG5Lu5RE5Cn25Rgmi7UihXQOEjMC3ddEifMlQ9ycjHOMCmwYG4tfqE0BGnUirn
k0teMYD2A+htSv3s4XLCBc7QM6ZSSAC/WOrbpxQU6QwDjk6wUV5+buDt1cXVuSihmyvrXcUd/nw/
WgY1eIAHndRFXc8/TvRSb76nqZb69tqbFqIyrdUr7mJTmx3+oqrML0Y8AXaGCPJ0Yfdhv4OlYpQS
V7+WXmeNOQLcpvKO7rs5DhIEYh6pgkG3uGZ/rMyngMqJ1eykKU/BOeREETVFtgcp0LF4nqkzeJWm
yhbXbN5e6Vh2R06DJmbpez25Pl+aymscMmnlozwriNTcH3GCg2A0xLlvVdNB80U/6+Jv3mlm0HCZ
GOUtzlcH9nK5V5byoHUAkMBwLTlHsIHGE+brVWoHBI01de8IM2wAX3hT2x1kf2X2ySypA2FKXCfZ
lqmZ1j6lf5Cw+pkjQvZRVNrppVk9bhV6isxm1SyyrmPc1OhdfX2NzpGKXG5egmCfO6yFkY4TbVE9
Y9yGefWO224SQtViRcsV16aJXhUG94wnOUXXrJ2zJN2wawJeyAOJz2xyeyVcEKPhvmtAE66znury
pnx1X0bPMvUbP2pZEbHdZzNC56D1rjns91l5LHQPnGOFIHmzZ4OhFEm151DMEf61t6CuBdMw6H8E
grS+tGOY03AXE2I0forvGEaxwC3+2Wo7WMZN4EMsGoUX7FR7WUFcci4M8Yn2/wEGHppfctzslsa4
YPVJMJ4ix/94vHUpQJsvuwX3NaRf67G2K8JESxbSAK2m0V4DojPfhruAS32A9zr+fMk1rAFW3yIb
E5p7tri/FY8TbiBLgnsDTe0LGxuMTAhpDDrruOnl7ECwOSSlZrtgmCgEUqoS/8vLPZ2QFpVOlnAE
yZOFoDwhUfWrMh6cAOkS3LzCT8B5E0ZS3XH2glwdYLZay59hdq+xskT76IU/WkL6usblsA5fZvcF
j8TkZCxYn1ycYdFOl/cYEgSu1VxAad6Zr7pBaWOASucEKawqKTkOr3AuCjGMmJBFqMchqoWEhljR
Ep4xgo4k7MDv2Z0IDHnqhPICzlhHIyy4YsEr6gkjDncn/qHJlpEr2wA4B/W6AquEKThg70AFlVah
Dr4nk16LayxqOrJ6hfQX3bjwANVV5mu8+X/juN8rBdDNuL2po+GpZyLVBBN20TR/LKJIIlcHqKCl
fYsqrX4WRfGA7EnZAPqXpM+WcrIjarJdYGTJs47E93jc5Lbo7CL0Q5KM+0nZEikNJR8/6KiCB2Sl
K7RC7QfpmFm0oq++pbbqbzX2NoYB4QWCqt2kfIAbVQlNYiX2UWGh31hF1IAm/wnIL3d9S8VS1Ffx
51Clozx6XqLuZYMvTzOk3kLNMyHf966JRVUKbZAZfzRRDZp59IoVkuynCpT5lUuYQ8nSyTWFqgNa
xpG0AWvFkhVqoVD5kbabQUoNB0C1YQrQKtD5EGIBqxEBXQ0YOb/xjCrRxMajtGbGn1XxitgNSkKS
wfEM85v7bu2q89Yq/XaMP9+3NreKbX1rNFM3YdpnpZ0dBAxhgrkmQQqHAPieaVPeySb3XTvRzano
JSx/JZY2NMOZ6G5PpRnL36YBARgZANmDEr6uRLeC02WQ4I0yQ6JPQp1Yp7vlMR/zSR8cA00UqlsF
BkgcZ3f3i4ATiQTQpch5RALG922vExuXtJbaqWdkGMaY6NeTAd6aQy0HX7bAmJxh1jVHFcKQdjEE
Qa+cWnSDpBDrsd4iK5BzcEY/QLLYVsYDrt7mIqzjOXvRLfCx3ydFFeD0m7JWiX8WZzQ/plYlBshI
R+kKwJcxeh0fomD9/CAiYYfNa1OiDEz+++7XitBHzfB8DY7NVAJNBa2mqyxxv4dq9i8Lc+cyMd0j
mO+v/1awTgwsE0eM1IGf7bzveqwN5eUrk9iTrCUuWdbZ09rAXJkjcuogEvb7PfaDQ/zKDamlvn4u
rnY9lAAbvOsDsUy3r71hJh8OT2R3ApynirDzGLcEV4EucZ0ODHtFby77NstCvU6RVWiFz+jpF5f2
s6PS2M7SqffhZlvYix90FooDHGxoop63r3/sK+lzK+I3jb9uq0m1FdjFtshSsT3rL+oseLPYgf9S
FOzOMBjUXa0HMfO3a0zhBEvarNLLLbjZS+/WUXSz0TuLvaJzpPnRcpHGl66hm21QZ2b6WLedcD/+
zW7cI/rUHOSavgsNDc89v+MYQWMa1KKEoF1YTJppmhkGxBbcs7a3TvYidFNrZnsn4d+I8Dcw1C7Y
be63eP+jyvGw3AgYA6sbIxv+xeKGIlG79mz2rmzW26zv7Zw+b9svtoARlcu3KduDWFdyz90xNpkv
2hiBBqXKcaip+AgU4ig65lZi3wgUpOHTepPq9GHh6MP5CibdqTf0hre0xzqkd6ZjF9GarH/bfNQr
odCoCBtf+Q4Ob5zUpXwgIVBdpN2Qe8CDIh3uuPcdQRYDMoY98spXGbgD804PzaqFUicJyirkEcvg
7P+58Y2gvRAosSEsrmRfVY6+wmuVKMPMgHb8g9BTzXCKqKsFoSFM2LN3OiGWu9qRW9kqntTgDZWQ
JxTLICkULbeEOfwbI9oCKNeWZmIOQpmrw0+It5dzknIG1hCCJxI0XAMm7vSAklnpkHKb9gfz9LA2
0YqGnsikDzpmBAnoC/XPQv9l6UYAKyt4IPQT2KPQ8RdnxOwcoDBxiNuoKbbVHFPuZoeDZHSy/3JM
9u7ydfZ+RY4jFVOqJl8nVru7OWy04MRNe576zxRUOPeGRbus/2tOjnCL3d2E2g5hHSd25/ygHUnF
1UtIYaK55mjMocMnxobRYD4P6iVWtaYvcEVsHnhEjv4zxFemaarTJc1bNdtaom3tuDKP6pJFL26T
yKqfVJ3Qh/3g5kxh4l30o4q7zzx0sRfM8q40SQ4Z1prftm2/jJkb7e8C8ch/Ds4HXYVNJk0CXkKs
vSVTxKe7nrByVxOQGBmFkOVXIRpXsdN23P6iU0HHIik7f1fPDZ2nGO+ja9q+EVDJ4B1NI8owBm++
pMMiNW6KVzQqP0Ruv9u4iJ7YF/Qc+/4BFMsO66n1pzHM9mhFzeG49DvnBAXYgpmIc+WEL1Gmbg3w
rn0Da3YaljCuYcLSietYGIDUbGl3LR89QPNnzpTobWyQ1nTUMTiOv9OTBLP3oyATxgFK5iZfvfP/
OGUQmkhju7Gk9btxwfD/WqbuuuVd96MxN8cXFeEKkQBsyyLdPI7cIp1JrRZjxOXGRf3Ud55Gnlr5
6/Q3lb83Y+NHplyRtGV8z0dxi7gBJd+nGyQkiVBmDrtLugUIyTSdlkxoViyjSVM8PIPMJTyCaiGE
YzbHuprUBr7wpt1wgRuwYzQQ1ZKWfVSY2gHTay25M1uUlBBvwv+7iYLil/U2GsIDRhtwPQXShslf
sPrAlC9NdAnIkh8dsevSopRQaVlK6xWQESbjLXSjeDlZVpUA4qzZPoLrcgWGtNM1LC6RtoyzVlkc
h7XpfRy5CRwfx1aL9/n7beMPpEtlxAhQ3H43vjx2KBPExCBsAWoeu/81DJTs/zqE1hWioeNlO+gi
TWStATjlFU2m4PEQ/kqs9F0dAEh1RqQLqgGVzA8s1PNLYQMIanyrHKPulx+cRki2UEhrtUVLqqZD
e7/Q+cGBp7Z+8oyVCh09PZai5JKn//Ex3QYHAUpbgtniUmVelH2BVctDAAXY9W0OFBayzoAfyraa
ldBXklOC868pE/Jlo9hqEMJfaELe6MwWDORBJVJkZa5YSz+YUogZzBohVWXfKllSplfsobjJ+53p
AVYtu5l6iBuOIHbHnPJOJmbbTgJxiElLyWvhwqbsH5Kro4D+I2fRUAkoasviFDYi+vLMRs5KRfsS
2hXtgYPulA897PKEXrDcDFal4t7n0qnsmChAS2rzFUcPqbaxWO6Fv3knCllW4Mn94TJYE4ag40lf
lbL58/dmWAth19VUc1XYRfi6VSEPyYtTF1N10N6uzywkTVcp0VgGI1y/GaxMpiKH7gIKy3Reo6f8
3Re2gwyQgMC0eEBk/e7wUEW05l56C9j6MNgMTKhPwPMUlXSYDlBXtbz4+bUD/roUyrIp8LtMtGHB
2kceXNveJmEUuOzwOzo7932mbB2LuK7pgfEDwQuZ5w1YJkbu//B+Z+9GsLEY5UcT7DaCi5gBdlTj
2ut9xkiLtR4bF8ZLXRN7eVNl1KZGqMftX23dR0Q21BjygDvTEaHRbNo4lP68GSyhVQ8Yp4ZOb8OP
+8Mt01hz7qUn23T1QGj1iB22zBSwQFhjryeG110Hp133mooQi9x4sSGt8Oj5dnVhPQrpyFCTCOwF
coUx9c4cIe2kBWlIY0kCsvmDyt5v6O/XTj/qAo0gXhrK0ZScxKV/snmWrPt6+2xLym4fEetA2kZp
LInWJDE1KvICV/EffYmOVO5yvJzxaMYfvj5R1BwOqL3+TmTddlYjcSsnalyZpzEEr1985goMyIt1
yfnA1nq1oavWfjyNVR4o+NTeg3BzDpCo2Z1fKMB/omv4gIKwo8n48xbtGwWz4a8MDvanXKhARLOH
n9/fiKwY8UzWPHw4nS8aiTbkB3znkVx0y/A+M5YJqkhjNVJ36c05brGDWZ10uHA5s52RUoBr0X6q
3+9TlDrTLarBG8ZHSGZIek1xMu7RwajqZjRYBSDucvv5rZHqoaEAkF2Dow+Bk3mIr7eE1Y8GQgoX
8489VJnpcpFQVGcpzGWlRqC4kSIFevb/KdSTrsZDsbTyMqCHGWOkXICga8bq0uq1v9ojgpJF1oEF
9RTzd39qEbJtazBPm0i5cjMT46ADRclJh7cYjuGHdJl36wlHQ7sTCYauCidzMIAjk9uFP0j6Xj8o
/1Y2dKZ5GMeoJICiwE8vANrC8OunRYpc63pze+w7m1scuObjcUIuhyzMvtB5VM2nU3i8mD2+Ji6x
WoA2BZjhTVUpN/HqA6PhYZf8hMcRqQnmFdaOqbpWnchUrSV1K7N1GH/vKOG3whuholnfneskkTp1
NTCMlwJApSy88R2SCy9Djtq7nQzzFsNh2+PUNuiuacXvi8/2G/Y/EhTHGm2au72e9a/P13nB5Mz7
zGg5pZJx343Ln6nSjeHJuVuLQ0Igjv6mxF7TmevnW3BvdA3UeDT4HkPEij633WLmpxVccnt3fvOk
bwydWyoGxNvLMkvwFL0lFPJ9SLIocopgalRzfKg/1PZTGpa58QBCcpa3wSH2NnLoFWypOx/lqJoK
2xfMQJK+oPbzL2TnP01ey6z6H/hpYSdAsnSENGcivYsCM4S0MwK0wa2w6uOYu1mHQhEOUW7H0DJP
sCrnirfi5gr0fH7QBz20V65P+lSog5Y5Ccf327WXHc0sVIoFcDqGM1WGGpA0wNjNM4zg9p0VWlqI
zpTVSnGUUCIfAsg09of2hW8m+UKimG0Akh2hpfy7feqZvhh7eRjEcFsd2HR12Up8H7ye6KNHBbTt
OJpg0eCYg266eXyo1Xq2hFgex/KGGo9Xu6/hHbkG5dK+CLb9tyKqYLNSt8HNzLIh2EbgdsvmnlnU
5qUti9KMH7eirMu+6CqHOdxPs9h2IRWUnnuIic3WiXWZLoSXsKc9WkhL+6jPGQngG68LOJQQealg
mWrPk0cm0uGByKlkS9rmGeTjDdXTswINLMCPH7sXzRPMDxXw++i6My7+3JEyHmlV+cTZBSYGZEwM
bGUo8meCTR7gO8f2OsxcWs9jny1qNILi6jeYcDxuAiXnOhgTooeMdaZH4TX2mRePmVDpZ8ajvO2+
1gLxzHEIscXzLhq7gHF+1qXysPe8/kirklGgCdXufzcKpfGkY9SMHOhWF77b1iizFolvc6O6qXe7
DVWTVe/5Xe7bOUM4L1tG2gtHmbpb9uAA4CdY7iyYDjOGNrV/Pg3ll7TIpyce4OZX/7605kFsgTqB
3feAFLAWEGMKWdfqQkMMUXCNlAfOTYi7g8e2McQBkGrLIRLktvmOHarsZoh5dbMJNm2/x1jGM/cI
fkxThXfetz2bqfycuI2zNtM7PKow3D3bLfFfc28hRB0tOSgaH/4G7bAGzKWn5sr0Qk5in3hG11Hw
s7kkfV0EKSktTuJdwIZfYZ/mTMcb3/Oxv84svz25Zt6Axf8d3H+5nZh0JwZKMHe6Jyu4SxVRqreA
iSBX2g9QmI4uQDKrzs8MQGeanHsg8Eml1lqjjX/AtRu9wwtVAypT4QtzNs5uYp9rjK1mvevHOL6y
4ebn1qem2Em5E5lhb9CjZGdYCtgrn9W9y32RYWhwCkx9V7fUouJ2QyiRZg55JXM95m2i+SVc/mf8
XqjGax3ojt7RAvY4C6dI3WImCH8HjXhSLOe0urMM6BDE5I6tp++MrWMhRI6D0T6jtaIpH53iiCE4
q9y0affb+PPFCUacEytWNGtSGC9UDjwSRJQqFdIf+NJHp5xskrJZ42x7jKYIXdrkcygtm4jAB7lC
wXYja8fMhKEs0Lacm6hMEQvuTIwp++qxbf+UAv7dKs5nhkYl8hdiCL9hBI4OSexfDXSE+Qfv+vSe
ahTAQmqECxIWpTRi3yAeTzQycSUlpsl7QF1OgevqHCblnAP4MWnm2JL0ktYjigmAnlsjKtzdD5jE
soHKgeTGI40wOFcnvHviAR4NnxX4K555PbYewcTz822DdOR6lKpKfajaMWvJ8DoJZPQyfc74xZ1X
jwCa7ZBVxZcpc2ToxKkz3NlJqbx0rHUAELUtj4Z+10hTj0uwLCPrtl8sPN33ZAyM0zNo+agCWdXS
fCeB4tRwLp2LnyAQhjD2Zfd6FCDdPPfHQfjlGWO/vM5Qq06rZBhMbK7cCxeAUJhQl96h4UX2EsoD
+1zeAd5IDTnYrdVrSklNYdJigwDVyeraacD18QBRWUOT/SlsvKO/ey1RE3BqGUXcMkTK/CJ4me8I
ThTInN0mURZ3bQw3Rec+nWx+c+JG+jjQ2f0ElfKZl+qd6TIqGsj1E6gY8pI0JNYmKjjA1wlRYl+F
Z2rBvYwP9wbTw3l4v+IVobfbFRyELfqdd+XP4kKr0BflQHaHyBcqoMfgyy4rYvoosC2sUi6T0Ogt
y4JHpGm/mIcmnNiqoQ6DgmUlSrlublNT7wbQgyn8y98Y8n81c7Ayq9MmgJ1U7NMEb0CTFbJB0MXl
Vfz7NckuJ/POl1o4Z4S7Au4kOP24nG41tGk5Z1Ni2fhxmGCXc8rZ0lh5MbnJoCXL/n8Ekxyw4s8j
C7G/+CKpV1Cfy7DLXOWFfzUxVj7XjOiaCR327J17beKOd/+/E/TKGU1ddWzYdLft8JW48PHcp7Z1
+VVLYfx9uZ8z+3E8sdfA5NHaUN6XyIYc4PvBFLudYRKAWKMC6rVTCV9w480fwAK4ngKXvz4Tauss
vDJb1HQZQbIILhW3yzcsNUehLu2AjP8TeI4i49YSeWLlY/gYDoDMurSVIpa8ZpMzKmtcGGRH00ew
Ifr76SH7g3pze8zbQKDwRxvM/xf1aKePnBJbNwn3dJeo0zQiwHtnr6S++ly9YVncVG0MR5KoZHut
P3nUyQY7SeB3WNKRJQA3owd68uUYcYaUdZuEbgdtt8csIL8AGaHgiKBglqxXJOAhxY+cbssR1b0u
EHq0JCQsl3QKD8QOogEbOBA6ghwjKcYVe6fueJNYMKyK8+AF69pc2rxd9r4/YQVCpONQ3GfvqAxv
pebQfVbOaAoqacKvOLDIzfx9KkvzWghUA9zC19lXr94l6x+PQGXA6zSWfygwFZZ2r2+vzmXrFU5Q
Ar4dEIBG1yChrt50CPeCsFdFRiuaTIhALOynHW+nDAxRdPf72sF9la5ODCGn+27bt+E48gKN9fj2
gS3vv+eXmjuUp2vBLbL0ZVOmik9btLpkiltEt6yS6zZNzlbm19rKRBYqTLUPBf8VmCf//jsex7hC
2TVZyD6WI7SnH7+2PICTgy2eeKrkVUiMJ2miIAJKsX7Z9AcWFjfVDZ6ipu7Me1eYAKplM7Fv5sHI
lNGdcWz60UG/b3YV5agXX977gbOyvneKv5eIYbUox5GdK4V7ji4r10PaEAB1D82HZEDvGhiqNJ60
RDjXB8aMyXNXbx3DEhiaZDRRokNSgbu9Te/oT/v7xtPdGkZLaFqagiJSP+5oEtno8UzPpzUbchWa
kLaOPX7A+TqEfuQ8nmZmowuvr1TjHeHi/e/yfI0UULWc8HNA2NgSVo5powQ6QLfcZHle+BT9kaeo
GgdujK96GHS+uhWlx2KhxHVPfAvFwhsvwUEBSCT1l9BgHo1C96KlO4VRhDfulzUPUfN4BM3oeEKZ
/smobKfhahEUtnWz/pPCX7Lk0mM4q09bVc33ii9vqADbBiIljCuz3epPWGb3aLrLo+PkANOEGb9X
cV5BKR+FMPQcut5zu69/eprYdnoJhTNsXP3frs/K3tCiybrIfUGgetyeT6W6aMh6DwfhY5vu9FQp
J9+zM4jgo7T4zWi70YXU+idhr/kEckCz3tVf4Ekg+j/6xWsgJF3m+vYVae34WX5r2lOkRy2lbdrR
9cFI36qboUuK8tRQEyE+epfIUt8FYMCuprySJIZ66CE7jKui0swqk7Wry3ohN98MzZxxDGzQUXUF
GYHDkRVkVaqhSjNnnjgl+thUrAc8ykJG46TdRsSQzbQzdZbINrFViRh18VoB0Jg0Y5j4wMHsoI/C
ApunXtdROw1eUH3fn4jiCXgincEWmNPX9C7q3SIU1+X/uyoPw5qZXnrDF4PNnxDEE2lnv/7FdhHE
P83sDBR8sbOk1kOQuzVYNZ0llSLr8pfB8FU0w2rGW5cgEq3ft3ATlnZgzN272PF+owDSXu3Gco3h
DRlBoGTeCv+f53c/+hxLQrWHm9dkA6T2g9drkUIuttV3SqFJCWcETENgsaq8W+MTstT6u9DyEH3o
H1NmCuYVjIJ/bsMDmsI8B0wIrsuD2pMTfsvruWP4FSbxL1e+3fLoj/WIVko0aywZ9oub/Zr0aDNQ
8mhip4qYipNhYKxDxK9qDk2z55AYdfFVm+ykR2Xub2l0EX+6l1c6QgFVYXyEbEEq0LK3jufPTfg8
9kMAJnpDx9443eNMywne2drsZjTcV35YblP2cJT6GLROEWdYJNoSmsDhD3z8hgZGphUoQR6q1QUI
qbciM3LDNCB6pW8XqGcrUEe842zpPAizi81mTSNyQ47GwGhjgKmK1Ps1VoX1zP3/Oxc3mdNxKcvm
JmDysjQKwSSOGLugthgUMUkGKO05+zsRDu2xtQj3oZxxooccV/q9cbn8SbAXMiV8nPKeAx1usFzm
T8YQxJRR/w9cGnxryBlqnYD1St4OpVI1B+Iucbntt8aoVPH7F1KhNB78F/OG+GLUS6sKeDUM+ion
8uhRnD+N14pOJwnwLXyTRVi1ivm0sLhwzzazGsMnwLSDmBQxqWqPe5X8cWxmOuCyvLsyL7Mtq2Qk
aOkeQ2P/1N53EtzLcuDyp0zl/Mhx+f6dGeguRYMLDqmQjGgFZZmdUTSEbflCHj9DCoUsdw7gZjXD
d2RSJ2lZhdN+5ioeYfQzd2X4VnxzX4K0QwvMCwPUNtftxF3Qpnpjh2bU/mPCMu/8KQpbQwG3VmB1
INpxjuJTl0zVbFzA+Z5dKq28z0cxFMFr7ER4zckOQWPuKIom/3sN+gXaHRCjKj+mkMOJKzmFMuvV
GVhygl5DfAYSBSjb8kH5pL65pau6I21D0SB5m5xQ8EEBl/bHaKFt4LRIHnQoRkKurtlpXZ6Cv4VN
YHBM6AiCvpqQOx73yYuOYcF6UnoqH27rEtN5erbLt/o8c8dLYCXDV5/RA81leb2j4Ua/4G2n38n2
mcv4e2BTwodMFoFcSn2VfsgzmtbTMe4YA39rkzIMWi+WDZhbaBSYd+j98pGeCqqIO+03oZvmbFKv
EDcsrutRqozU0YQ5OrVl1vZTwKxO4N3sVBDVupxqP2UbmspUoHbZ8WNMHTozLy0ngTfq9a7m8Tu3
II0zsE+yBPFw27l/91oM3/Buslr3vaDuXeLn2x6coBy7g/AguF/G0SwhteEX+MzYWcSar7duuNCX
o8f6ypzR1rKswazt2I2vu3lHsxy+acVd5cuglASz1vFRbhJeTRczYzxoeD+O6mI/TwORE/6lyQIv
x56N05LviI7iQYnzNbdv+3x+liortxDUODFJmUYT9Hb2N9WBjOw/8HQroiwNVDh7k5s7kXfZCuJW
JyO6I8TwPHs+z92rk/zEWT1rDU+lDi2e4xYGLDOoAIXxtriu34QeFoissjFtJpFumMkw9HAKSH5w
OCzc1jO6pjFnxhDZU+KCVz/7ZzwSwTK8KHiSJwQLa6VHyXUSVqv+mnxq0RxIqNWNVdBtRsBEHBE/
M9WeIqIcrZoL8g9GothJ5FLhCAwnFbQEeQpXfzBDhwFgagsw2yqbylNek/D1Jy5oO3Jxgv7z1mzW
pcSYDNIGo9clPGgORz8l7EoU24xtyiW8WpuhuWt72R9j1RvWYX5KingFgJuGuiyZmXnZ+6YDOgwN
LDhI2w4uwT9hy+u/ImkUvR59DD1E1yaN9AOwmz9Q0ZOaBJJacpXiSxpGWGcsw5400ctdMSOMYjor
KBHBcsqcwNisbTzqT8zZTZnVj1vLHOH3bj8qJc9F7Wkh+DvVqXQfznrsDepbevh7eiuESAqrNXbN
gdXFwEYTULOSyq5bBMhzP/JqWXRdxqwOfLJi/c++o6ZyDNduedxw68UpBLnHWFV2aUAKI8DDsCVT
I23sMh0H4CAjLXGe7w/J19I87xSHJmPPO7JVDzHvb+5T7Ds1m91KI3czM5iKThe+EukObjBeYEhw
nK9fZ+MKCJchrzXPH0Mhv4DtLbiCx1Io9l0B3XPI/ofwSlOZqEuZgTpEYZRgYpy+tfc7eR1hmjzz
QPT5j/WvjbYhmtfZJXh9NAr8SeZPu+mzCQDDOX0ay6fiP2z/4qDJzOTnSoNmlIhfan+rACTf42Ml
ifTdc2/vLwolPVTPPJvZL14JCIj/DSKMkV3mtPJpDSwWWV/8cMGfvaxJNCf11vH+UEnSHlXaVVnd
CTWg1P/MZP2i4RcR2TGkGPSJYptN7vLAHSPkT+xbhXFBfnO0EZUvV5z+DY1gWawcw+5D4cCems2U
aw3xroqYn0rjDPn1wULphnoQ9wZOlHCkK9YEFn+sQf5/4F/rL9TlGNla65UFkNDT9j3lhsN5q8xU
0Ln4cUEGnveipjrWM0UuiUREVhFY+WMltn9gmqHt40AmSviP9VqCGasF5p43m6LKa1ztaP5DSTWk
ZjaMaVjPipD/njzTEw2y/01/C11qFDqJI2Fn0TTz0luBLHDBcBNIC3KdfQ2wEyYD9g23Mxwa1TFh
ufBzYCfPrVpwAHD/zbsI6tJHXEpv0EIDCYdD3zXkC+OTXxC6OZfmFFtmRJ6pX29x5wIwfYjDu26H
nT2sG8F8uic2N2vRmq5DZkLpPfvLJwucc0zsOfjKo+q7XYP36gQ/6NFspNO9YUGrc/GHNsjsWYCN
izxlhtc1ZH8WwFyJSftLt74GEtRWRwa/ifq2wgaI1qrKfXn2mwlWveKZ4LqxywmzpM1TOrpxhboW
UqPhMaa5l5W36KV7DScs8sHeX8bXNUCjCFAW0hv6T1DOxautDRGMMwwiW1Gb+HjZWHim+nxI0wD/
l7lLhUJO0oa8EyuBxZlg6Zp1/qTLrmyWiGnjH8AYaf2aQwdVN+9KY3y7z/YbiL/Nn1q14MbHpmcL
KEmuhSnrj9hkFdnQQW72W1l5uhaEB9IOvtvObl3UFougN7At9np1asLq+MkUGkUnCxkknqMty9Sm
TBtgfamAMBlPLotL7isb3eI2QxsZV3cDONVC6VOvHj9m9IsE10ox+L5OI3U2wdyL0j/+c8OMcaj+
7Mx9CLB2mEq0zjDxSxF6h7aUP+jBV1rOIa0HdOon2DKLC1jBgsJHXP7xW/URVtpnu78jZJDTl4th
McnMXhngVKEamEDFrLBG9r39LojydivtlbQ0cj0F0aHnz8P/lYMhS/TRTmVWIzaxvA4CmT9BL1pM
LxeUy8aO54/6BhbNK9E9RcQF/6hTM3hi8g0mLQWpZupcCn9na2Yj6Ce4xbeI8OW3tE36u7dMCo7K
cwGPtj5SBS5B0I/RWclVpqXY2vUNCVPao554qg0pBfcc5O0tOOjTuOnHXfhM4PGSfrBh1EPqlH07
zoGpVIYSJfyDTnE7VOqgzfDbXpBMaIGOAiymF69+tIuF1JAk1mgPxPdPUGDgc6wOHbIFeWH4DB3B
6suHuc7jMuTtGNSQjbLAWQfhhtddq0RSVFrvgqvb/DW0qelr8iQ2ez0kF4lJBhI2AwrX/fL7YTFj
1VNbXdcMhhPvQd6ezBC1eGX9ul/ofSv5bn6c3Xtlvix/bK6/PV1V098vyGXOV6Idc3FVvwBzrEsl
NuSgi1QfxzSE2UCuZiMqtdp/c9uDi7QBnIlZAEvi9qNn/Wc3UnSHpjhv77OZiZtH2pwl1UEhYVNm
w9LUfGFwQjf4QIZ5Uj05WiCdxcH35AcqySE9XWAfbqeJGdYZq6I4aZ999ZvfINbZ6SSGVGCelcr+
ITn8l0E7/9hdVj+QWGyPlfKF3DDRYw2ZlAyEHdTkxALkVhiteEuPfmXhmgI7Kt2IBlCGrA50B3ZP
o1VV1KFVHfkaPVJeUOpn5MEdflGuIwoWkl0lx6g2JhqvmlqofyX/txGzM4RymfY20HKp4YdWOq5E
vH9GRG406ewifkqWne0kcoBRK5SuDNLBavbiZZm3adTllJAwiHDrk3LFDPpK05lspnp6Iq/ScJ1G
RlR3i+/c8j6In0t+dCqoqSCwRZw6z8CJd9OEGfSZ57mBtdsoVh+nf/Qrvsj7Cf2YUrErRCWUQbYd
8v1qwOf4FWLr3WJXuzQ3KbM5ShXsSx1vWoFMBVLje4RetIUM6swbwKYOhYQTymguJ2nAFf6gqQKj
8XHBea23DewmIfoFh+IpGyb4MJDeBW06ydQFY1zlT4fbch9nS5bJlUjNOeecYqQaxMg09m/VBjCp
MWwqBniLZav2wSjEdsxqVuOfkQ17gUhfMkgpDmY6UorAgfCQoWBdCXojJURno2JaLiMVxPK+3BRO
SJBz8qmtVautb535W5DxRqxakzcBekektOriDwJvg44sHriyLSdWz4ewozs9kOSrkk90ca8rlA7p
cB8wtxlqB9qtv/VQn7Z1iUvIPb+UI52NKHX149F0tGBb2SsTfqxxatxI84vTeBE6ma+t8pgH1eEB
puQot1kpQG2mLnA/qZz27CUOsNmPjdWGQ2m9z45Frp4flDk+ySJCuXYtuqAAtJVplg6gE6yxyJs2
wiZLR9BA/jusTP9I3DChpsOmucENr8himPm6kaAWmVUTIuwsBIpf0UMiUjyOzxboie70ySBxXpbB
ZHIqTNXShY2umXyLEq155E8K90eE9T9E6Ox6mo0JGTDjtOuqosnRBd+a2koL4kzY4RWkrnUma6sn
6IRY8lKtM/MoGVgKogGUvxrj+BzC53cOkmw5g16uQ995wAsqSfqe8PFDJkJPQ1d62dJwVivsdekO
5K3MTrhvHFgNpgFgTIbDjpBkRV7CCOwWUliC5J39VqqBagMV7Be+XOBs1HeFPLz37oWWSvS2W1zO
2OXi1/QUOCQhDW2DDE2YwiYdoz+h2UMw7Szne9BkBpsLdgZHEgn4ma6y6eSlh5wCLVyAsC9C7SAH
4IOwhcqUmDxLyT70+j3WDslwt+Hc0qvstVA7w+DbsMQpwS50Fhz7+shJGYYeM6QxgK2qW9G6KER4
EO07ULA9Rey8m+N1XgIESD6jhdEREL599NyyefzNTfk0LhiI8Nhv7pxk1XwUfzuGrNZpv77TRwbY
xJ4UW+OB1sjJOnQjqkjm30LHqfLddgOSWAx5q5ov3GwVzYwvttt6U+dxx8KyV+ePAOcD4SP/05zB
igGAb50Ws6glKsyimh/nqK+58mz4E5s6QCcHYoMf/EAZ24Z/WYPX9AWzrSv3i8j1nhXRy2j6zMAh
h6dVGUXfXSw7sgEKI97UuN+lwzQqq/+WIo6RkyHgfSYwMsbQTEYFI2eYtlhOC/PluuQLCrcOCT8k
OyYxe/dvK8iz1y/6XqNfqtHnhl9xqY3Aii9R7bFkE0QJGOF3tQKnz9ZV+La3eyLkMElAOWp/Ihte
vCv6KDUDWXIyB5CED6FQ/tsGTEAikSOsrGIUjRbeNTigVPnCuKlkg//zC56iKxglJUZ5FoRvmLBl
EMerde8w5uHlIL09glfR6lZaGEcDYG901mbcmaJAdHdKyrYvU+VkQ3ZssBkctsouF0TVYD8h1edB
qYJMi41kO0VhRvry+eb58DIkcCTfTk4GWfwWAuWhPHwh6nz+stHzy6vTa+KZ5SNNTgzia3TnU5q0
FxC++edTo0w2w+f6Cz0qE0IZ7h6Fw0BrslGAM1XsI6uceZ4fbEGNIWnqcccbS2RBfhyCbDVzb3Is
vkvF3vSo9LFoODfoufOR2t1hBApafMXfTLD8MK3BsnXhVepTj5+HH4f3fH+ujhXgAbhFhksUQig4
yAjt8qB3IQ5ZoWYIboJzu+bUSNPfcqQTuETDOf01SOqNcQx7tapjL9SG3Zzh4CFUq5TPeKiZZugp
vXRVtdbEKTXwIWGZWcBMLK4+KpgQ96oXrIeQ3NfIS2y7haDvDSL7cSAMcYFKyBJC8RB2JVp6DquT
2IYrCTi3rqOSPTtTRtPgAA3rMPJq7INjkGjTyUcQxS8YA8p2DkqwRK1dzZOrkmp7Wn7jArVcx0ir
QWkKKtXQa1BsW3zxWw0Ao7D+8K+q2uAOfKzvILLwyIyFZ0iEKNBYXfknpuG7/whVM04Pdm6oHyb6
84G1mi5FinDWW5/AtCS7fgkdATuk4On2SgaY361OAGMmntZzXBbptWNc6c+o/j7oZxDU3gfw8hxd
a1z2eoSUJC0p5yL28M8DuRkoAWEl0Y4uxKhdYAbC9lSdaO5h5TqTdbUvOslIxL3vI19uDDPJl/ll
XQo37Z/a48xxAxi0+Ibv9r9ZJfkdTfaLSHErgOxglTqXVb+qGcI2glL+Hlj2S/CS5+LczATCgxTK
XeR1Ssd/HfyGuBPRW8NTN2qVoNs7VmQoOaqCTLKkQGKNCsVZsBpHQdaEbi3SxC7JnejJ6NNpKOwz
wCRTyGElTPGZ3h/vBMksnXackT04n3T9GKUA/O7HmRhB/zbxe53HI4ZnIUdgWgb8oJz+24Z5SSBS
9EY9DIeploaetn7QMGrClbqDPpQl1qtRXHKJafxBKnpR+Rp48+Q1JwEU6hL7Vhh4MOX7lkTVDafA
vVOX+AF2G7TNM5NX6keLH24EDKG+AMbdrvdXN7ItjcdefBqC0R2k+DoxkgUpcghh5FSb1AIy3zFA
qs3d95GSNVaWaZeqtv8fvCxDEHB+XHGRZaPf2LTCYl4BfCghRT0MdgyK9IX+mOvsXWQTqdLKEmk6
TlqL3pmHuwevGECHa8Eb1mvJWAnxKIidVxKwnbttY+H0SLtu466zzBY1qdtTVrg5dupJJZgGrxx7
RN9FX0wNZY0LZysN9sztDjaM3bHioWUHyJ4wd3V44pTH7xMyF1BoL396csfl+HLu9ahLUBV+dueJ
dfmqmSv3phdDco2r1hNBNNsS392i5D3yCFqB4Sij8fLNXFB1N/NZqlxvFCTPxjAb4DNm6f5md7X7
2dUQuEcQqSvnGaQCPVeKwmTFmIG3nSmg3mPjJXK7TiRnW+2GpxjfwcqsrmGoApKWtGAQBe/HcJkO
Lmp8L20zIMUyAwnuxAAng2sjzECtPOueve6mHcYwrslL2WmRZUVMsOk/MPfdtOaxIkTqT0fHHqTL
BeWLGhlAEDsLdsdGTxcN//4whCwBJzkVEJql+y0McF/Tf1ib+SsbhqARSmiuDK5zCO45ZIU28y8r
/u8O64c79OLZTDjeI1iY3T6h8TBCEq91hf9mj8XBnFgR8Mt8fl+Rml22LpJ1Xp/AJ4R8+DAx3GcC
j5Ev8t7AoYgHW61JiPL/2YCXaCcsZd8HXvPquVpsB5Jhfj0Rly+jKBBU2oLpr9ItGlCrsnrY6uDG
5R6nAwjTNj6czGHFGsC+brObXBoe6owxvhjESLxSeWbHpfSg2vB6kNH1CJh8tsZQLusqUVOj0PIy
dbD02ypi+oPgJ57QfTMjbNseaTLu10NgGwsLymMOfE4qEygDA8Kx5JunER9M+LdtHAK2yTXbmap8
b5ZISRDIbKXHOVhXcbezFFDhF4k4bW15gc3VxXV7CX8rYaVPOFAdqQ9nv2Ozbq527fMm4PYyykgn
KdmhjEfbLLkzt+XmVTmDsY013Frudc8u+cBq8pcHaz9l4wVSS7G1bEL0uRBBEv+esL15cI7K6MFS
alLrTe8Ra6vR/29bbYRitak9FXa3m5oZpwJwxKgYnDJBupfVuWw/7jFDXqQN3MTNgD9s1z+Zm5cy
F0Y/lslZIg3/CmUMVZvSCFSCXYt1qxTKPVHml6Tpll3NW4YZ4c09J5uGPp3GcMoNFg9cjoHi9eDN
O6F969J34bnNFK3s/G6rKgjhs9XOx7GZ2fIfsRLO+oDEQNMBvo8cV7oJQKe1ZOEGLACx7O2SUCtY
00JTAicptqWz1ZbmPlh7kkWjGACmQmBoG4JZEJyzw3MvA9vtg2xjiQNnn4ZG60jws46Qo02PV4VH
u8E3Br/mojQeOzYlqkniY3whvDVMjycLp2nhfgJPLikZYETX85chVj689xCovuC1ZTFCSrkwXbl4
5WCeggn66nTQtR8+ENzkc+h8yPV07bKJMNcdgpTQh9ZBKffXrSA6ocrtO/dyPRGD5rpAEqulDhCB
dFx2uZc2rbK2aMera81XnAOrS4ZKZGxjAPjvm5aMBfSgo/a0B+v4qPf2UEIyzFRQtBJ14cReNBLM
k8rcergIYLZKunr6814Mg/JFBpXrE5tXCb+u7zmnAS76LyiLWd5TNjmupBdyXXrImBigjUGekv/q
xi88yO6BIucpUggZZi4HnJnBOKZz8QaKOIt5MoHlFwG6TNs2JMUz89ztUxy1YQr5zxVyjLefx0B3
/WnG78OpB6SX8go/xNsfLkE3fVPhd21N6GgaHuxBKsK9ePXlE9wdBdE3v4ttnKcEkdjAYoKVR402
F4Jq8TTZNol5Vv16mj/Tq6KJIHPbAUKMYu8aHTazFh5CJ3IoDS5JqYnd7iA9GHbdfnghaYvk8TrM
fG3bg6/BQSshK70bmKQ5nGW3KWTxN6rAF4LkSuQje7hYdXtVnwkekw7i6dxEQb2/xsaep8Xmx/0h
CMR0qQBHUDRDce4lqEIyR7uL4ZgH2bAJTYX1BjpKinHAAaKIlm+7Ru4weKnUcayvPKS/opt/ZMA5
bUZ82qsvbFxAL2DL3YcoZIAGhfSPhuGBpaFgtsaDRwRxpdFrEP6Wl95rX/e0RN+ZLg2pSzjwwyqg
v4WPYT1DTOexthb/41oO4YQnHwWGufwO0kdfeib6IvDTdohzGbHW9K3RxiRpwg1BLmoLVzuKSYgl
28G6tB5xuTFNd3qpJIfoWHLVqinG/d3KcEYtnFij4yY5YVsX9TRdWcl4WxL9XpmZ0g3/JRFA5+fg
3kUMOE6+5/SZ/IzN4FMrVeKQUBVxwtdfUi4e2X2W3i7lc4rl9k3riZKKBGQ+Tb3jbjkkM58Pu8BL
tINKYKXJgbp71qqso1IC3EnRMoZEH6VO6bY/LD+JVlv3LwWwOrAg1ALQf4iU+DYqLtm/4esrI3J2
vxaEmmtVLIq3rLEOlsvvCwkommpttZqwEuOZHr5JsZTb9QSUStrwUPo2fFDSHeO6UHEmSmMA2RAL
VgJbRoRZAI5YMxv1eDHrJwYLlJ0qk3/YTRgSPjlvrplqjCD8qRNLbods16azHx3AS4Fa+rxBS1GM
5iLEmiE4wsRPU9LpURLOcxuLUZbMbfeYLlCjsK2deKxjllVN36cnvfut0GnTg/WRQyZLWh5X4t8o
DQn8jAGrdUh3AR6G++g8jA74+NTH2uTEN3qbwYKmTrbbzpDcoClycGM/NOKQSqYFteqXBTBM8R15
W+NzeyjdAopcN3RJViF5pztMF0/nI7etSWxH9wXA1M5ZcMQInCLSG/t8U9KrkA2nKah0zp+sNsuh
Es935hm0C2ZIpkB6gkT+HWvuRF68QdzQiTchXVY5p4NGgq4ZPQa8uKNhjtYPgjGGvD2SRk4pivnb
YbFTlOU6D0VDwGzVPGofjx+GmsxXY6xtMNlIg4FgmbQLG36osB2j62KPOWOO0Dbmh2nTXhEPd8c6
NqHR1MkKE4k2EtBxMw/ERcrSeBqfg+KHwNxgTpW/1syZCvPN6z6yMU8vGal8Ibt1KswMT2QLpPH/
X0MO+3dFf2g92Tc+h9gtUhHQ0E5i1SMRzaIrsOquRlqLmbJ/ZTxeVbJOQRA+XF1KiQO5VUH+wFhV
Ok3iAM2+1m/DV8dySK+Bv+Naezm1QUW2PTaOxALsS2rJvcRdWGPMYvDp3fHWJn6L6WZbpgTqZ1ru
iDLXvzk0TLVzCOy+748XZ8QIwa188sDquRPp82U6qxJfmmaj4ELw9E3PYo8l9R+LIpHp+HCAUL4P
34gpkQdCJxINcOgsoyepIgiuP58pjx/SLkZYDPQgwox2ViqW6mg3dEy4sYpp3bbOAljXLI+GnLsN
/SbwQ9eT53XtE7woC3LWeOtXdTkrGV9Ad0j5zN08ppWszDgIOLpjGiLdqWjIvJG6UUQml/xVMw+S
2MlQCCF+e7nS0f1vtu4ejKHBLgTAwOt2zsgvfLKUVplolHAm2TctHyhXQDvw0h6VhL9+Bw5uyxtV
DFeD4J8WWMNhCh42X98aRtwwchtGzFE9RX9R/TUoUQbeW7EorAyNHj2fSPnYMXa5w1bCL8ja8qo2
3Z0T5H+JYxL7H35gv532ebGTkAQWZJeiOpoPhJo9ra0Xii+Am+D2AcIDh4qKHtY0bbpy3YOGuvaw
HPt5+HZCkvR6u6vaMqHGfbUQ6voQ8hpEqTW1S4xSZ8u5dnc129Tz3GJr+NgYOxkcACdaCMIGBh+X
eMQtzX5D7kaYePofaziBfrYP5TXfC0zgmiW+h3ZMMS1HaY74136U7m+5Byplwe/0eEzJUicXmQAQ
OA4HhzI2m0ivFcEPd7F3kjqrIljGwAA0SLnErUAkBmgNz4G1AaTyVHxdeCIjKOZIB6UeCpe7Y8u3
bNVhVgH4sOGPp+y1B0sAzyaMczUxFaSblxaYJwQwYTPQWmkyo8iu5eNvRWP6Ibf9NqSFW4pXjH19
pvKUl+DpJtT3KxdYuqxPzDfGzMhmOR7Zuc0fQUCgUHTRJs27MhQRHWXJ/8wuxhrQbyV/DkMkDbsb
6mFLGwGwwud0OP/6sj1nDALOwjU9Htyz+LwHGUa9s0Iqvrjnv7sMSOWfkykmfNrfdRVpvmk2Uque
Cyq98QrrPJxoY7+sP20W9zNN3abJTAHMzcpCwpRnqgmgnPZ5JetUDnzTnrx4Ii70jZuTfJfsglwI
X18u1ynjoqqg812n2w2ScmnSPFJgAek2XRgGVotAbBfVScMiwR12AwmvvLZzo0ijtmF2/qJ7TUck
94bBQgg36+VQPUaZRuM00ImGcE84KBIXPZXPGh9rlD8Zbv/ruQsrieOxfHyYiMSTtn8f+lANd35D
zNgTJLb6cdWn6ykbBm4sVdwjwPEJ0V7NHjqHGpAzgZLWcuENg6zQoguN4ZpOydmFWONNM/Ih+caq
b13OtBnfx8YITJC+I6nByx7Na39FXvt+eIviDT9fygcoqKihH91gcBHrEXvHeqH61MHA3Tp1LLh7
xEeCgIvQNij6MPlNN+OJvdYy/xiDm/lUIx7YTJVeRFxC+lV2Es5h8F9sQAN9yeXd547UC0VDhK9K
Q755cNo3rnc+YZ5D4a8eWIE3NZfA/wWbCkZClxcVcQ5sPxi7yWvxhg4nItLfxzrtTA449YxPdkbK
fTMuDojh89TcfB6qP/Zem2ibSpiSYzps8iu4PXTpjAIEbp4D0bY67bt5YRwS3kMtorEKI7tK6o5s
nXZI8Loi4ZWI+kcDk1amTuiQgDIpBY0UwfPxhKw3DhfKTeXtvi+8beoZHDM34VJ8iIIh4gQ3/Did
SmUaowsEkXBrAArOUbu2ZugOVPwKS+4OxyN7B8z9m8ikgmWuuUt3MfY9pnilfHzajiYfvsqrnkHD
I8ec/9dZH72s0Xw7MUUL41miRBysmKT6by/7GvkJv++RYH6mkIn4gHvQrsoFfks3kengoXJUNuhW
jO7fmjqOnUeefLGijpGS9I+9rcOQCLSjDIFGobqemMLJsYaWZX6avBHnsag998DZ1UGE+NmFR5WA
yDRtSHVUM+Hn6tcPltfba1bG4spw3F5SPmfop10IKtaP46W048FGbnuFIigVf18cfRIGqZ2i87RP
3RD4tz0ITITO6dHUgOGHBofhHwpMI0bXuzmthWkGY1L1/2/Aq3USLLsinvWw7kk+lv0HlsI+MArQ
TQB6GfVZcGxzk7KlZI/njH0f3oHa6YI7fU/BkjOH3tXMbqIXphM8MZxcbCPd3c+37/RZGccLFUnJ
DueY8uLeXLJ2feOhaCpXf2RYhFIvoEawj1n33BlhaodEkGFYbZywOgqll/mGnp7HU0z+oSsCbojx
MAnomTHfen/pfG1cQTFdKXsWtYN44gugAl3xLTp1bstwYN4/2JV3lFj5eur75EM40X9RLNXqeFsF
tErp2vd3x9eIxiKIxYzVMERdBhytzySEXEWrKGswhKN8X4LrU82t2eLUXvELG1say4kaB6/qpPHe
qCUVUCkGv72gf6RKYc1pnMQqt58Aw1otu56jZ5iPXLcDR7wbw9UJSqeueh9BTVDi3sHwhS8hNYeS
wif4eixdtS8gm1kAKkRs82CVujMOuzMUzJX48oJ31WbNZ9ZW4l+B1vKVm5CwwK8KXBzAng1hGuR+
O/IlE4VTYybwMWCO0Z6TCavfoD8DI90IHlJF5toNlCy0vFyiKhU77jWe39LDL4JicPTM+stYe6Ps
kXPZOf8Cn2nSUbRxf2P0p69s1QeBOlmmRUP/aeE4iyOOCIePf2axZgB9NM1WwheRGB4+eO/m6Qps
pjSrmbirR1dmTwtz5OdnztwzT7Fmgof24rRdEzym28v9+7mG4BGF9427d33wZBJu1qF9HCJvMo4I
SdrXm51tA20DnyfaL1q5UTmP4PB4QvcSxyh8IvFhmTQ80tlzw3xoaiOFlaNCHLqvmotMMlNzEsBf
wn8+uwsO+Ih2ZhnzV9kJ0l+8JHQ+O9c7g1xGRdZ9VJOd4Ksx6zQPqQN82xW5m/6xKg3o5FekoUg9
A0WUMCjWNAeGD7WW30YBwNl1f/2s3oZBlfblFXXs7z337ms7KNO46HeHYbRJZSzyJ4WbL/huYdPP
Y4hWcTTD8ekOTjgXPoH6A4qOwLKTt3ycL/xgzvsh5vdnHvAfXFPDxnq6bbXbibGidZwuIXBeem5O
Iw38bgRleAZdhLS89HUv4UFKKDqURw8drxH1mnWmQzacIDowmaKqNteMDg/YV64WS2pGobWVJAbM
DmBatjNiKtHEmAU5NKNuR15u8iG8x9JRI7JTRfu08KOKNmIIstV93JmcFj/sGiccLSt6kNW0AvQz
E/KOAqSSvD/OuSCjEonY3A605L7H5Aakt1VV6vuVS+hO42erV/wVGbq1mhzY7UL+h6vHWOHd7j4m
hPBaDO5H/mvy7FQnylwwGWJZKQ3e9v9/jzUCR3R/PIQ6LgsyiDQIADTpGtDfr/Ms6VW2JSJOvw/X
mNBCcWnijx2YAXWYyfqu/I34NMjZ6QasTJhYl4q4vtaSkY0ZggmeKAmq5jkhFxGNYL2sNQLs9BWA
4mL7w7v78nXCtM2BGlWu7wc0PLIR70bAJb7vEi1w9FF7Z+863qHUotb1YjAwDx6UTojoLol7g3C0
RbE2XBqJa8HI2Q6/aQmIJD8dfmswHhnpbHqFLyDqaq3UYUg5i2oLnZBkhjk085xnGceS6yT5xHbY
LT1PL2GP8N3/Yiauv9TkNH/tJ9SKDNj+qLCF2YOyEgCSKn89TMJcqoiO/FDvvlivoO5KDBlhSknV
VsSFd2ofjTvSwZ+IE1cJco9H/vDxTYJk5IopOoaRJN2JAMagbJV8QgXsA+DcLQ3EcjyeOH0d2DDh
iZplxFp78gVUBwNbz+JzgBgws1rXT3FsJyHrWvqngY1MZSJGQrlRg/F9xMca/sJoyOoQopGCvUNn
DZvvswm4+kmlssfOr40lskCygAh1q1Tz3Cj3wj8bcdvXVKxC5gMmLSVEUBYsMyCkgLhVsON6NP6C
gFzH2PiBYzeNidpjBI1CJMFirk29QXf/RhnsjxpiOm76fFa61VuAUFj4XxNa3wcsTWteq56jxHO+
EuZlbZy9Ol76apvM84z7LDsVERxAjHTLnkZBL6eaf0cADmxSTRfNEliOgM5gaLGGYyct6DU+cxEg
J/vymkc8F6VWsI8e+I7/uHIKrF94y+/shoYy427GRyTArhcp5gC+5yUHCg7WcYKFGQO1oEhjK6bx
kknQtNaUvFw76pyKG7JhvvP3kbqtZxvlDAGlNKCn2gcnYs+dCc3QnDeVUCwylpDmXpKSzRBJCYJU
xefDxQe1Y1dcGiXuEn/pHG+x5yiH2RtG2dnanuz0RT+OxeDuJA9/OxC2DeQkX2790ppsF6W1PfiW
Cut1sX8HDlbR1XCgpuhqIClIuJ7rxD05yEpx2TFtw0nT2wgNLJD10mOP16d2TMEODzWSZIwF7Sxk
KXC1K4uJ5tqo8PHQltHqWmrEk2eFboe9+Bt1Sg3G1R5l1ltteW9ABlRmdxbi8b8UAa+mouHb8jMT
pXo3ldyiMl0df5Mr+anUHWAfGJqAq2x0uAN+IFtd/OJacA5By1fvPeIhiEQlBXZsjrihtpKTsciF
ThFT+KBTc37LaO5faqf1ppeQg61Nlan3N0+FOLMBcWhJOknV72x3L0HbStH52WGEuqsUEFRCb/yv
hK09za5GGP57QPXKJjv/PeXo4V8Z0S9jR3OwIxnKSp0wDKMMQk0I2vgTr0+NY4Qehz9Tg7T846Fx
4E+oROYYo9LpeW2e8bt0iRtvMulhAr8SH98BxzhABUQY8FMDhqyAQkEXJwnalazQmzd9jcIAVq3W
0sNqta74TuQACS6qG2fsOPFYoNY91NdLue+60bTrUhVREDqJOCWWNjD/OlkEceS01BEObo96as6s
UjPDcTrDBOEo+BjEI7DdZNVVexCxmJJinEUMDVHz3H2IjRZX0rB2MrO2Md7yu7hBkFPN57WQ1oua
S64Jt2DkPOZ4f10rKG4lTQgwbQCpGW5FUxNXmLtNwPv+E6zFAcmxSD8wNcG5GDNOFwmYiWGPXT3+
gvXqyrO3xUuxjgxuhJkhOJePsN3XeK+wnbRtmKTAbFiw7kr0IIEN3yzeQq9pFMmb0q2O6lCaRLbs
kZdsAmBuEyDs8/dDINGiOIo0d7TOucRnYJlc+wI74cIJkxDnZ/BzIHQeteBzbwjxQ4uf9HayUeY2
SRKl41Nhb6XOfwb8I1rD/XpdMCrHwL43axcFeROio2Sfq0536Ny91W9L5Moy4qh0IqqZv6k08Cyv
PsUymQXfG4K/fABypEZAV6N8bO6oTYE0+ee8mRH+syr6/BpsxFojqjEYWvVatMTgXy0rsFgFX6dv
mWuO2S+zEHZ1EkXnScUcHRodka2vdmK5XjKZkXh7TBaNS13PULBwqi4UuMijZuSFXapssfS75epO
r/5GPFn8TL4WlOpr14mwm3aRbBrUnWwTLBrk3eVCZp6H0k5bIBLUM63z9f//X0ffRoRLTyg8yYcG
OOgnuV4njZcXKIgTcecEw7FnQW5mBzmeISf9Mj9mUTk73DGRgv0E0lX+Zu+RQNA2Q3PPTmurtr8o
iZ1vbZ0+6BJDAOG2/wsWsQp8xRl8sIUWW4TTZXcqhBVGVJK/6ud6AXhY02+cXAIqVmOLFt6u4Xed
rcT/l+7nayCzprrdI0zO0sls0cLz/OPWCCha6dwikOFh2bphTfex4g3z4X1ogcs8tWx7SMu6gAIM
VMo66xGAtm/n/HRrTD70wzMRC4yEIUCCvuY8eAHD0rjanrehTaDCkpPK85Cym2tMulo+cj7WtMTQ
Ws+LnkrIG1R1dI8GdwZZofCDpeuPe4rNnVZ4GX+G9h7qBHwiKCfUpnkTUH99YLqmNt76f6ZEEVSr
8Xz31mioIqndywbKySx0LuGVTmC92lHzt3p+NENHYPdIHystMyYxcC3bG14+L4OClWgsDAYKQxLt
Uc/rTYNIyHGPi76njfUhk+4sMiHYqZesrbB2pQRynxCAomdbbeMAwMltaP9TJVf1eY9kfVw3mpSX
sGMHTMs7bxDPkUnjJ+CtR6vkQg+NkR0M/FFmSNXGH3MnMFMWsCFqInpOtbaNnu3nAkeKNzjHBC3X
pdzP+qU0AxBSq4J55RqEGkEan5+zv0olXovE2L5yGFe10ef3lNZZIpeBFG8T8eDc6V4xTq+jTMyD
uNRKoGoVRsR25NA0KkazTzS3ttLlFzqhrIOivFdXEgcasY2Uqv68UbrmWzvQyTq0Vd3t5tnuUU43
efXf61Zka4m/0AXHXbe6QEgiU4rL02qCZR8xmEwvl7XdYiOvCMrJoE4Nb/Wq3Xhn0ZvSHaOqmts2
jbxmDmdlp/e3+p0X9/Km3f9DdBYJrhRViTKY93HOoaFmn9Rea4WQOciRce0wxSMU2kKI5eI9xl/1
/LT9193bLmbJj4z/draectC7MXtXW2Zc2GASol5kqx2h7IDPqDOzb7NmkBYisO4hGy3prgSWZE9L
0zbP8uAYPKp5jIQkkiW/lN07LHJGTNQ5AywDyv17AMJizAcAolnGFjwbvr/0+r3YH0qRTQ6o1Bio
t8rt09m2C0paPj7MnSd/FRvMiWJ6B5rF29XWzO/YVb7FFUnJj/BCXdDH4/kexTBVhkf4NCT35XKT
1Hw0r7AA6JAtz36d/EwH10dd6La8U6rftsJTWdznQBzxStpse+hO77d3aFxJj+IpnGfRfZScNV0d
a+TKSMO/6Q2FM04FYJzF/oBdSthlfucyYWdmj9PN6aYQ2mesyxGPCucTIVpB6uftTpoVOvYbn5qo
2UdK+R7tEPzjjSzKQ6sQs+XxnxJ5X35wO+ixV0ZvbI36l+XN0j5Yix6srjWcEZHuhtT32oQ36miz
jXztXiniCbjU4Y078zTyS8bVdqzDmQ/MmA2eCrNAUTFgDZ9RDpyT9OYp0HimG1JostN4xd9XJAKr
dKso/DgJA3hlyVEWzkSyStmeR/XXkC7qYLRkWZU0NIJ48wnk5UL/R1+3/uifK+GaAOZJ443OWk15
ae9rwMAy26+PSDjd7RFZF2rmKJaroLMI9YQiTnaovn7eSL8RVIuLGUAY2MlSCoZXdDuGuUPMZeVz
yAFbv7Stg69e9vb1Obkeyple/e+bfyHw93NM6/hVcsqpxj3WLHIAzqs2PlHgKQMeMFcb/CU15y04
ljKaRJihHYEHUSGXGwEvDx88T0cqZ3JWamlDzdoPehGfKPJB4/nLxp9rlgbSZfTbXhjweWEvKLEU
LVofEW+RsWJPApgmJj7RNMI1kCLBNzWfApwNU6jk3h8bSp/vTg9GxknC0kBJxWEweoLjUYf9/kHP
tsh3KaN/oxKbCYj55RvNIp1AA0cwT0DWKmvkv7B5NVe4++fVsG4hwG9Te5+XC5YByycKWxap8hnO
9gU3xbYWVhVGnmK1M8aNcskwzBnYQomW3St8wAfcaDBmGh8pZBtqvK383mOSNe4GLhmwMSrAy58d
vFxeblnlAH3mEGjDxv4Vh6t/ClAZxEeTD9yhJSxFTQ1F9sMtjOkWGF89rC3qwKCjCxPzeMKk+MGj
TC6bb1XUN7Oj/c2S1UrND/I/LXFMr5MCZjtWTjUGP693Dzcbt7RIJxaGcGAa6fx5Hu7nD7ae76UH
6fKiElYcef42F3DneRc34NBnO4GxeVPkIo+LuImomPaPFfQUR7sJzlAlyPCHY45v6xp1tBU0uflG
pGIAy9oPJxTVmeIV2DF0yXGDaZIIWYJnkKefGsycx0Llvl5w7i5WleiKW6q1E9KqUmWZxk6+mre8
IoAnawHUx+fx12hp32qcFdWFFCscpnF2wpmHzEBldttJf1x2D6xjnIsiFZEGjBoimsA7To81vpmc
EDyeBLSqHx5SMT7C2NmWgYAEdEf3XCnj4yXda3KZpEAtazz6U+OlQT1bf/fdfe3pS0Egj34VDc3k
YQnF18cwlINBSadttEBmp3fdFeO6Gh3FE2V20MYBzXSYfo4U6bjHABjNvb8EM4U2uobzrSqpPeie
UP2u1WmSAOcVScEqLTa06nZiOIpVBaShTMNlPhnc7uz/7Vo3tFxlMlTkme9LPmIqgQdgcHGYHIbZ
5O+4YAcEMJJ24AIi1ARUNPpkmF1xQYDUdmMOKdJblVAeh8+nMQ4pwlCNDwcIc1ynglscRn02lcxK
23I7sLRlrwxBFiJVj9ovye/DEY+YmttJZrbqQwyGXMRKhfpkOPOb5NDbD/YiFEeCnFoxpuq7gb6x
kVJmLGl3Oi1uUE4AEUcE+2PNdDB66Jatr8/aDn9Qjs8y3cH5ynDTbHGbxfC2SDqdHfK5RoJZ2yNU
yDlxZp6rtRurbEhyiFtDFzOx74L6LZajUPm6fq1St1ELRfrhuL3Vmbd2119BHpt0sJJq++nKtCjI
IKkupW4I8WvTHauga/gykWE1CeGzeEzyc72/98/yGsDMS3b6S5HMMPDNuPgsOtYQYGiF6WpJFIDw
MGDFsEz3QvDtH3mxjDqpBed5D3PFN9//fL44t0km/jXcpNdJd5tCNdryU2i2TpysMJJoryRT9vVy
Jxo2zkQoo45WszfcwaMAhvvqJS/gGjN4PJTH/lqE92KLGwDs1WuPjMKCOR6dT923ON1cMhELfWN7
cWIieIMsdopT6DNkKv4XfhXBcHIVAn174qHVEQBDBWYy4kLRneKuDqBSvkhGJJMeAkW1F9I4Lol+
PXzf0wpHzg+kppOo+fAPrwkdQSGN+QxZyisesW68VRmg67XWNteo1VD0TrDX7n0/YRFYnQfHHweo
Ri2oSM/53/DJy/o3/z7rN5mNDjdc63sI8wijiOodsMFNSX1NPMaa41I8fBEM9aAIMMxQ3kZMOD5y
WE6c8S5W2Jo9XOt4GCB0H/+TbmG2sp/TEcubDkL2yZyzTrkbhXGjzaWafPXtaSA93l+wz9kI/Pt2
gQR/vsHncsw6CKG7e3THaCNByBa1wuy7CnplVC77hpKKMMeIvnNYOzYJYzEiw+UygCFXt3512757
nNt+xFEKqM+6rnZ9sfU19HHUXng02+lvT8GbWanCC/xP0He6sNSFMMK/KU6dN/ewEuagzhiQ/+KP
WE2eDWCvNnm9S+BUbukg2WqkozoIEevPD5LYQvrrtISrO1LTsWEYNvJflPmyyZ8Y7oC1IZfE6eRL
p66xeZFPyvAmMpcMeblORi07xNKvusuxulePfSbx2IvgLpK/PngvblV0QNTn81Kt1r4Nw2ky+rJv
uBgQUK5B4WimcpHOV7cGJ1VD+olup2Nu1xyWBYeL3204gis4wWHe7+E5XHoJFkU3f4q0WPMQusDS
nVgbhyfNeKAkTfFBmgLEX8ln19Jfg+APE8bJHwrzZ3peZAeLjbs3WAJioYeVZA/lQGOEz9saew45
kN/PFh1pnQMoTzS5tVUwtWwDuFIrC+UoPJqYx3ftAOerpKlCRh6EHp/WJWcDwxr9BSFlhl00aQQp
NlEnv18cYHXvRdla6LYzXlIhPpOZ0A1UFDQ6AYBZX60QxbUUx5XU3RzooKRg909LsGunPGMxeMDl
nQovbKI1SXnwBPEIbodNGXjWIpLO67m4osTHZjaM3XKqU4MlmqJTNKWb9Ey1+EX9tkLNCnAYxy/C
0UzGGg04RN98lUtFsM9GAfAekgmoXLD/ND+Nj1PkS3JFU/lbnTJ4GLS5N419CuPSNacBD6yrZIWC
NHCmHXaNPnTdHfjPIgiXTZwPoB6sw+q0qZID8cGUfF6+XW4pOBgh75U3jx1fV/Woyoa6mZO6WHhq
fTl92yPl+v9fDYhPlcj6dvGAT4yNQtpDSDKU4Y4D3xPzhXglleep3YAtGLK4M4b39qG+g+tpdfnx
qNVhfR0axxkN29SEoiYszXIIyQA1b8edZTuk6DEqV2XmXmbEiNwC7mIvXLQNEiYL6BPikyget4nS
CAQRUkb7qW0NHEFuTB4X+kqGA8125z9py3GCXTsO9eD2GY1T6bdIqowbxRBoEgVCNh9+YJk40lYc
9xyZnZWliNkfJlSewwYyuTFytWZDUqCvG2NlbLaVju+vnR8gxs2tYdS/4Scbmtv3ZPoFJq6ojQu3
iROsBAWWXN3t4bAtRJiRFZMvyiqjTtEywWZgwpUD6AZEWe1tE3464PLRuipmtq52zmHd1j91Mn7s
BZ8v4dVj440bRoSKvwfXxhHJSBkLuXwHKQxQwl6L6uQeKIkzauLbaYLP7s4KTFjU0g5W6PiS5XHl
i4qlsT/SH4XobtfcX8iSQJwGCahO5mvHBN2uwZoMPkisjgQBlF5qZkqBWakJU2jfah7Zmam/HK0H
VAAYsbns6HC/9DMcOoJxc5uvY2MlkOfu8HNeEQEjBOpOFpx7GQUzvTQPnA+Od1KAIhgPEgzh9GHO
71NdQUUkw0SGKqjI/t/W4NLHDjesj73+EGPVMFXR4elkcTSubu9cAGzD3izk25mCC6SoSPHkIAAa
6j3M3pz/DWad19CDWL92aJzaqLHSsYNBMUtV0P/2fFS1LTekVl3gY2ED72M2DjpUuXGp9i8SKGla
U42fkd9dBVIx8bClmTAzUfDXX73Mf4YQMZLFlquJ1unXmn3Pvgz3WGHEp8zZA9/doJqbvZt0+4ty
v5ZtU4X/aJIC35SRD/711kpXBTMcIpM0katCAbWX/RyPRRtAWk3oY796IJKBdS1KDHmSSqefJeZX
F0lVRlus44+dTwtvwxr3pB+0X2oyUjLWPd1qzMjm409yXsy9WfMAszHCMxU7e8o9N5LhzbuLYIKz
tY9BGldDVjbCHHUvYsf/1x90ItpnbMrPMLTYq5aesUroPdPbwWdDQVFJztf9gioTxXkidMfsq0w9
bVWL3iQJQYNkrcyVGERqlB5MlsfyD0ayqNmtoSNb1fAO1S9Y4mSK53f9X8jXATAT8E1xnsLt0/Op
QnLt6xh+0LqtrRD0uqf0ROzkLvHY8m0zVtJFr8O3+quGYQzilSjCgFp0JnVk9TBhWNrjxat2LVE1
S0gBAEMbYKAotrgDLqVHB1jsib5HkbH1Ucbipl30zL9283ADNzzJ9UA2nmpzXLQrGlZhjTDNxVFz
ct+fk22I+CTj3nN4hk1usg6eE7fDvdiN4kqA64G5d3FUdrAXzKEYqqEg4mb/t2LUU9bJJ6ZMbs7r
IHxJHig0EERqtGTvzwUZlC56Y3HA5mblZzdNOpVk6aukL+kU/fCJDfL5stPe9JY1zev6nzHHciNu
fmD89blnaOd9MvZKvG2d7Hv6WnlqhKzd6VgDBPQLCoAWOpxH+wFBGlc3r9itTC+l3LyJwoNhHNs6
3OTTtXFd6MUEeRtxbIOGNFZuTYwy5UOTjXDoKjztzdAM/x61YormREZIj+8lPtjIiiF7Nf+/oWU1
1KAPmzpr9zEbKWH98WMf3ujE/OB0WvNqammW48CVbSMAJoLIBldljxUPkJ+h1AVL86runDvURDK8
aDu1D3luRJtWm4lD5vZ9LMCY57PolT23mEFw3vXorK9Q242fVYlcqG1ZLz8arw6CRkRHfL3X/pI2
zq8vC2pb5raw7xDRlcjzhK0cNymFy6x3n1cE8OBlM2e5Y9zggnklwYcUaw2XWZINQNjE1bkPBf7b
cM68nVC/R4J48SVMZdoAaPT6gG9IucA439KXiHHp432yJ8KrfxwfTAIzzoH/hH3nvTiYAPAAMj68
y2Cu/EE1sPk65NFdM6LFZQV/uTYvU/B9lqo+MGDDq9K/ayCecAyER63oSr7s7oBUUUftVev5XiBc
hW1x2Z9O6fVtwbzWnR1MQlggOOF3GogDkENBpo+m8c4PICyCzSE2i99WqoT6o6B1EnnXN6mXPrfl
CqXcj+/25bbfGbVIp/cjt7j2t9Qt3Y4joo6XxE3bFatc6GXyVuDQShHw4sAIjY15MHZ2nSJkLCbw
4Vhm4V00GHZzKWwUiE7aRN/v1XsYr4KRtAsP88DtlUXCBL+1QrVRYxbs7VbijCnD8dOsjRjrQyoQ
XjNiUiwcOYiyTsXIbt6uZJZGuG7bVWx8T3reLhy4yTKZ2mk/Fw9bfYS8h/KmWr4ITVlOHv8SAQAY
Kd2ryzkHeXR3LxCs+gzyup2XyLv17R0EAGQcDdos9L7L0Qikag2666Fu6S9qYUpdRJBvfrtc9Ys4
PQ3bTQng8oHumNo0IFlqG3lPcGfpgYIh0DczJDynzEyqlX53vsTVnZFHhmrNx2VyC5FySHE3cmAd
1D+Hj/yIUFSgYALm2SbTulANQqhfuxNzko+EmylAQxdP00sDFeVOKoz25CCGaGxYxGbA70YSHlDk
XbPd9e71lHAVD0M6c6eUH9+g9fzdgcWm9fyxd5b6kXE6uA5R/lRcxlJ+5U6crJ7c/EiTIWkaNLS7
UmyJqikvY2fYAJ0A50GNcIns59qk0rSmxBaJPlgCRhqT+OG+HQSI2gtkhbg4sgkqgbm4Pl5JRo28
qD+j4rhRPjCFiBLTamtON6YSxLJtrktNP/Ra89SltqGf+uXEvyU+Ui4Qs6DIGq5HKrPRfMj6a5EG
jW04G52PwAhVan4d0GXi/+jgRPxJMV1HBG/iuXfkV/Igy8wLtfuWBX79ZQnOvxJaqnECCof4xuHQ
d8aIgrST2Iq3wMTRW+2IdtXTFuf+11PbOxMtCK5Erfvr+LDlrGmPPtlhRyQebwmw8pLWnnewW0eh
FjKI6CDmtp/Bx9Jt8KmHl9sNwbnc6BN09lvVhyBP5DH5e/wIF01vKsfcjTkWm68v68uzn3N8L5St
QeeNN/K9VAKBq6//ZQ4/0RhefoSHb5OryT/Xv5MxWdn2rYXioFK7pID1lfuulqXbouFyxkjg6CPM
XZtkeoF4anR2uktI9Bwr4tw0QI+FlPirEmxMNmeI9lLLPJer9SyXU2xmiIaf5W6JzLU4xjqYcnTD
B4DkyOB1r2hs7jo+2eer9s3ge7vk/iwlYXNJE+RtzcllDPOa3o5iiikvDFC+f6/wpnwMbRyuweUk
W48G3osYbrWL+ycrSl5dVrk97EI5PJ9POJpC8oGmlZ2JcE62XvyrDAPezfbBwn9BxdzMgCWJ99r1
EzjbIb5/bcGbTB/ez/vCondIkwg+ICSt00vL/EPFWSri10QVmxsYrRYuZyPrXzhDrgm5jpzokE1F
uWpNnZnLjsHvU74bQnyF2Eb6SIdrM/tHgT3LFWPYrFU2SVCh2kQE4aCttJjeLy0qnme9ltv9yD6c
YErjt4BTIZAnIG9OyvAugKTyI8VRvxxn/dotNNS3/0J7orbTTqbXLJ0UhcToeiNhm2ZKbrckB00D
DGbHgBXxGS3MhyuyOyCq49UpVYtLX/TYFaPkEE2LRO1P8h11lmmNR388k3uEOV2UyGDGk4+UX5DY
fNVlJ0315AlCpLSmIzUWaz5X8lIfBZNt01pz8AVzXD/6Aad4pNCgyWD0o4h8Z3xeGOpvm76Sgq2t
7aZJNYA/Glg45+m70aOnvSvfhU5ao5xqj6wJjQKmb58nLgZ8qw59cL0GHByHYX0BdRbJGkcvREXr
MpoWFin7Na3wznQ7Y3CwLb3Y9KddX/xUE/gNXOxQEYXqUsJU/MGKoCIBegeefAUOLw0yl76pOYwN
CpWn/Q1A4G//uvngtklRCJLTIGsm5sPUXS92RJw93yfh4XS+69uBNj1ajCY8goiYG47SXjJAad8r
ZChCHoTCyBqFIfj8AY3EXw5y1N80ywAAE4ixAze49tdl5FiFUtzuHeuXvbq9Vp2Tn9Inz/AT4epO
hAUJZ/aL2g2tNO/J6X5BXVlU5A0vQBqIbvHmKsR/l9DIoNzJ5eqQNhvDpnabKlZv/TbsyHRYaflr
m+mUMPe4KqL/xuzNkh4YhSfHTw8BjCx9HSFbVvWtUwSRBQ1dSSyfLLet+X6EjuO0/rEMuhh9DWgl
3rMW1WTuac355TcpfKVU1/eOIds6auRhn+/6nSej6OpDC5lRSJ7OmAPREILDt6KDzFiYMGdnqcjw
NmjdEqOYacV7F220ByDYW7SQ+bFeRF/dOIiR9YrQGkoZ/qLq/7i9M/GNAtemg3S9xdkJru3GhBWH
UGG/30rJ0oin7cQJNeKYrO3Tm0tbtUxcPSSNRaCgxJvNUK7lFvq/QOYPruhxZgfLphEOdTF4yKAa
45wXmC+xLVMPpnOyp3ObdjYgXlB6yPYEi2j8hMZ7tgVM4r/FW0E36VqZgNtWy8nQqZho3EwGkE5V
/KIXxW/Q54DQA28hUsOBIfIJHyLgHWvVvXRV5BClaqbcfLcZoUaaGXKWz4t2iA5iUfyCqnQ+dBLs
FE1pXdeUBAppqh/1c7n7p4wqv5Piz+naT8hARXWIPsnn2ecUsTwg2oiA5+B1IlQUUa79i0sOYSwI
a9KJpmHBsfHvlhIk1VoT+hXzmh0AjKuajN72br4yav9NTLkU6Jd4zzeLzvlerehik45+EH7kEwyh
Vqt/DLFd21SEm+VX4fYsz0gKmmxsMQOLoEv/4xEYPZ/8Bcl8/ET3IPBVp5HtsGpXwJRJR4Oj2JoZ
6FaZzwd6D4p9+H5DwX+ya+9f+DdeSETuVtCJtS4UrnqDVmSKKJjqqgmrVy2DQIRC7u0/BhsY9bvT
CrPMMAIOr448sOzmA1S2C6tU4WsLhIdynN/YBsDvXX2ecW8jNAw7pTdWJF14G0/Sq7ckorxGLPN+
DFQjlG4gU/cC5lx8SUQ4NGfwzVFc5SJkI93raFOm9JtXzeUN7PHal8sWkzdKwhfLG+Ma9sAVXtC/
DmORkYY8nV4XhVBJGIVyJajMjOM0jI+4DU9y7p5dZsOORNUj+FftVGF9hWEpnLPvwp4MPJ6c7LQ1
ssGX7J3wyTHQ5Sbm5rfSrBpQG9+omb1fapmvUtGIaBU6DD909xpecRC3LYwl0dP2rBfiFpxbBaSj
6fe5uI4zTqOZGurFwlA8Pxb2iGD7da3piyykD4TvYhYjBo1H/BWR3My2V1g32xM+YbnJ7MbrR1v2
oNUJHQ1EL0Qo3F1pcrerbHA0VRLXCNW+1WJiWvL+QG7JIs/HpOB8OfgTVi1GuO0Jc16+nJZyk+hm
SG2Xd+TgYE00n0cj75uCgYAk9gHawgUGyUbPfqe7MRXzuonyvvbwecy7BK6lOBoUfAg9MKFEmteu
TgL/ywivuiAstC9ac7snvfNB4fC2B0CFIYlcmRI7Yp828iJRTiy+BtQeu8bW0Ovtv64aUo1dUkHp
Fn/vd6vNBBofhDPoJbwyGRrEcY5ds/Q8rz0/FyKuybRMJgDM72Wt/fpct9TZE6R3oHGWTHcigr+8
0s9/oAqkYu0IabOh6GmrnoNhm2ZebmEm9vC1UwZz4mxcnOxFu4pKMi/DhCwu908Mo9SYNdBb71qV
/bk3KejhbjBTZm9qHobUStF7PKXn3Yof56Mf1Q+X/KfRxoNl3vE623J6r0Uj1+0NoZp0SFAmeH1I
KHmPdf+ffIwrgb5xDKOc/O1+KQlZ8hDlm/CG0yzhtbSYBStIo+8USKOnZUYhe6N87R9Tk2Ty3aMt
ROAkmmTZ3QzntR2wkfIsygL7pgrc+ZNs6vmtMj7baSveWluASf546uyWjlgI3TqEHxyN1KPXHshe
waEhHayGqh+wZB3VvkqJRyNABKvmaWeLtYBqBlXL+N8yatOu7pj60JJxYZK4iLp2WiganWPqJAj4
pT0hnUsbiVfJkkm+/zIQkE8savr1d1C6ZZoAafn5kE9aXmPpzvM9F/vNvyBjcY49kMvb2k5ura6M
VHkzk75/BMm+e89AmYOqVLY+JE17Xux3e3D1+PB6eTECHyIRqwjUYQO6dxkduq5YGIEs9Xf45C37
C4zthfTQDwmgTlwiwKqW+uBa6nPnCVyGhWrwsIGGYomeCZ8ixC031ZKrQfejJG6MO6OUD5Aw7u7S
QCndIKU0bUk3iiSGWLx0rBuMJhQp3wDD2mVrcNHinqEISc9Lf7a0eI1zne0JzE8HsZSnMU4/CsDH
7qJyBxAnmXDWzxeVoTWvqqUYIuV/aDKyCZHYg796/KcfyGnfNL33kZf553xNgYebxZwbb7k9P0MM
mFwdcK4kd6DYptG4vpy2VmYDHRLenKTc50GewXHHGCI/cjoQMvb98bpdMR2QAa/Bj8n09iS+D99M
rslCFaPxW4OLNDuJKn2J0e2bNatyBGTj8l6YAKg7QSFJqgpvk0pUj/KhRKpVvjTwxGCxD+PyRit5
5cJ/GzMWRiJwmtQRZi0zNZ3dAl/PEWRslItYhfcJz4XafzWIYqH0PdxCi9dtjfEEkW2M/ZlsE9R8
S2oMJgZNmjCjIZyxnliP1R2gUxJkEdp7uPlyqc7AirjGLlj8CHbq6NkrF/4bI4vDduIzELg+xJmE
fS4cSpBtJgrTcEaXJaigXjlsl97ayz1Y3/sMhQDtsS8Fx5B0Nn5Inn8kET4EIyYFjV0jC1DPIsO+
CVnsxHVO+3ejmCIaotvpjbrYGp2wbDtvL3oGVH1KroTfCXTejNqU9F7XxJ6qfSJWOiTgMOZMZMNy
1/DOyX4NqzY64nH0+dKH2KBcxfZ7seZZw1qHQ2819Gh4KK6nso2pLzXCYl3wcvrntLsTzrVDgE26
lHsIA2y1UegZF/J4tmL/XcuHZc9YaUJ3OJ0EJhMEJjPM69448N9+DrbX+Zjgl8K1wer2FnBi2vuL
wb5Ufkpbu7/20bCwREMZV5y+GLrB06AdYWctX5XpEw3L93kHk+lSI5OySLihczCwVwXnF0XjkKUU
PathglZdmEC7/2qtZViUQipE1DMr/z5bdiRfclUH+NY86yxQ0RYilJUpMGAlQcJuYkeKgiaXDxd/
Z+v+TDIHVeyzFg15igIP5UuIU2BYsGZb4262Oqf70cbxp6CXivZoM9oY5xa2GEtudgALZsZ0I4jo
27H1QxJDu/krLOsjr2rSVJ5Av2iC70E9FtzqXcwdJs2p+WPeLFkno9nrlE/K8vhXR7R2hZKcP9d2
w3mk0gsTKJO9Gp/jUmQX8VKZ+k4Rlz4dMPfsBGJr1If3LSPc0mtMrCkv4aBPjXf1xh8lbpjoWVE1
2VKumchIlWHk4iL33Kp5e3eONq/LWu5REvuAnkVjswRnW8WQQQWYl9oELyynIURCCDIrVShfTd3X
n1D5z5d95PlA1gv7YUsXlFxC6WK79mDi8p1LL8kOBE41+35uIy7f5GNTqX+Sx4U3HuJBwSNHV7In
277ra/DeJgIJtmv5N1/gJItmOYJ5whSHeleRVqrfBvpT/wOqRJATBgusHAu/a5NscW+uvZWda5Es
ZtYhX3JyGij7Qzq7wDPnxjRaCKBoNm+JX+UmDG4zIDJRfkmaGtCIbj8Be8Z6tVg3zxlwz3tktkMy
w7qFmwtn/MQGpXyEILuE1ztngOLM4ApOsoflHGGLOduO7Mrhzea9qIrQOAAroLHrNVDyEDvmz9On
rfZLweEZygxzVPZ6R0IiMp2spr0vCqlKDb288xQ5ILPhL1eRUFN8Gg3dpFWEjK9xtli7yOyeVh1H
Z8yExYJTjpu/ekKEKE0Q/OBJmuQM9O0jenasE687ycrJotHaIeUSPdceie9fZd7xhy/8t+uezugX
wOlkMCgdQOCdaM5ByfaKfzQs64q1RM5iCRXyJG5h8v00WXItB7dJt1dnSF30bZ4n5Z0RoBEJfUkH
RPyUxZ584mpXaZDUbvafbkR856qnyrFYRL89K5DCGRlCEhsGQUevyuxG97GDgkZZcsMxbj1vRpQS
cZGab3NoWXfsnEUb/ELLZMrR1qi/+U6p/DseJ18IhYid9vxzHuTYycpkfoc4F4NheTPN2WckFLNn
91wDW6Q5OT9IjzLGGx2UPIu1m+wGbeEeXRLZiv4HBaWi9/kBCYAOt566t/Lhya/aZKiCMXdnbOtB
KBcDZ03vgoJNmzjgnhsr62yTamGXWNzMO9qWDA9gPcBN3zgGwBZ1HtXs2mDldHfeqXwNfEstv/r9
BhC7qt179Jlz1ZSRqhj0rSkw3MCo4wzBbdIc8zzc2kCNBDYCE/opYM3GTb0wj0QUuZZKJGqoOlrR
8AKSqD2cgfc7H+Ccp3KoDwTrCQA8NMgL1L2zYnNGj4t1qAMlQWftOaKvO6IYa0ZXtrn8MCz6fqEY
Mfy6fHDEbL4mW6ZYZmTamHT3LCSghSIfOSIwVzyNl8atbMLIfsegwCJ8WobSlRRYlxtZ2R6WW4UU
Wmj8XNOR4f/+4gMklm7cnFfbJf7kWOCWUddbqjoiE9neWUBttwDZxotTrie5fKkw5lxBfIQtyghk
3bXIP3iFO39zyVGo8jl/uJwPVsKgVw+FqeYeNr7r4IgfkL4IqRpVi/g1GzU9pS1tTtPwrcEKMXdL
EIvsXPTldzuOOlFZjBHe456Y5qbgZOMdR+E+zMvpDFQJ/w7b2UIP/OiAiZsfXpNb8vpJycF8ecGk
lUZx06gADxP9kCZg6fYUPHvwshtMXLnfIqFSby0XGxAtsUjoUmS/6B5V0vOka8rTv4aevKl0cbET
s7dGCr71HQ3atWrFDYe82rtoSNHBCI3u+voACuYvCDDgyJRbtGRPe0dLOV8e9gfYWV7zJv787dbl
ocfRjY2tqHZYwsB/4rxAeGupAFWJczvUe8uHZMPKz1/EWDkikGCOOQKlLP3IFZZjXL72IvpbxORt
RWi9fOgW9mYYpcglGR7eAKE2fJgyPw7hbbqcaY4Heh2pON3jEL452ZzXgN0wzaHmQ3ilHYmdyzZ+
hs/uRYDaSzvAwmM6GO48I0iaW6jhfgdZYRKs9GvuAyuvMaYLehbuuclC25J4lPfUpb6Mfgu33Md0
KAyzWJlJ2db2Hl8OncdM1dirDlezi0EMOL0F9Wei7rZTGDEk4+55WSC+9Bjzuu3FqrHm94u5en4R
L04n/uZKb6tV7H02RBaHZf8DMu2y0qOMEplLfI/ROAS5TrRSG9MQ105gbp4UUJ02yI/x5sR/KhWA
GjG5i/dZHvCjnAAOJkN1CrxV0IV0Oc0CN2egO8w1HME2SK214t6aEfUZuix9+0o9udE9ckV5GisT
bbMRZ9XJJW27jeyLXijGiZnWoEDtWHXUGHvsuZa0MJxSbk9eUk9eTZP49onpVuWv4/q3yN9SV1SB
G/yjhf6XZsuigH2vXaD5quClkWHEV+be7GCMsghVAgS4b4crsLs0p2GF0J5mEBoLwCBoPxCWwZ+x
l0kyP0cgQvgktZnijQ6AOy7j8zJ3nWKX1UCSkjOfcPDFp1qTDm7+0M4wJLUGJrOukG5m3nw/rDv3
trrbmJ1l2KFmmKEFVO1tJJLMcjAnzk9uxK/INQrdQbjnFK8w8VdGV6O1tvDDlupkhUEgjfFR23+1
4po2gbqvAajMa36mEgSJn5isEzaFp64JflsZ2sJyz7PrcAcTSwu3vlfJtaDsw2AUJvW5Cy4NUBMS
XmRASQK5LAq8KhAH32/CtdbVnq6Laq9GyRbr/6a+nIV29EN90z7sarhLDtXVsgMGugYLTbYiidHn
f36txDGLlY6sRTUIleZVpmHPUQt4FhOr3g4mx/FlSnBhcTa7I+HL1+JbXJBLuj82X5kg9ohu+leB
MMh6ApDQMHzc7vbc0pVJkaPJp1IdvUdWYxKezECmRpB/RnrzzBpixBQBvoxlmEuq+2XhniqdxYM6
wfffBP9XVWgDxHwH+y4ZvHxxGG4SKYRyf3HUSOrl7xWfle8UaIvoQs1LjR3oYaT039ZuPAMEEMML
fK2w0Sbpi4O8bTRjlIjfWZJqwNk6XkiIcRiSZYrABZOz6Xr1RXNFs+YkEhDNTd2OM4UO2vFvrzpc
uh5Wn8bCpHMiEiixu7tJUdYdyCm9wxpb8FZkS6zuTHP8qoSTbBf0ZggyLVo7PcQV2XDzJt1YmecY
eA0ze5hdQUfeCERI4EgSYDClWQicg405TGSlLJVtMSQqFVjh5bQzfsPh6nY6UU3JBt96fyYhzYD2
a1dsvU25LrNd2YLzphV/TLq42Xn6SHQNmplYuFEeaO4UhjbJ5i5SZ9EiW7T7MZRCpQ1P25QnzZ9l
78n2uhk9GdUidVSa6sMcTjPJvwaSCf3O1CnXrY2dgeOaBYxpPS2TgcLGvLRFF6tC+LoCDZpHhCPA
mAR6ivJAwfHvLJK/PE7ERx9+t4EGfKGd+kzbjx6h3E6C0pk6wHbVEwTBiLz/Ahj+k1RDOU5AInOx
XjSpHU/lt4MCu4Xft72r7d8Ky9/SDlz2jrZBhyJ//dYMvoz0TPajWpv5A2BPvEt4X2JBc1Bb2Qzc
mL4n7XkOQtRJ9xXoR0fOYcE9B5v+Ci4szrpk4MT04QyVmHxc1WeU3W4I/R7XvQM8i3jzLAvoBLdL
IpSPZJfhcv1foj+IPj8EC00fhgPaTCyZTuClwk0GQn04K5kfMBtKCqVwEClTXXUpbNBTbCLooJle
1uSgyCiCEHJO//mb/r/acmAvqYg21k0u6CSzEmFaYv0IuXvFxMXlXRfisik+bG52UWJvgjuaVcrK
nGDlsxR86U22mmzHsYs4C29VVPynHbxMat8ZM+g7UyM+IAoLHVOcXN7Yrawo1j4Na4k8dDi+ntDX
HVHhm+Uf8Die/AFCLCp1JMAZbm/+UCkuW0MLyKrMLOWtvQ7KrN3YtSvLe5JpC80b8I2sVjecSS2w
MnDX336s/PBLAF5aSPMaIK1Z6qpJJEFnwRxmiuMMJtNG2BfQ9ZLD4FbRobcYQT/hbvwJ3v286VxT
Osnl2EPoC2Kx5+0DlIMuQ05HGplPJBWfzt7aYhDK2ZincXbzpf3Fk9IJnuoHxgwKuR1TKtUWVLvj
9i2IeTdopNQ7vIfWhMvcLrP63czdjbmtttBM8FXQYedHAnLQGGcQKy8umzSwPU5j7bgnmaKRsO/s
w6kgQpWehINck9PRgmorMvE8l7o5hcpyITzskKgv00FUMFnwrui9aWEaTkHwPMAkWwPmVMYa/Eye
2g6TNYEgtrDW1YVlDmltvy/OMUW4TIASDCMKlVIxpKZ76G6JAvR5lRisQcPZEvPdWuwLwnx7N7qJ
V/QPToZTF8atWt9To47y5Klc3pGg4tz3kKx6JgHnzAwjQz1bEzLkzyyfGsDdkm/Fi51psaWunn6k
o644nkui5n0bxTbWP+T9VfWUvEdfUOmDA5ESlYywK6F7YQXv+UqrAZeI2l+T7E9Qg0aO13mhQkTB
NNvyooL+bU2gfbymXM8jHwMHYmcZ0Owi5Y1cY0iHsUKjkikyxRCs1A3vosfnPMKDu4eUWz8ELaeW
u3qYkQDFaO9Bkka3LGtSfOqbG7RLDnA9l46zHXJ0sUE+jv/oMElRuggf4T0bpCk63d6Tcvy7QiA/
D7rk/zoxAHRsu/DnwAb2rAkJBWdyzIqhbUxr+Ata9e0oYW2B4ywV1iFZ59nhZZXBvlsmQ5JNje6W
YjAWOTCX50Jhy4X8seb8gSTkEXuy9vW2glHFiTF2ll6cv1dAWebPp0yR0hDCMluP4NTnabx2GU9X
pEM47HYvcQhhpuF6NnqTrjxpY5DaMb/x4flFBAcYiOiql1tZrDd+iM29RWTc3eabSWYi3I/yOuXr
eCj+MF7yY+G43K+DAggoFSLAbeA1kgk1tn3NBbfCpWVlPmClQEG2hXc7Fm3mUcTRPYXpIyYATsZz
QxOgY+C1ISzMxdZxRmcnXalZvKRaDfI0FIF0BmLGsCEF9kmyXXr3GZ2UGV7qlEP49VFktcNhqenX
D904xu7lR0gpe463ruQAoklk05eYeUtV9ewdkmyTgf0InMi5OZaSu0SK9BeCSsaVPitvnsIWbr88
QnVfkU4p+tmM4oIdya97kHO8btZCVgtdangn9bXZTPm8GhO85Fz3Wlp/Y5sL8IW13ElYTGdtfFeA
VTpXHyvW03EZeE7rz5UQQuy8uqMfg2S8fIUEc3k6rO+qZgTT1YHw8qvU/JADLjlwbYTgDk24t+cH
DUDJcdQRY5+Q7fdiPsqZXaKkpQ+ptUhLyLoQEbzmIPNfDVw3bHPwRc0U0IbRmiOZY4/Px/P/0S8c
y9wZjffqnIFPcbg0MOXBQ+JwG3ipQ0lnuRcGh7TK+5sp0hAd2JmokpWpoyW7XZeLDMcFDavAfB1P
PgzAMI2eWH8w187yxDRFq2lHJA4oooKgsCsUv7kO40n5MA8YYEQcJ4UgDURvjtgYb4DC47BlWbBh
WwtQ8UoU8NO8KqJmpCfD2EFpyepriu8BAtmMgSJqP4aAfHtjsz17zWuc/fO5LxXS4yXj4HAS0Gtv
3b4Cr/zpbGg0zXp6D3469IRGYxGJWmWb/iNVUNnc9U5a8mQELXfgnHnQH+2p7Gm6nYHG7yCv0re4
1SqyZYXOyxUUFcBoJTAi5FwUtXmXJ2BeCV/wL56qqR1VBJ0k/1sY7FGCbpt1VIQkw31D9Qkaz4SU
tUStOr6SvQMilp5L3EeQzA8S/4rkXwX35R/T2lWobCKbESYenzrIcAUSKJ8okCEff87qeIi6wPA8
2AlL2f4mw04M1X9s3eBhjL9XnTGwZrgR4xFfJzQhd3hIRLrHxqgumBFO/69YUuxPvCXkI0ImK692
dFKwyVe48RQq38NKhAZ2wRK9CjhOl8o4V6PfUxmAEMoGo3z81ZTp+q+Dkv6mJPJdNe6Fr3HxKQ0g
fuav+LkjkR7yGPzkwJvF4wbrYW6fXvPeZbsw9lsrUvq+/kQuDVwZ2nphVizFl0STa3kmJVYIxyFG
B9OJTj6I1/g1dDqUXW2eXMN1jmepZnPipvFq3eXWffDfhynpcgmlSRE/6xjfVrcUnDa/A2La98iF
NVo9OGsyaYIcGsIKvLvhspxT/3Sgv1PDlLzOA/vt9DKXjajVuVOxO966bV8jfdCRfMEkNFp3o0N1
s71lfhqb8mDZM5SGCq++DlPScd9iESA2clBJKoANKs1vbhcowYLconbqnG1Ke56+GDe5KgWWgkB9
PvZqikDRvlFGaymMQzD12Ryaulzag/6wT9TUSAVQ3Zbak6G0zNnCoKiZ8LiHbRtauuTBQC5zaqKo
CV/bKvvUz1/7/RG0tq1idd4vGn6qLlf+pIiWK3+LblgB0sHrUmdKHh16u3Kvyr25sGrG1LU5dO5B
3hMRYvwBbRNFolPZPNh5eMJLl5Epr7GTdr6gXAR2L3nyPlruslzWCRlG3ddKEgzwXem9IHjVDYEr
DuMoa89hvErK1ZgW/tWa8y3ay2TITV7d0D6ShWF/re75qJiKQTB+7bn4QFYqUMEd+hZydqP0NEBW
mgrBW+2wh6Ol3hkECXUwZVSNwxXIvPpbvh8FMYn8H6Ds8aTS7/dRysw9dAFVUHgFL2i4VDxKgsS3
1+glorujUjcz8w+SXCzM9WP37aPeTLd0C5aTOpswCxJqK9jHrMwvaEUQePcr57j6gxnqPatcGMiP
nTRf4wYL2mBKSI96+P8IcQ4MCpLNNYzxdq2yldkz4bsSYipvnWlnuTYgaLAs6dc+vZpZG9EzWvjJ
mde4ezwW9XgWDrtyJ9kcDNZLB2lIPbyDdi55HiqQ82uts2vuRmQdDQDPeV1g0MASty+PF5Z+G0a+
HmrxxYW5bN0QfjHw/iFGEP63vQYiLiATsxr0+dcH7bN+jvrDIxcjGbXh6emItoOAR3gUI57LPhJB
oO7Q0MHSRS9QNNsS31t/J3wwPsmsP/RNlS/hdoh4rhQpM1V3xHR+azcJQecJ7XsDU5PPdSxMecTu
FbA0EoO20YnyAHukb4RBWTHDrqgaZDyiU/wifFJ00oAmF0I49SrE1xsjPHNPT+ZaLSwkIxduzN5z
D96RYCidGfq59DygmZF/0zAdpsncti1tfqyeKmHXtdc1eYTRKrCpAWHw6IPS11ulefB0h/IH8xg0
JnopX6ErmmwQGz10p8JxMFJcbCW6aO+0GTxfnE7UEhrM8RK8Iqp9hyQyw3IQQmALjrCOhmANKaWM
LDWf28u2NSPHx3ZprnfRERlPRCaaBEYctu6kCnC1iGqDLGAdA+FTLgpDsXuQ0JGDN5f9deM+acsU
Pz/ZfzIQ/CNMlkzL/X3PracyqBN3FClIjwDh5suoguNltuHMtZNSs/wgZ8jFh8JycYS4zbbaXrVy
nnJNz2XrF9/6NJuMskbhb6inm4RFntiO8WNz0gD0R3hz6P1oc9FLvgQQaXb8bFHh0ts9CEBNLf4U
y4jGwwwiJgJXk4y7SJwZ6BJ0Q6+LTlywSvPR38BDpQkQum+t9DGJULR7+afNgH02X8ODWD4Q/MjQ
ymgcwZOflGi75I3k1S1z0ynHZd+5jSk+K5ayNI7bVy55Ezg+NV3PwVx/HCRf/cu9LbTxEE1lNyyj
RmDWFsQfq2tTYzIWKltOm+jUAUkwNhdW6dp0dDxuUe1oIOQHEDizd9usHLtxt2D18qZHk3w5QVkT
qM3y/pI0vXnEz5OeCYaMoVQWZct/RC8vhFR7zB7LCQZD8/xl+ahFpr5Dnm57LWEv8djBPxv7Wqx5
WzU7FfZyNaFlWbG/nWtK0GKQzWBcHX0vxTYqhGs3Z/DUzV+PyPvMZB52GJJdNX8F0O98HBAuUX2h
/k7h7GnTeMaI6r8tcJbfeCZhEN21ZDocx/6DZ1WKUVkk0rZDfJMQA467P1GT1kRTLpxO1GxxY7ke
hUcQfwjlTzQcTiN5/vcVONyeOQYsqn9V9XiKh5A7b8ycTpaZongj+hRNw8PH6ZW+DJ/IaIvzbk7W
43gpAXWW1lX5TfZKXa2udw+7lsQBZF8AO0SWUheTRF8ymw9UlTzgZYzbyv6rp76IELwnklb+tIsE
h3zdrV51HVLQkjn6cFK8LxCblVdHZMCTFPHPGXsiQRKWpl2Pe+XbNg/uTzrBEklrbUH7/CwR+jfr
Cnils32631G61XA8VBgsnlK8uTsE0J5aFsuit6HznYNbNQeu1s8tuUjfGlnP8jC7GdtlDCgIZFWE
RZRQQiTCXVse0NVFP/ONpomgTLsYC+10rhFJYKyvqmj/beSxBBhj7D9mxmZQd+be2V/VZvB1g4pU
vo2G2moWxspM6jzre09bKl0yaaObSKEgkn5/VCs/v9b9j7ljkIm9IcQM/xxsd8TFkzEnnVQYr9lT
TnRE1Kc/ydeb1BX3QGZYsG9wfdX/6N3BlMx/3zPzSQfUOqRy5vyZz8f5zAycwc2pzDkB9qyMRm2j
GeVY7BRTCFp6uNAQVM3bNbqlEjGYZYKv2kdFznVts7jk+zLrnK8ER4BDUdM6jPvZi4dHHax/pbyF
EXxFsmOfscN7uKeFhCH8lVI4pyyL90zL9GbAjtBH8hV5baCeVOrUVdda/H4NnTd22PK+4gUx5A7j
8hZbwwmYGNP+Ky2rb+9Uw2oxDWd6TP3PsDZA35vVZlFd8DEJyqqgNnTs1cFVHmquifHOCSrontET
isQRCeSKkPcBGfC6wFEmGKXAStHUeLhLO0RKFrF7BBU4wdRo6WjR7n/8h7j6OQFmd3dHz03x4x03
R2RDwIIkmadzSNQpgO0LPd70tEuig97VSMVGE/89LnmZYOXPVXn186T68vkzmJ7vbHNUMeoxgI9d
CzJ9a7uvfpb3RszKNYWq6F2hyDYGGfLzUDjo7zKxbWS3oVff9kgtrLhCYOrA8zeXxYEB5woK8iU1
FRBKZlzgMbAPCGAJG5bIfzcaXYU3AWdA59d4nRnLYVA6/WXJX++plARDh8o91kojTnM1BFc3A1Tu
EEzY3cUyBl4qbGTVafgbLlonkO0dVTptelRA86TZJCwx5bYJFZLseYvWi3y1siDj6IGYtMeD2EVa
sosr2v+BQxc06gvGUS/RGPul0Mm53CqL2Cyuzo6CN5p158h1PfeIUSd2HUxkFSjRZSyZlX3vEKXG
h1nwGcm6lTsi8cmSNO1qY7qhsIaJg+0LceBhQW9IshAVA/7NjNaXuoTEKkVGzfRQNRW1S579LMbp
CYiOcD8kZ53QFbq+rAfi4l+WrHjSeWUrRYTnFECh8yumNvcsFr/B+oiqtiIFT3vNtWnDsARKpHM6
83NOJmmx4kaymm46TFi3gDtmCuJNDJ+YJlWqitTtDbpBKq7COVdTOVXHQTVo50kMgX6L0iFX+KZl
ha5PjstXYRg+HIFanmv8xmVrCDmg86hAAOYb1EJ4tnAW/TjXzT/oKCJ4of8lb+WCGRAPDH+51DYL
tmmvm7xZK57/vLnTUWXp4HrpJ0tGqWXmEv9sN64eRvSsrwueXbhVEI0E2RLL6JZEBvlDvhRV/NqD
TEkc8yEWtEsBCeKcUyIP1LFrmGbJIPzuYpXB2tUDlLJ+jKjLhz83OsNonpLQGZ4HpXOvcdzeKrxy
fppKEr1i6dAviyOBd8/qRoE7T0CV2MvsSX9CEAgTDsuk766Ho/MwsM9b1ajHKlbgGBLkf4ijAGbq
4gTltwQ6ZAN+mExw7RtF2jW3wD3jiABEncsGc48ewnoZPXK+I0NS5kl7UVVddwLfMZDAbY6zknI7
EzFsl8Jtab52NFMGUoy+e9hGyXK/UJXZjh+rvcp1e+DHuJk90/aB/NU5kLivnw26UvmhTU19yjTE
NUjNdsv1xujTeqfyib65FGEPs9dS1F9pnfhmeh0ggABBttilGFsegbpBG3IX5GWZtaV/dRAtYIP8
7D5gBhKO1rYgexFRfkVTGkuYXUZnlEFjYeKmprbrozUXu5vo6Dx9Uaq/Y4NGLyIyj59MTO7USCzY
OFJ0HQtK3+IKVHTvWTaB0OvwZhrkfs0x9PVVI+X16eDLbHKUvyffOzZJanNEaRAebNCV3DinZ1zm
hNmv7Igz2HucmvyZc3AzJO2SzncnSDBkcs4/y51VYxUNaq1aTh76K/Ut0gp2PgtERPfiKl9AHLOb
AlPl/gc+B85yBvKmNNbT6giXgN6PBh6yLEnb3vRWh4bD6V3xCXa4CA/yyk6RllVYj7vWvcYKSL2c
Sy7zharv0bpefubhSdbubmjUg4IhdH6JYRLjqLJMX7zomxa2oLlZXb/Zy0erRKjoQlY95PG2BcJJ
ReTO5QF42kTAWmaVmtrAbPEIii74jDM2sBG+mMHLOcymaGzaEeO2vF41CNnny5cz4l7cJR/P2XA1
BrNdfl+gpoTcJs/we93Zb+qPkkKICcxrQLPsRF7ba9WHSeZHB32sA7W96EvSsrTXfyEfRBvb2u09
AOYJDPP/6vdEB+yD8vup24VuuiwDwC01SVSyfnyzjVvhjwwMoyNW3x0VKr2Vhiax/M75gdyeVuPh
qWPvMhuGYz/gFLbRBUJ3l64CpBfxpvdpI1Z/3gvrE9fjMXsWhh+hhNjulmqMnfSLm4VKotIwKdr0
B1BfxqTQyRM0zEDNQCDV3E+6L7Uerj6G/YDAKEhUJ1iD4DKJ8OPO6T5LO1J4nz/Xi/QwOpubFX3W
+jbwLd+BArTbkmPM1GP34ROKWhSAKa1I3DOQwxRTp9E8ijuon423CCq4UQuSvBcgU5QJcpvZM+k3
DgSGmrTxmxXDgzZymHyl9YD/eECYCZc283KQpmfLFH8RLIBzndmGLoAckDmtG9Yq7+s1wbRnEzLC
rzcNXnmwh7n9EJXVpD3Ea4NGjaks05JZDxtGsTx3waGRKNIjnP2PbN1P2NVwhIuo/QNoPqowCsgA
W9w9UM4aafvQ3dirDXOztDBX0rkYIU0WBWsauxYM6BPIV6MiMapxt+ipF9GB14DxvdJo2bIMq34e
pKzN00LLP6PzS9EU+qHzhnJRZzBNUss2VyFUFrP9F91wN+I8JLecolpmdveROqzGnCo1AYc7bFMq
gf3swq0/rrOBcBm+32A/i2u9MpCxvZcR56bnMhQgQuc/PChqtOKPIdt0J8XA5HYEVB/7O4sI56I4
egMhqpABf54xro3DelpmjL2+fjNxXCYP4AcejZb9rSWyP4GumjG1yJHHOF31ooBE1Qx5RPcOzK1Z
VlWItW7iNeUBq/WI5REdwfLTszEl2SKJkJ/Z1Icok8Yb+jjF/2eIml7gsWr98QMr/bKezRmwseQc
p6M3UD1pnBVzhfPWogh7/7dFSrKO6VocnQg7Tyc65UzmIelD4Ralzb5Ip0b3z4aJc3+J9WCGwa2/
7A6nQD9zNNFjXp1lRzFUoC6b5+BBDP8pqaEUW/Yf7WMgl0wyXDjshD8vKkUsH2lNDurI7HUVxHFl
uL2q7ieDjSYuJaCjeTBzhX7RPXivxlS7zyCXRz3LUTi+9IEwq0Le5ACqUGOR/1Ip86zE2kjzbV34
BFmjCyQI6TXpB/dQdaV6Xrw4sQXDQx0m5kxTHza9PHyRdMiUsScJZr+BXI+ZA4luHjt707ZChtlM
X6vqF778IRYhwSdwtjPFf2DQN10vKfHYNQZy79rzUN68hsInKwqWnxppoURUja5HF/7C0dt1JGvy
pDOdGor5OdDz3SEscgUYHwolZoqGP/p0U8O958QXUdPEMEig2lV7Zay65RnJIF5IVbllFJ9vaC/o
76qrus1qqgf2YFOPaV5XnCu6aiYjS7qfMw0IIEvS+rsR33WWB8/X/zKnBm39yRGLUQsOSF5xcllN
Kdv2f+7tDHv5jxpv5AeJb/3Nn4f2wRLPFsnMHn6D5cl4agbt9zK27L0KbGKoBa0Ho5Zd3t97Nu1k
Or6iH2mPwi0vs7A6X2OAv+QORbEBdrpt3KCcGrep4zZmmaLvd3vxvGufyWtU1LZ5SVz2kfkob1yF
EO5PreTHlYMgVrMzaL5G3+BEpbSD99xf3WtlYfVE1ALkT8cjQOzXaKbBDu/z5vV01fAyjGadFMwb
zhZ1zzILqQqdlMoTO/dEDHco7ZDTsmERku0f3vn08PYAOBOO9z54XVd/BgGUkFI3Fd4hZq9JJvCu
DkqxZ8QM3IAukOolfxG1tR9hAfKnuQwJGvZZteZCcOImYhHzT58VZm7nTKP+f35ILQnCGQgG37up
TVfsaxNl3Bc0GJNkOe43BRW4Z5QVj/dFjOUFFiX0PVVPZZlUtBuZugvu63YuAZgOs5z8+f+UnXib
ewQsS9xz7ra9LqtdDnMuW/lpbj8bcGPXEgLGChat93yHby9lSoBsAon/rnjAaGJS1o8f5yD3X8U9
lqSHHnZ8i71C4tzkK0ancKaH8JyUwOWFUQqNXEQDUYAceQbzqVffmMjZ6uNFkTknHhKm6u7Gppac
HOvKdhHrVqIXErfPXG1CAiEjrSuUsdTSldDg4G6AOfkF0Of5RBvmPgYA4wlpCsqoZv7PZmeUuGPj
uYiS2QbXn5pke5DFtMyghJGiZULEcIBWfGBVMje32PYLAtietNs/bwdPuR9HKpyVho0GmQmnlsk+
QZ7mZIRJSphN8k4upVMr6K0BaV5bHhcsLnUpG5op2XWpl+OOx4T7lE6/eCHkUYVRlDohTAOGmkNU
uo/6ba0iOCjJAWDIimYgafhqCx98ginNIckdGYlw4sXRKdGVzyxChel+X8ek2+MSEqE01kdwv2iF
0YF2XCDXs2zU1uL0stPhqajt4IIO/pGuAa6gZLhhYdVm3+7W5EWNWdTWIIU96aJyNsucs/1+uSgI
UzRYDG4HVIV58Q9Gy2aWAAWmRkarzypnQtF0thAwM78QAztfxw8VFWYJgnOKK+mOFneFRiXfp6WB
tOVmJ8accpolKsfSxb9mQDYmB+JM1CWQ5j1pe/I+HVLGhNQDV+rYOAwpqRLvSAklQy9Lq38NbGNQ
ZQxnD6n7TJyQLjTu4xD8DOv5FQwGPpzQmTMzsHVyrE71ZWCwQ0Mv/sMX8CEqqu2rnotqS1YY71SS
umNHEo/6VMNuLUYSGWjALLNxdDpqcfeEhAWBxWuCVRnZI+4nGYOyrNWh6W8ICW9WnUH5/kGY11Sw
bT0ah+/g7CWIhSZfZyL1FVSUEjS0kStFzpG+e/jkLJ2DXVZ2mltrGCUJBhGjTkFSfSqWLbTqw7nf
/8s9rV9fOVfDVv/pSU8+vxAa8OET3zgcMShy31nqDSs0XCswWCiq0t17eVTrLAl+3QbwNe3fVO9J
sr7cV7h2nha5lUYLWjqVfGN8S4lgWp96PZBHlUfllLM+oGMngg+T8kmqgeMQHaX846C2NeJcvDmZ
Q42V8xaSB8GTEsF+udqQjKxfGw24kmzAoEdGrpYmAn1M0jaEFyH4NOdMVT1m2G0qzjaXo4FCMcbF
9vvqPT05IQgWI0ep4+Syzk1Ks/pczk5yx+/zXSOX055bQ6lQMlIoHQeuuKPC2Pip7bjEI+/w8vZG
GeeKbXd+Jxg7KSUw1zB6Hn4cwIGqXa46oc8RMkGOJQPlwHiPFBkWd0JQBeZ4fIicLG3ucoU9I1Ev
7Lp++8zmJ4bcYbAAxwYUsPexm4fTA04gkeRBfpCPuzeYglt4p9IXodXvvnEXSm6AxBx3FPovg8Qg
9ocVeasJty6n+2A2MWsgYA9A0RL3EmnUQDrhT0nBsDJ7iEckBdVyBkw+RJZr28H9HMsYptX36yZG
myNt234biLkic0FEoVYohckgsdOO0FmXsF/HTrx8mW4FKvEgJhNAYgTvmNgmHfOoMPYMBqY/Ois5
qpg+nMds1wXBhjL8IHRz5VhDqRQii7+Apgt77DOo0pD35k+duh1MjcOTzNhlIT20uculSswVzVHv
mQaqLBQZnr72xU9RUkOyL/Th9NqFEnlZH54oE6TNNqK22pF9dCPBWQ2LBWL/AU1Fg21t8FE0gzOX
C5b4p6o5ap4pYcYCayHlYF5z1jkUxmxUeLG4R5pg/56AWuBUJ02C/nJgmGUAa2Nl/MzfLJfOlHV1
mP2fsdDB6mImEZ7G1ah4L/l7YlwKSXknDJbSAssVSK+ko1DCOYkLGONNC/FUZcRBN6ZysDSrsEbs
U9XDG9n9QFZWP8lzUV89b3+FkAhd4eytkG+aax3MycYDyqUnJIpd8VKgnkUcvK6zKRuKwpMpMKvy
kcjaeyQNcEed46O3obAdPQCv3+eTMRbaIp4aObuD1m2V24RXMo9wvjHEDd3zsgoS/T5fsyRXaza0
sLdKCL0Z1t0ncPdkySs6gAJ4SUHxJUqj3bU8r4HYbDwlDxt2YC0fNii4TEjD/cK6z4WW8g9v+Ko5
hipRfigfen5iB7AFH7GIQ21/jYCmkwf2ZUJRAgfh5mrfOFsbjgmxGoPqSnAcYYWXnWAwdQNfYevq
ia3EEOt5Q4nekn0oQuW/jgh8kipxD/f/+KXIvO26mT5UAstNHcz+zSylHR+Q9PHqr7WM0rH/ltHH
e15uzhGWOqFFMiR9EGftYKzacoCBbzpv0BGpxv35A+UmxxATbTaU8ORmJ2VjpmflxfeI+JsZpq9s
aZ04eFC4qkDa5gmNlJ6zHa+VmeafmTmfIxmPrbBJpyx+8Q/ii+97IAgOlr5FqrHcDZ55zWGuxWlf
D4LlfmaFCigwPMJL4fP/80cZDrkfSdiqOT3BSX2VmuzOmeqD6w0jAhXBrlWKmfygUuIbbIWK0+TG
2p1+jeQDB8H3nKqI+4ZQMypQH0u+Bp/3rh0xZQWZCcZ+pZLQAUNGN7U073ohIb42DLW5zDwhKXQH
FfPhm4CLCckzAdJ1zpZPaJsOUdajfcbX2z2uRfLLqrfS3P9lj/lu6VEzZQyDJrJfJ5+ZlRYuvoj7
WpaNGvGWeX1pTZJOZkwqzaFCVCoLzXxLKssPj+0YRVIl540yUzG0tMyMYq9y+6F/YV7rqOpJu6mw
Ux9igHe29bT2kGs8LQZyV2v/939SIyhcI487WnhP6GdSSZhu4rJRCgu0zt7IMbYY4k3XaR5UGGfV
oxg7VoCqSgganu0Sbun8ZPxq4vmGJHRLsp/5tGiJtJiXkCC/dPyQoXGPZ0KvCBy3ybDjOKUlLBYb
AaODOl94xFXcA6hH3h8VVb0pyeT9lj3rin2sHt4yDguVmYN+QmmUvwJBcUASRGSfbEDJEYYh8dtU
18IOQgqZrDeUf0jZprvXv00Ddw+4gQlD0LjZ0t+u2tJIi6Nogqg8MQ8vHuuZTqt4BhExq/W2hBKY
O1zGuTrZy1w7WfNskOK0jzXyQVSi+HNmgaWl15tOxWZxVh4Ak0VU73cYw+BIsXIVw9i5HINqUon9
EGMr/BSTZow+nccYK7732y6wbAZWbSnMjevwPUo0D2aKLqpEp9RGElxf4Rrvwm6Ir6zsoxtFROpE
+2E1zQSBTjocQBzE3uBmDnuA/wB7Enz3wGJ3PM1KNzPHgdc1fkwJykGU9Ar4EQ8aZC607WDRJXdc
TOGiNm85Ozkky08tc+8TEHMhzd4Lnyv2gKISA7+4aVMb7KIwvCeqcIwx/3CbqqctR4/A87GEINqA
OLGBrCZkYWjcGckCAaxqHfRLMl6GMwSQKl6eQu7sk6OIBAcVHVkIb8FgvKeYI5VbRmN0OEupFrEW
GL1BHrwVClmYec/ecj43TdKOW0TVefpond8Vo3K4vVz2qkIhiiQaGpKg5N1dKID0aLXBNG81oYUd
bg71I+waacalHcsTj9v39c+k3HjLwtcBAW0TV9BDSY41sH6+mQRsuxhthW+UFNgm03gGnsBM7AgE
HD8NU+6MPEjxUeTZ4pv6MHuBqurEiq3g9A1NAyOYWGKP1Ky1zUf4BzcZr0UHCJtIopIJ/PkBslbi
xDvwIk2JKAY1TtXPKmgzGCdCIen7TBrzpzGUFmCtDrDevP7YZ8i7wzPufvBBiON/AseZCt+7goqZ
clZv0awQvR5o4Gyq7Fq+7ZcCzbtXFGJby6xn97LfIqkgPdT6AwrzyR1Y5eBRLm3aXtSYi1DHQi8V
wJycjnVLUpz8ctl+sO6VkHljyyrpBaBBU7LwgXCQwATp+9ecmBdIKh8+3SZXTLgDAo/JX/nfx5bI
WJQep+OUgw3kp6AOMi+Wjcp1/AAabZv3dwASNFgLmHJOthk3d/PV9DVDTov+jdjhcIXHTVLpBJiT
MtgJpUXUJTbhLc/yPDiv+cDx9UYAWRUBluRilPO7jXcfEqDWuJ3c7Ik4cSEHF9yjc+rsGIn7MXsG
kPJJIG+dB/DMHuAU/Lwp3mXTaps19GGEzIaMBzHL4M44xVnDXg5eVOTQ+kJm1U6xSbz9KgRkEkef
oGpXL+uuu67tlFuLthLSO+Hn6en1oweyrRuTt94E2UjXVyoOdEAHLe+7zMj4jn97kDn5nzl+e2OB
mC+XFyoPQopPhlbNCBuA/ynDzNVJ39OJUkG4cEauB/Xkefoe9f7wx1M0GOXyPsVlTcOpk/J9kByE
lnGK0ncND03vqZB6mS5dTP04Ty0dk0eAxZ3Y6Ulz0ofaghbweNzt7+dWgYwiLgl6iCUuF92ft8NA
K4dTREDSGFTcnhbBYWXcp/0e+kGeEjna6/j2SLgQCIwsM+4OtiZADMgBt7EvxOJE5cCJ8hPWCsgU
6TNuCXvXcmuRtI8uSJBL3jMFiy796p0CVmXWnukKhwH11T0hnh7ILY3+EWqxAnNrYrv1Q/tPtzkE
r3/4scII0+x9gYvA09uegqp8XkVpr7aEa68b2/SdxOpRBvVAFC9MHgIiJ129prRTqZj7bc37pJoU
HHMr5DdTN7Lyf3Iy0kcjq3qQuPM7+kO5sJ2/cQFQm+ky8G4sOMHrbnKO86NLdPcMYYJzGqobH+AH
N5+59oQTfttxs+zsLCvxIRem+resJXXmwE8FxWuAn5Va8fW3haVzK9hJrsqVfvCpnLcx0Njtod5p
ZOzXV3/O55Fcl2B1hQ2bedObC6uhvl3n+nbWfb9e9/1URIWXe3xgMh5CJS1wK3Izz6vsEycG/IQH
IwIDlbTFLUYy7nNQk5vljnjVaP+zZnuEjbs/PnZRhj8V15tJGTolbvXl81kEvJMlX9jfSL7agAGd
AKXNN6yBSht5yChBiGLw9IsOLmRxD2jO11SzKn6UPr5Ow83MC02czoRhYgrQhYQJc946m6xbYUB0
Us15arcUNp1WYNvqvKz9IP85TqWhmCjvKFYLZUM6u+tpC2u2qB8tsPHXUFiPujS4tdgQ/4Dv4bE/
qVgjFTd6bEYgonv0duI2p1PHoqOu9iNmyZVSkMegz6Y3q74RHObAMKUQWCBqKzIZhj9qMCMGFeE6
v3KGgnTOKkEqUBY9iBLS54otccRxYchcz3dlBFksKDLosSwxLUouAx6DC4hVggfAv0URqnKIM+83
va96ADdN++j6TnFEfLDwzw80dCXeauSC9m+tDlG1C/U8WsWm9yOtOpLnbg4vPzAwn5awKl2ET7Vv
iAWMa1d1GCIIUohAyb0PicEOHqLZlV0nqkmB/l7wIOn1MvCVPVL3TklSrZyn3LazGjkMdTg3R+sl
Lg5TrMgxh2akVg0RDsSObSob/CjuMfL6Xr9FyXT/HwvscpWWKiXvTQ2hQlHKVYhXBFRsLts5+U8U
CpoKULArIb4rGbAlYqS2Y5Hq0LxzTRsdaWIzyfdqe/4VmfSCTC3W8viZt9TIonBcA8F1v7xIoC2Z
DWcwsNTwBcokKzWuJ4dlPyg+zWpbpyMJpNdQamIVxS3MbjlbjUFL20Cpu999oowvU/zggz8k24S1
jIYQ7y3T1CtQPtXTBOmJIcvFqv/hngwIHMkVswyz+QqFGQz2t85wHsWzxlVLMefAflrdDm4+v4Vf
gmhqE5AropkkWw8Y/FmAM/A5V3Z1HOpPWhCEbk2QFuypraS5Yq24vFurwgflPvpXZTQRr31FN6tl
rKtRQPdv21OezYl2QAIbV4c+WmVW3kGIImuaKADEMTVY97xPhWCTqxkMQGsPrdrz47SqgvbVdEWa
xAlhm5u+qENCQ2SqVebN2QTFeojAf2T3I9IwR9P+vc7tOAp0W1dK9MSBX0v0Fusyng17QBXPjP4N
6X5TZAQfZxYa+yKrVjEXOqGCnu91PNHsrW4q2Zgq6+95LhwqNLGAhqmOYdhY3B2OLahtXMcJ8PaW
04bveTQt9BjgjW4988x+l6o3P1225Pxcb/qQiB1LYv9WxUuWVPxz7DtftZc/0QPnXbpQ0sIqA/oV
HSFlZ1v50FD5r1qfjYrHuWsctUT2Yiib35CDsfIkM7583SIfQVpLGbpTj8b3Gvt6VuQG0BS8Nxb7
D/rkL1LGvrIBD0FS7+5/2d6n10jR5A+aAxF+Oj0flvhlpmg8p5IhdcAnLb8Jt+gPxvrr9Ta/gLrV
dWy8JX/p7lvAXU/t4lLHK4VmLTQ33EvSjogMESTckN9Wfgrjw1dDAHf67xcYyLd3q2lTDrGV0C7l
9KgLEPKO7LdYoUQk2AT6JAsULUnU/AuhZLpskUmd+2905mZFz/kGCbpR0N2CzohHPhmmFEx+jGsC
ypzmENWxQ/zcct3Guo3g0PKqJJy56qRXtPG/QroOFrI8qO0LTxqs+vRytFHtVRo5hIlkcDMKfyDu
PhM3vnqfC+qvdpapQMseQz4Gzd7gWGK4Ii+UAKI9ud/PGVI0EO1Fj+ideejfVs7Ds24J/OLW3yaK
ZZyBlaUKfgIbCt3L3Bh+d9ZJu386f8gQjtCDO4cVLXdZtASBDfrljBVAH4TCBOZOcCT4EIHmHmer
E8f72CqBJAZHIDnLbQvK6SWPTos/BvOAG3TK9sUPTbeX273zCyvtI2ZTdqZugDfXaoSyUb1mhdJX
8B1xcJuDMZCW0CHfIOeZPi3Kz0ScIaN+Ozr942ytug0oBb1OR9vzOQzagKWqdXAyfxQvUhaP1kiH
9lhoDA81ElIWNcLf2rgKY7DkgYCoxKBIVRU67QW5Gb4d+/Dt87hdtPW/fAJwq1Dqc7KvQRFb5PRc
x4OxijwKJHQN1C8yX4BORK5ATBUNrLhYJtp/a2e55/KvxEJ1O1mVb2aHtKNicWQaOSmOAB9hGbep
MrFy/KusBy/UNP9G/8uvQDyOaeoaSUnTQzD9ZBuMF+dUX2ZgO4zKHjliI0RaH+oCmBHEEuU5eovR
VBBPus0RMP0Y9xzjR1hXczx4+IjySFOTeKhSDUFLIGYS1T6X+7Cpkwoi6dPZw4TmYrDtoO1G4lmt
gH5dbph5PeAx6IjTcXuFiOumx8I62qdXDSNL+XnRX23XS/ZARpOLAMdnCcvi/N9G6erj/8PKb3hm
+04NrSdRRqulZYyUNpkGAabPk0U+k4m+DSVVDdyj4onp+OGjVi2NBCHyZIWLjcsJ1VuEwoc92VkE
UsWsX+f/R/zfL6jltA61ghQo5rOugAwZ2TEZIOw3v1RhUb3L70wkk16D13z2/THjb2027tnLfXLO
tjMAefSzCmRATPJkUR54L0ZCRNVUAOD9NpQPTUEZygs8IFu/tUVwFtp9WL6tSfDxgATVHVRBxAY2
NQsFOnsGXbO2BI9ma5Vi+WYD/QhA/P4m3jotHs1MJ1ZgP/zx66bontvuSMjB0/5rf1u8JNY5r0fF
NvQBjn3EKjR6OeQJroKZtA2FmsyMfAeXehOptTPa7J9oDI1fm9w8X7Dy8gqMa2AxKwikNaEPdmfG
K8SK/EJL0DoL6x71dXI0RUXE6XT+C1JMaUDnxiuXv6GxuX3I/Duwv0mr1UKPGdRdG/mZP7dHwleg
S2ONtqT3W3atqXQ9/MDaycREu6YJU8ZiNzeOkbEWSJ+zwEQjZOHUuuOTu0qkeJOzo4isl/ROoZ7i
BR7z/oXGgQSRF4ZDKOFtzVhKTgCZ0KuRtmUAtw0dbMjlYI1SkAmG/aSZpUj/v9Ecp8Zgc8Vs1ddt
IllY4xH2TsKNOEcMrjW7s4p0O/VvcIjpWToPGsGqSdzWJEK4TNvuZRTxQG5QbfCwMgY+DIOGT+lG
AbKUgHxIHNratToBOc5tezcy8o+4PtQCxe6Llrgff0Z5s2kHfl9KJyidw1jKr5lB3QiEk/ZWna/y
PVtF4Ff949kbu1r9HXy2K4IMkA+yjOaC5oW10Ee2aFGOGOsie1h6xmiiPebmultO5/6sY+9Hx9H/
ZrDHjF7ziphnVmWXtk1mqiE7nE0YMbUe3wN0j+jX0gPlDSeYi7pbzCSa1tkgSopbM6pDWrlH6I2l
AS8+j8z5d7teueF/PTqNK2mT9jBkDCa5mjUwTbnZtEKX68po43Pwf8LlH3HZiY3cSgT+aqfrDLZg
6iFrcPn9wxBmAyseiXvOYlprRbmdty5HnTL3rIGyCMYPZ0QmVH4BALgbMvqoO+thag2HYKryOJSV
PGSh7zTZLz3tZS1v9yV1x/AcPh0aVEDCk0b20vW36j9fLcaHSgx9GKziNDgwvWC8RYmET9ECX5oE
2kI5S6P0d25LdjL6KuJvVRtSpPgLoDfsHFyzWnV3FISRykSekgoMhXo5+ixestWW6PbzAD1p+UrA
0IoLkR6nmV6+zOvwCP4JqazHo/TNcipM5DtLhWmGc5Tm40nc+jdB+0EZiShOtv452UFkUVLJ/YPi
DmYf/P1k0D/DATMN9/irKEufzTxmhp0cDoeV9NSBJHQvXmyaJFOOzRaTBpn1+iMiXGL4jZUlyhm1
63Ce7p13wjJH0WaakF259YkUv36rpn1hRz+9T70BMCoDnWi20VaVa4MQ16g54ZeDk4N1z53ue+O1
lmR/uPNFtmfQzXLntRJhU2vKelBLmhmigc6mEUlxFGBEGYWq5i073KJNt8V1NN/oZMcf4XyVXsJn
YQWuCuh3V1+Kjd7H9zkEFueacJkoCxxouPqJQFWo6jz8kCMEaTIuEPIlEGvhChPgsJre4e60shiu
u68H3fuloevWPqQP2Wrl9uNSL9qr0KKgkHqyCcebFWa/yxugPBwC/h3LeLZ0nUSU1x4k3MqnIOsV
PKrlvgDVr/ti8vGVOYmFcFHqg2TPnmTVUCSN5Pptdu3Bzd/dXxeIhUpXBwh7eFE/kejT/Sp7JFaM
4o+TujRmx6apwnEffGxrNIrVpFc7cnwMaA9PgrmXxFuFnOBl5taZGgoGRT7uRBHNHgdcUNZWufM9
EYz/LxkrkBWzXV05ZL56Mu5NmhVAGIb4oKCSo6EPEFigNRcGUw2751U4riWtk29lda7j7uW3yBlE
oxMSNKMJxhBmheot+iy6HMBEvTVF80B5KZt8f/xFRyBnsFIMRgGYM+afFqQcg855RktYKoEU8InJ
ol2HfVOIynbi8YB6pufORa2wtaIrCDODC2LaFcgbjs1l1Hp0r/2EdOs12vi0XCTwaMx29g7cXAvf
MKFSX3iYjhN4bhOChnPKQpNXsyofACLYQKAcRd8gKWGpMpgFRPjmtNDAcVbIFLDswpUVS6k16nYF
bDJ2NrqYlEBNqE4sSryxNxx+BeXJ/hGC7twdBudgJC5hR0zR6klJ03mt+SzsbV+KUJtxT3lXBpje
1EfutkVL8g7HUaX4fMdFVfd0qC+KJNcMnZT9vnI1tigIHcskYBLLPG4TfMUWvTLlntu9Oo9KMaxm
wuE4wlCjpIoKYOGygbCQdo96geU7kHSAPbh7kxVvI82zt4ZMSVlpnelPTShSlzOsgf3KNWe63+UM
VhoBGnbXkTzSMs/lgvVbJb1hvoCb3QIfeNNLEhbGlDBtAEGcQ9QBuHfKmqd+OoUKaL/wbotFvQx+
4r6KerUyIRcJ8/vCBsMQvRYH8Q7Psf/kwu5O188oVa004vbkzEWHULVNFB1fcxAxmDB7mhCkhuA2
9i/k2asfwgpBVwFldZOVuP8sQH7/dcta4IuXQzVLAsz6/PaJ+A+exL6Ft3Q26CaRLLy97KWnI/xh
sSza4ucNymBJst8I09B+a5rcLR6kPneqFckw1nNaU7oiGwzerUFrwFhwoEuaB6Tl1zS4rJQ04Thn
LTdUoWi8aJAp4JTE9pVG/e2giAWXQoW/FORF3DOvacrvcqpmQTu4XI6V43WsXq4PRZ9+T6evMg28
lI5HsKgFzxOWZRagtbxHcghDRuXRBXm9TfLgGjKUWju9GyDRebXbnLz0jS4whKgBqJ88OeHqrHmj
5P+G1tGlg9f+4aVpEyX+Lkn59NifrsMV4oBGaAJfEUA/nuf2v3kNv66bcRuBYOjMXcszyIe+5emT
o9J/y71xCnwzVZqh6ALTRifFN/BDTHIxdOUY3RauRFUOGzRC87shHPmosWaCKr7LEFu6k/cLSh8h
lO3fL17GVxmqH2qq7DCE4dEPu/c1ltsD/Wvnutu5wx+eysJSgVgiFUIiAqQGiJXss+I7uEgZ0y/Y
57mzeqah8dhlLNfwq1cnEvrjlO3qhwFj8hLqPpK6Cq4F38gvjtzFcjbNiVNYDWP199Hs9oC2B8Qz
8xHEmdiXovklXc2oCZ/aHfD/kJMFPVOOo6kNnTHjJMPFBYI+xXoqE+qycAjBT6H6x+9iSwI4aI/0
Yj/v6dLE5w80JPCFPnx7QSiTUtLLhO5cRgi3Zs5yqN1ZZj2EGGYhXmjjDpPVZbzzgNlN650wCY86
CdLTCBm9Vvrb4sdK619K50aBgcm38ZxIR6TEh/KxXrAuCxh0qgtJhUxIKcOXiR7QaWaAzKUEBLUS
0yyHmBNwDonaXfr21jFT+lEA9qMggzwdSC9He2X90U305gK0cjQQS4sQugFMFqc6SX12IGs5VToA
0iLcw8BM7LMZIx/FQth8jV/+c8z71KfX1Qmz5Et0UAMiTzOez5THvawL9VJbeGnsp3y2yBL1QYf5
fYGq4qpLEhDWKB8KQ/3u9OCeDUdg1o/RW2xFd8DyHiX8npT4uN0q6eVykeB8T7eoLXY9T5OgRmS3
3HoHeZHou0SXmtKBHygHxUx9NAbHZP4rJBcoF7ZNPJQ2vLbqpbPWTQRQ60w82UAtebmYLifNq6P/
UY8AlPjnzEiab8Of5PbdYCCdMoI80OrcXrs3XoTzQ2XGTDSnIcEboYp4hVxAwVaKzPnJ1ObA+jB2
1XN+AFYsDut92xJrdhVduXQPNlwgRULnKGAC7dwDiVhhciPttCSuBPBMhHBOBdXChx2/WKjeM5wp
uYtAd7SMhIU2AV6Vlv9IJxZxjaqYeUa48a46a/Tj1jRgfnB7nGz8Vq02DI8T19PODFqZxMJKFuOO
cj2E1/b6kz1rww3+wubu8WqLQ2fQeDookdBgL4NVun9XPFqwkwCRTYvNTaxNAZMAgWg1REB26wbV
tLey+BGz3xu0RTAYJWdZSKTifgrVKsHmWVLI4aAzHWKEC/k+PDuniQt7ij6KCIkOblCutZC3ByhJ
Q8yuzGTq+HBAnWwxgYvXbigiKRbnVWzcuzF5+PM4iFW9zgyJtz7+ZAxskWx0Xi42DsPOLbTCOfbK
n2zlMHJxmdYAH2h6Bu2jIcBymLgX2AtGdMlI+tJfxvzowLRQh4LluGCJASgxkvRHhqOnFq7LNBlR
tfNYpAWfbb2HeqhBu5vX9hjU6HOOivPNhOMvwW8T8X0GKYDNTjA0GqKSZCLy1xlorqBATycRSBeN
pVomXfzkkfEwerU92hemqwXX2asKIP64Tc7lDCuLGOmMp+v09NGlT2zXjjwxhuPmLwZfXOTplCU4
3sql5SbzghynXFdFH/50GxqYB16qFpUd+rODmJWaPYhETwjJIkJb5fdBMBu+6veBT2nMH7ZXVM9S
8CKZIiVb1YsFmCR95Wv6c+2dD8gQPt6mmFTYDHLDmXs6mTKcTyUaX9Ty0+qYhyFbSSvpJDZ3LVie
cjzMMSd/8K4wqtjiYpfEX7CblzcPpAO6faQPj6Z7X9I48NnHchVRmThGIA3cvJMTBh7vWU61R/5T
yCDIm1ELu07pTymmKS5hqh+T+iVWPCqTUMqPtUs7fRY8XZL7H/l4T19tTFg0i0EWkkvMzCDtJZ4W
opwpR6GABYU2e8O4Nl6PY1q6v01QLfM4RoHWcXzht1ZqyX37DYFXd3ZLC1htjAp4AdCNFoXmUGq1
LmmdLp6mrnruj7kAPYN42xFd0sHTdui0wNZY8lW1PKgff8Kk2uU5YUNwoeYZq/bzfO/B1eZxYjH/
QWOz3N2aw1PcLNU9gLPbltVVqvd4ooAgCI2+UneCXJxAZGRw8yiImcdvEBlmyXOzoWx3WNWqt0L7
PUofkHIthISS31TDDOnO9p2d1JTLNypDOZEnXzZb6NJKl6wdHt6MtOQm6/9e7isy6SgK0rRUc4DV
+LYxUrObWoKKgxz9n++3mI1LBja8TyAlUqwlkT4jpQXj/jyl6qjNnZhJ4+vElnkXnoCwuGCkPYhw
zELPoOPpy7HqAdazW2J5MVX9H9veI9b9n9G+6pUM7YwgR9dzfGrSgb7fufp2Rm6MKmJNzFkwpcKJ
e7dlZQAopo+CJeoQN8Vg4JzsFJf6c6dDgbjYvFIy/bdT13neVT8BJN6qBriNP7jvQwJuRmQo7RPf
s8RjtsBwRkKwRF0NB2LldBkmWrTp7KxZoFMefP++GMsgqEAKmI47MtZXsTtOVAXxHFbYHckbUgFi
ENEQxmNYa5RNFb7+F8prVAATABcCY/3Tu21yp5TPDLw1/pCdkQhP7PxRFkmjA8VuKOUIamn0gViJ
RUuRTuhetVY00BkMV52Ab49qGwB7jLprkQhRqo6wtaLCteqK/sriQlIwwH9+txA5IsfwyPIM1IJ5
0U9b00i56Ivh76kjdPKwp8ijNPgvKOx5jq7Y61ywoWELFe5k3tmaxUtgaU+03jp8XUz4mkGqdvJl
mJMyvw47L8zSnA6DTuJ51hgrF0N/ob7TLlYZEJWTqb+nygyZRwOJtwLQDGsGQ/pbuvAOjuDg5LQj
BJk4vY1MMPNYA+1iFU2AsZvA0B7wsYMzN5piY7HJnOjh6BBuauRLaKJNlrQdFAjkqKuudSOkRT4T
uSqcS0lNQ1GGszd+4qpCCOmH3rccep6qvvpND1kYGw23SHJUtIFBdIV7tnTWNwRufxxKQPOxZgcd
fR9JCWlkD3NlEGBiQCN0Hp2G38glGt9UMsSXFqbuPM0FZwtEv/Dxa3HWzA5ZjG0923D8fmZhWhnd
lYajqDCv8e0DVzuvCNtMOASgvMq6Hk4aLbBNFsxGRk9nLDxf8jm1zFQHaIOF1S3HRhQnXPbMtFNH
pX/MwLHr8zrH1FWdBA9HavDvLtZq5xDrvfPcMXM1zI/0Mh5Gg7EvXh+2lwF5eT4VyTXddb9kyjBD
nwSJMBLgVLqu1XABZYMi92Y4MANf9nRGloC2bFpewct4iVwOtiI0dkksuo/KKmX5MinEqJx40gLz
apjW/KZTnozAKcJHTWrmcev2QVpT0YeSNn56Tin7a/2KqN1dgktXDg8BcsotFYC5BPFna71/HM9Q
XbyUriTlKdOGs17C5FH8XEfafYEP/Kur+E2ikMO8bh5egH0quLwFsRV/lUXTONFi0FgGyV6raeAV
n+rS/7ZeEH9dLw41L2dkAmiUDEvg8Rg7S2ofuq9pSF1fSIy0KuEkDGO6z8AvNGrbnbSpN8F2XxQu
NlGdE06dSP50HYCZ/r/s6A+q1cQtSNZ97djsZ1OWcV38ods2L6xV6ruIsWjOJ5KdUzXXunMnAIWN
2mZR9XiSCY9sWo7KHJAshuCP2muP6v17p2YauoL3Wm3pZ1LQH+odJ8vQ1oXufW9Ohx7/auNUKhFS
29aZBk2ISXM5hihFBA/7bABkcAupeWk286nLTpJm4B0Jg74w+AWASLDpZoHXHc8ExdlztVb/fg7i
uK9JYsVT8uPL1/jBz3qX4Ouh6TL5gsGijJ2cmDQw2rFzlCsIO/tjHlclJ4gtzZnTvjB+H/Flk8Hm
XGApqGe7HSU5qJVU99NnoUHZH9AwqvdpMzpVm0h+CBUfo0gBdo40M6+izNwgteTMNEigPo2piiaA
osQZyoS5d7FCVF4GAvfzdNqGVCU0VJ6kJozXP7jIAVpLMNr1Vjjb06MtxYC6RvYWXNYiADV/s4iV
EPazZQ/zecRGFll3F9isxed9jjL46HL5FhkK4gpZTA+x+bpJyUD7iDhySbaL1MSNX2rfbBQTWSEj
tLoToH9uqt8qnhFZhGafTLAWrLqEDhHym4eM0wziFZ9lXAnHwxsVbq+bSPl0AeW23032y/iBZX+p
sIFo9UYiqQ/O7QZHXmOUN/TbFEgPXfSW4EVbdCjMzQ+hO0XalXK95FrBcSwgqpifeNfhrqODBbsm
U73YkPoyCFe+lCSeEyoqWal1ZvKNXJUlRMxD+zq8mB+ZwOxT209UZu3bEL0EP7VOE3FRKkyMkNO6
2VEwtRR/Lpon5/HAYb8UGu/LU6ZmiD/at1sPuhvf6M4/R9AUwPDIJboLBUu3oe8DN4F3PWxaUbb0
09Fk5HlBEyjC8valw84vAz6cowbRgw74pedjATlKxcQn3acR71HGc6C+DbYH52K8wQ33rqrsAObC
Uhx5250USVkrAn3j8SgHDr4Ts0J8OCKP5vv5HDPLma7WAmlO1896agI0wnZocHa7DGfVbNlQq5vk
5ue8Xu0i474mf/D/axYTUGlkZKhZ5hQMGdVY6mYCrqPt1BM+0P32nxjknpW6kgrC+f4UeiCgIUtr
eIEVru9hInwuF8Ip7PyiZaMjhsk0prTh4ctimQiBh9bIIJT9CkDodyq0SdYgbIZjiQHazZktV1GI
vlNpwIw0GeB4lWKGgF/WnMbc0pXO9iN56EHM42HAtWHNAQ9HFGHicnRBbv7KYvVn+bkIoSHI8rbv
mqn8Kei7DmTMnpH37Vk/RAOEieBU6+34LYsG66xqGIcAURXqtj83wmgs6swan0uEZzwhrkSj/tTT
UDgXCzOgVkDEU8i4HFrvAxsFbRFaZk/swWG1IAC5/+NvgMdkIq2URWgjq9n7CrkaHtQys3IlPm0D
r7BaIVCimdLzIehUaQRUWf9aa3pDnB2nX1KTZRu5RpBq/z0eNxqMEbyYJZrRvpHd77tuynexQ56P
K9WYksJ0PheJSbb0A2OYY7gDrI+yednnqYdY2MwL7RmOfIQxTfv22XIPHSCWYR5Agky33z01KGSv
RnV4CUGZXzDioUKInMGiua5r/Pg0o1nfV4DxUziERokX+kyPs/snHam8bX3FX/oV28lvMHvMb/cJ
Yf+S6I6SIiTh8JH0aSc4lrKtKBVlCMB9pebrmsvazqnkdPqmYH80EeQcW1G3IjcX2ns1vPDSwU4r
ZYe4POedsD/iWF2kz9mAoFylwRLUsMj8DhUkc2vVSiGGkLwIT5pdOsHGJ+qCfZkta+rG7lYb3CK2
YByW+mxNVdkKLyzNYWF5VyR65lhPnF5BXIit3YY39jpomw7INi9HFx7OJaOBb4S1R037FYcBKg/n
jgFFMUc2/WjLAwph0W+tgUZC4NwOmU4o8X7/P6N24XUVVp13TAqsU34SQINK2+mouhZ3oimXpqmI
Ba/QQ5HXZwdH/yIH/pJghr9wQYvnus9wWsb3GQCdWyi4LitEvaN+x25mnA6o2dPmbGbOJJ0KVf/I
BpElqW9+AWCFFOWOUrkxezRBnzelZqloL/hxpUR4SCZCQvOAQLPGxJdbnqJhem99BfdWIusKWZVx
5ajPlRXFXIgT9UJYbAK1J0l+oI7lOtlgNnLZTEH1GSY/LoeIO5RdN79qzYrokKtRek1hY1L3jNxP
1d6WtBGdvcGLoUSg/U5+jiViSEUmy+cyvvfX6OnZNB9zmwCDkdilZuXpsDhdkaJWEC0pi4c4CKXS
+2pkxmcb+H973aw5mk8lpORTL4zKZxaGNuecJeiLu6WGu69NUqSLPuPkh/Tok6rdk/05o755YiBp
GozMhCwEF4QxHYzE0HEZ9QF94bLnfeZVCfrIaOPojGc8BzqS+b0A4LhF8YKLTyHvNg7Gt26z7cRs
e6CVVhaldpwoiMzhPPlOdH7hAwiEM7N1HZ+4sCOwVx4suFOiuMjCRgXrvWhT3i/oDpBRnjaW5CtA
lyhZRN8PoovTvJzwRrw3RZMs3wfKnB5I0IGiWP3yEMBZ8LpeTHdS2Ln7sobsQZonDxAYnyIVb+zn
qRMo/uxov43Fhu4p/vXvysDkDmBp0ypRXaOqS78XC2KxdaCQ/Q3Ls6kX5bpKOXah/dD8WDTIStHv
ArOJZQdQ7Rpx4Xp2qdWeeiVp8z6trVTVLQXOjLeBqjUmQBgKX9WfpqNH3p1gI0IVwdcOcX8NyXiU
rFmyAeJDwoPVWM9UZrhi7ltLkPN7hRJF+vxb7aTLo9hbSJntfa0++d0XpjNGxjr1RWJQlOyBAFbe
xRCOkqGda7icDza181DyCnM93sULD8X8GftIJhnNpRLL6ZSBzrv1cD834AyQNxF0+Y9c3+DFBm6Z
ps3pgkDMo8Xwp2q5zOCpxEnTzm1+zYwBudqS8VTwrD0sxfpabq2hxV0EmGApbfo5h2ce+vNCUpib
nPCm1nQaWNEC1Tuah9XSLlJomEgGKHGaqNIp8iXpJ6AjQFqnaZ5avS4UwtbUkTRpHOow3F4p8Set
b/pzWFpchKbHgrREVMmtkz29NB7VQzR1vnYH2EGh26QEyvRt7scfarL+0ZpWhysjAUCW2+jcwmtg
RPxn7diROc23gG+ePBcAfXaKsANfaF6vQAhagiS11VXEzajb/d2gFOpkCkBFqi+oIA9AU5/ocBEA
RhEG2dZNv0GntritwQQQzG7nRzvXs4AR5l+LVVS2SmdTZrnMTLY0c9cLeMy/KKOBJo2K4cJwTrFU
aqTcvuLrtToqn7w8J/i3dxMlhlcw4KMZK6wadWEBkVvd2zIr4mnHPPRaKzSR6OlqPH1yBTaOdwAJ
8N/y3Q0EnQDXpy19YV7Cqp9PzcG9KUYCwwpOBFGyyhkLpGDMpRG+1Vq8jIPOCSeRepdIZD2d+euZ
v6OdQQfWeXHS0s+vVxhf7fJwJHryPSlD5Vm7oxdZ7Z1ZuKBPzy6erN+9rUCRMOnu8m2sa30hOjr7
zNEtl+gAkF8nPvjZfaRuVnI8USXRVvK19lFfpvMNh/BI2ubG4rLX8Cqg3EBm3pSyjkHCFn5Z5nsp
LOXBS+B579WFFm097CeooAsZotG8aG8ITP8wNsykXrWqUyTuF3b9BKEZaSQ9cQ9pa4T4RKIF+u6b
nFb9bLSAkBY0lGjXu87Ai3YbGdX4Qwk0bdnRI4aKWhPS1HvsYap6e0uzeq5FEna3vyzkPnO3DaNU
oeCO5ZhLA4Mj6sM9MtuigzF+fJag1/c9tRutvmJ6+gB8BWJNLCThLcQtAoo0OXZtFZjVuHgdLiE/
3HJcDKF2+DTnaEv10AgzS7GkGO/8Pa7rzuuFXrGUsLV1Buh8EwaAa2Bw1KC3njaZemr+/EMvnHgG
cQtflqwk1/aLU/TAozq1B2Cwvu3IFjoGuG5bA8k614vVzzgpmblX1MkSXizokzUia1B9LpWhPaFQ
dAuYSUEs3+pwi/lPrIy2zbYm4p7CxgWc1HNCODTs4yMEspIBTlU3WUfcgIRoQE9uyZBVsxstWBRO
Zo0SUzGNNAJssb0R9jWUvOthqPr2H75stylzpqTyo0ZNA3Kv4U9NNq9QCnmmazXOC72WOp2e9Xi7
AgjDMmNAY7dMPDaS3DKp2McdpCipVoWV6FVWtYYpZRRuTgvRcnw/v86K6wcAJmAI2kwitM6o6QYF
27/uYr+a4JVOsya8Izig0Vc/c6c5MF/BSaamPNPRkykY8Mm0qQd2umdijo47kv65bG6zs1nJYRMt
FJSUTBrhsQx84HUQNTPriv2+NO8ZSj7nEheIDxtsMyfhFPOrg1r9oecxCanK5FzvX0jFCgSqY0m6
6ek7iUwVS9ahcJCAFPZ6DCtltbZWNlKdydF85ZK+AZfrb6i/TZi5eqbibPc9jFdCZVncBdi38X4E
CPw/zsNWPfXEriU4mhBPGWKCT8/khqAA+OzZgrwEQGP7tZbLPCUFfX4DWxRp3IIp9yeOjxS3rrOO
XwSYlIgjam6X5u7Df21+SoEuwQzsTXFpngU5udl3fOeiNEjYw6TvGdAYGublLPqi25ILf0Yjqhz3
KksaUaQVvmhbN/t5HK7lNRa7d9ZCa8TxqckGP52oup7Q/k0xi3fDYRDMJynmSPObU/B6zzN9ViHf
aUlt3MWepx7usXkQ0xsjwztPsoSjXFfLVkjLqDkjjiit+h1l+xTjNW2EWCb2g9U/zLIXGpxNenOf
1bCnd8zbi4QHQ/3FfNhs131XxuyH5K9iyMF51dN8cvddSt7zag/o6sIZd3fzx5twlhSIKgck1WWk
GtDdqheucfUP0u+sThhxOW5Fqg0iIV+DZkVc+byYRz64e8CCDPGEITIWEPHXX2TrM5yXjDUUPutE
ULmxYldLB88oSoEUoHKDQE6i6cXdv9GfOP72guzHkm15VWzNUwPdVYbSu6A9RK1KNxMrSJHHk3cw
s88JbsEwz7rxKmhHBCwqijmM2aDBrimvgYSjA9cDwEUlHZxQBNRVD9gW1IkV++iTb4VNZTs/Pyrn
ff0NN+za70zNBs7Bfgz6rhdN1NXh75y44KFIJ8xQBDT+xFI9r3vX1dY2TdT6mkVr2X4ht2l9PIQ7
jlFTOxIIMGTUtrvsicitjVkKLyXzK6mEl/p8uiJXru/tWb0X667vN+iGWcgV1KRet3OKTD3Rmgug
kDFE0Z14/285lvFGIxABE6OlmXVjdXKaA2k87tFdW9EvUXUPk+XSN/kgrqoswEFlAvdR5YnXxEti
txdTRt5bI2ziVlgMqt0xLE9uu+fuw7rBeORLcS+8gy9lX+2wWMTG8Sgy1pcIeQblzudkelxp+xXv
FGEE2bXtLuUCK7yISbnaClnMQNxG0JL0FWpM+zIMJDjKqiYJv38DtJ21LzzDBHL7DvRP1q1ol8Qy
STm/tluGUHtB+WvWOY3dE2O1ivc3h6FV595Xs4a3IhywJb9SIa9ZVM7Cvt/VFt+YvQTj4QLxeFQr
Vg+aP7yGCZaFFr2gXFWbXYDSwXJrEyiZTzgBWVrmqLg2sGaIwbEMul1YuKIs6dg+cIze60wtlO18
ZdcsL8dIiGepWuY1jiX8PJNIwW9HEPBd68CShKUtmqFo9v2Z9ljubUkE7MPbblgMEed34p5uysTG
txckERrnr9+89j01WR4PO0S5ErMWQWGkBQxtHyRPdrVEUm5uPjGwb48yV7+NQFD11uCDcFmhuKzn
CVZZt2pbBKfYYLkbWslYqki/XHbPogW/qXL0e8lIcy/7wJ+cTivOrkq22hsy9QyJWXaTswBQEsXo
IQGUjRyqUZJUmsefNBxDZGgMAA77pvFSqxEqyyR8uWBL0SFQHS2zhVNDCn5eGkBipLL5y9ZISmyx
1vOdbzAtKm6i0zYvfKs7xvr3b4VMqTr9Km69VhU/2LoeCTRZygRA/hmkIfFTIVeeEVbTu/oX8Ord
5f2Q2ccLr1WM8Ama1+qwsp9Mc0ud8jVQrt7obFL22OH0q1CqfdtLMQvGcUuonjBnk7Utr0+BBcKm
0zNC43VkTUjxFhT8CwoQv+qGGrycIcdN/pyCbvGzb8IlZfQlJYyJVZ3Lp93iIjHAmCsvA5Wdhy2A
JVKBfjIQSgqt/EGxe9Kt8nw82iXxEcH1h+Sa6fnxfvKBaSGXvE/Nv7ZEQ/FzxxQpXy8kk40S3Cz0
HHN/QFVKgCWx8jb4mbz00N+dPzcLpco4xj21t2DTewC/AlBGn5gR50FmD2wpsW6nwbhgAw35e/vG
5SCDX5Tyd6CfytjWM4420ojdbTBPv/rxcZK1gdHJ/hAea6pHtuU0dkIkI2wUazv5kXsfNZvZ8kVN
uG3tYx3A6SZYbvmjUZQ8hmmAR16Vl277KC5zcEnovAozK8ZN0Ezis4+OAY1pp5Ym3b9CkM+x557N
8oa30CyCJ26Sh4Z8YjwVR269Km+gSq3ep7lkYiqBL8kMsnzO8n5rPIWNE2v4eAAqWqeNf0iqtMX7
7SmFmbqRbqvRcXIG0DYRFCtc9r2Ph7hTzI44zNnlwq2ftsVicAFhWMYtRQuhx24M8/0AnHHPYY2a
4GOOXXu1sKQjsCexILU6lQVqOj6eo0aBytmG7ftEEW5d73fexZahuJxRB4LtQiUNMtXU9qEsuThP
mG6kDX+DN8tI+rkpsbLXA46RMc2IxYS4ZpN5p1KdVl/dbJAuSLGMsHFGaciX2dGWEYEtPfGJ2n33
AjKCdii/3NFQe+WEuhgJ5KuFqMfn+1jMOlFYqsP6aFoC0GOqw6G8vwESaUr2PodUedUapEEh7EEt
3NbKp6huyHbgY0SLm9woq2XW73NzWT2D+sIxjAEf/dw1NeLyBFID6ZlHmW05oH9mMuxYucISlM+4
j6sSQC9++8Un4qGQPueJbsAKQf5cQ7IbV6k0nhk/KZ+vRdwQNg91+Ie9HuvloJeHqi7SU1SVAT2g
QqJB7yKTUjAdZf6gwk9rCBAMztYtIXDkjdqJDXFam6NmS/bjLnr+M6CWgAQEd9OTK7T/LhLjIyhr
+PAyTDSUd1Zffr1x9pnor3DgidoZp3eqR4XGJGIdM1/QDx8N0+E8szU34Jo9kwdw97tiFihOnCeY
DNHFjhOmB0dVAKRen23+3Y43Dc/C0OoRCdz5+3WGEN+9EeRGmo53lZNcnZbAB4u06/LK0go2vHnq
ChMXNQqGYfseOnxgZfaNNTLPmRPJONnGinQdXaBb3AK11qcJvLMxb/BI0EBqV1ED79dTZdVd5uju
+G8Onu9i6N5Yw1qSStlQlCgFGM71vH5PA76CzaZ4bKogHXwP9WxKkgETVQNx46l8C+K2VLvHlkVN
KorxFpF71gZ3P0D7pNueJKSwPnfhW/tn8COGrF2Bk6ra5Eccxt81EqSs0zM1ZhSKy9DCm5ts8OK0
s6mf9iXxp96otC4vRKlv7MNgZAK4PipPbVtasPjkBQkuofva60tjHYiXo+d53z86VXTlkVG/fvJL
f7TAyT2lNXoqWwCM07Xu1i4yLq15uxZu+X1Mce6f8rGcnFWjdgWfb871+//2jIz7jomT29SjFPJF
fw5EXu0+fBZz4LyKmm4kTkhOKi201lnS8gLMclDrlw2vTYENMj/c50RU16zW/9oD0oId5n/TQ8zr
1WTk8HhkmwDR0327FqKZOdjIj7yY/0bXznhX6d42mJfIlhU+hvC/PsJ1ZoYTWCXyqeZUfgyLQXqv
uy+vqk8UZ62fzKcaXEKJrGNOkn5hs3IS+fXiMYzoYpcfnNATEDAkHEPezzs8S3TKEJloQrPrVM3u
ZR8GttukCFGgIjTiaG5KexTt6YjUhMx18KVg67YCdkGMSpasUmbaPruz405AFN5ORYZNUJgFF9eg
r9c8IpRfX38GCWlnae942B1zNebyZYDMEi+7GhO76OWRFHbPFELtJ0M3xDi6bbNww8y2thhLRlp+
qklvVvkDFC3Q0EnLtVTwqCeh85p5hL/l2iWvv4qjIaDSeozHRTuitx2tBHBsy7QunmisfmXqRLM7
vKrBLXYNkitoRB8yUM04LfrUlkd5EjReHDEbZK/1/uc8Bhgsg6YQO7cxvLawEdq5MLyTAih2dJF7
ioWpmaD0eIN+42y598IYMNe2XNTdz9L3oDmhmRHfutr0qOxxhg4AxSJ89Y1ly25q8BOP0WKnhroe
4C3z/t1LQ80yWytEx86CvAf/oAiZhLM5D+b/sLix26qkOPjjlKQWzmwjXUNiqXQyHcL7dhNj+N/I
bYwScvLdkL15vOO6f15IW82A6kk+x0GyI2AEc93+06OF52Nw3fy7FEis3YVSHmlWCpcNO6v6CVFB
di6XQtM8TQVvnPqXEp5o+wexdm4yCHfPc4Ot5be42EPr+X31DflbxkOERzDW6teI2yW0OeHZ1Air
2SFQVg9/BmUg65xMMHR0Mc87wXJR8L7Ml1HNL/6K2m6Qnv29ngWZMk9dt6Ipo7B+8A//qfVO5Lkl
HPV8bV3gec5Rah9QlDXnPTrhQ9WxqdRsFcGxwG8pEsj88uxjayhrhPxC/hSVnwX5oKfWFSUIIF+B
JjJzY7ZPMNuas/8pny6a9v4a/nlU6y0ImYb3l/RcDHCGVB2Tb1fiG8DgZu/BnEjrGMb+PVU0rV9P
DlXQeXrsksHLuKtkvaHACEEqv6k5dkDaViTEu7NvPw++D5ShalOhk/bOR3dcYyhEFHSRHUTBirEq
tfn2xIF9IxxzeukqJ5N9nKnx+4y01it0GtoNK6CtHAi3s2vkuVGHmkwAzZzT6jkQU+JixJyoM+f9
OE3L0GIsnGBbmF7LQ5myf1WiN4fksXZqk48wXbgUWz+HcaDBqhV3VKrwU9smpGqQ3OT/w1zG7sw5
OxiJBOeFmMltVCHJcVgwAfcTLveX5gMbP9m98KgtZU96+Cjt7agrVGcBXMV3P9x58I7q9s1nLVaX
xkmGE0owLL0Zm5YdAcMp9wypwHCTBPpC24M0EasQgMdakqwIPpBRLcTkrX+FPuJsDYrucAQQDu58
Mj7+reGr7Pm7E+AUfAKtUroajDUdE2YLI4rBUil+mIEso/bxm2HU0Z1l3x3K2PNbHNWPKZfST/mg
e8L/EKlFfnN3a31Wk8EkhJRM8gAiP/4xSH/h6QMX+QT9Fa/W+ooDOIVftHu6GBZVl5idyxagnMNR
kIu4p11Bt9vQD6PIgK4OV2M2ZrmBbUezZHV7YeOqriuDmiVZCeyAdsrjkWR9EGC5KTwgLQ2qrNfG
5XQa92BBwe+1RoAzkaWmXOPRrGBLoMr6B1q9I8sT4P4hTR3oDbUGGdlt4gO3IfOuljYhCHLEDc4B
P2MF1ARKQXt+UqK+id4Jk7/Xmjkds/VLkFnOV2LdpApHCF7D1OsxqKu1jmVZN8/ud9LcxNj7hZqk
ixc5ehLsoqe02JUC3g6Fx08YVHFUPlD2JpHjb2whbUb7mPz8zjbCI0ot6KDU6NO4OuDZtofvn0qp
yESzBxdL8FeHiMDWn4fyJx9ADZzxih0ZizqYMNDtsUWQbHEniWercw828wM+Rxg6VOE86id+kApS
112rRDNAozu099YsIVzb3Nig42+IZFw79hI464FohLoeUgs98xN2MvNI3n2GF6NJJzAXwkSCh9ds
JFPmEPSdkCMwmiwt/DZM4/bmlEx3CXOIuoxvYks6RNFKD0B3Dv/iJ8JSPSLW9Q+HEGNdXmXJuUgK
u17MOZqrx7NZWjILv3YfY/uPgafdAj9BQKO1e6xUgjvEy9JXdCz+rycOxs/ztnrh5MC7cu96+uMs
4odHB28VKJVPlJLM+hDmqi4KDMzzDG8rNeuzLmOmwVc4cAcip901lCHVMQCQ/pqeHlPl6zb+7VVp
oxH4V+kwnbMQebH1hzq3LIOMfXiGTmhYgBSJIjVS+DGM9RCitTislG9XXe9G1Ry+2aIZ1j1DIXpS
YQyZOxRExxOdgwyReUrAoQ7CPMTksSUFFaurIqeIQiD9TtPfsBa1EnfLZmu9jeMtffxmmJUkk2Rs
cdJ98PkLo2MQoEh+6KAd9ziR3B5BP01EuNiYgWMQMZcIIwTfPOEjm8a1X9xWVA1UPF3ZMHLRonAG
VsBTvgogIQ/biuxgWbZ7LO6gH392r8043Zg6EaISzkD9nYsNHaGmTGg/hdp+NYMjsZ+KP7ScDIGP
h17/KOt5+Vxm3PETIH7Rzq1SViH2fpNtnmsQ1MjptnWPezpgIwYAt4AxVj2CphNsyfy+ozZQtbAt
PhisPLwZesc2WcjDZbyU1U32SgJSBspge/6LYaU7gpiSZ1hHfks/lmEvjmVDIeDHNA9VFb5zCOrP
exEn7FfmtBBG5MTq0BNw9a6znDL7w6hr1ytIqQoOXMdrl34mw/b+lVIGtI396Cp9Qho4TXVerb8B
seFHQ6GkHE6aleuInTRRX+56QqW++OoB/MyheWFzqGYKdSG5ImksLfAXgIumXOtstLI7Xbm2K3FB
PzMFW/REfXc6FoTk3TpMpGLzFsBMhU7B3jw13SUtvcaBdoIjiAmn+RAqXAV4nTrIdxkbCT5GU58G
FKPj7cKQugz4Ggr2ioJo3oSLJRQPU5d1x2IN1q/vB3POZHgG6FlByilk31fXPcsAZZ9CCyGkisVE
u9ys4uQQBTWtV4nhACKvUxq153iq1xo3fiEk//lKMrJlz29JOSm2BeNpChw1RAqveaW3sCvZo4Yh
ai6qfbSOks8HwqCA3qEdv2OxI6qFD8P+9+QU11qoGOkfpfXyhCLaLVaa1Ivgr1qAiQVnQQR3hIfV
VQzwjrxvU23ofxjfmoVOLj56RPOUzoftnmmFWmeWKDC/P8GTImkDWYPSxQskLkjea/vVlkTeqGTz
STi9l5SzXZa8qKi9QY5hPvVT60L992Rz9bfaI1otD4MnIlouqg9sBPsEJhKbPzO+f0cl2J7wiQjC
O2+0oGZXRVeROT/zwEPjViYmkLPjaCPfAK41FAbcvbGY2CsDZqaKbx01L0xNpaQuBbJjxavWGz5a
CKoTRbWI/6Bf0AqIlyr+FVTYuh9D+8bJcy0Tf8MEP1jb1yAFUI8iJxu8V2kS6HHq0SWc9825eD32
DSuLUjWUUX3xZJ72/Aq2XDErvPyvnSXaa1SK0SUJmmDX1Z1XlIxMy0fAz6X6ct6v7Tt5UCULGC7O
D1mcVnRreRoJeyUG9IlJZsoVWk2K05Ghph5XFcSoQRX+s3Bm7hX+p/rusYRyqrD3qiqMfnkE3S50
47TH8Ft5xDpk6Pp3JcwGjFVny6CUD4JJD27nOBd/VqDghwua6Ct2djwGlmaYaiP6yBwnDeE1uyBr
q0dil1B37U0OsLNaNg+G6Bq+JH2gdJa36gQC17T+RmM76fTc4AlIbfP1o+0+B/VSgGWTVoflHxRU
PbKnfIuEaCO1f8P24py4GWM/Fh9qKHgLsc0OxXNDVzuC4nnof7oaNfmHgGf0xbRtvW25pQ6Q548T
fqztMdhWMqUTRt6jrhS+7ct0CBscXRm/WzvQ1l9LvyA67ZhEsD5OxJSGSEFtHzOFQ+H+ChyC7YNu
064iuZ6X4m81+KCctbPOlBSzdcxud+k0Y9g8Tr9eE2WFS64KBXxlxG+xlQ8tKVIvzdb8huu++kmq
v6lt6lEptADtNA5I3FKrj/F7fgaNBeBFeui4V2NgMycFPIcepZvEfJkJ3JE2gGPrc7xdbVf6bqb+
I+r4UtQkLo/quu4KtXeMA8MsVviYv9Z7T+3FFx2qW8dczqf3B05crUrM8JBXoltg/eUb1RykYDj3
STl+YWRTr1oOTBK9RdyFFHFABz5dYjO9bJSvx87bUewoHPVO+VurkVlam6k/wyBOPI77S+BGEtcm
C3NhxJPB+lMy0yiUPBLYDxeEQjXbL/A8qwPPUwmULEgyl92+O3zm2PDIGce0WGA0rLN11HuNbCkJ
uASEdnKu5UsPFl3hdZ1JLU1rPqses3zAJxf7tFQ80gTc2kSO3+It4DKZWpvmo7+MH2CddbJrHguv
iGFgIsRns4f9eqzCX6N/nTyCkrF8YQOdu0xd5qgNM+yjxcIovzX+sKxpkeAyeUNrlV9B3WAOlSOf
h0U4V0eyePW7ohzXUCQvah2fRQysgTNeX5KhiFNU4wSA76nmBWkAJm9L32fCG881ByCZoK/2eMVb
1YcH4/BxKLEob70Vq5tRwn5VZdWLEcDMg4Wky9/9yG+5n7BOG7cyfmu6DOAglZL7HpWcjqIqs2ue
pN4KUmCZ/IiYYesYgakRCKAXP636gelieD1I1XdJ1hDYUI2QX1zlXBKIDYXCFlSnx54+AKwNkQhi
DNpzzbO8HYHY253ev0ZKFI/rKy1FnpmsQNW7cRMu+XI+TfbHAs7418Rqn9BwNGPeYuTvGQ6s1g4M
0HVsFkrDG+EjBYxUportdRez6w9U7uN0RWIQOacIcg3gvprCkLPs8dQSHs0LbL52ZVw3jiACaS3B
AwyTMgiW3vt/oCeNIde/yMhXJ2CJUH6FlxKf+5iKNe8AK6lq/0fylDiS0DFJSX57apJuMQVEp5v1
H65iFL5cGw6Pf75qiIRRzT/PKhP5FGRdL7NbiFf3ewx/LTew2+SaJPFBcuXt57c7hW2l9fziHBLo
8Yv8ZPsmNZz9O6C44Abq1dtKWEH42h5CYWgewKupiCDgQULorQFlXAglGGgjT8bQUel7Cjfn2cfR
PVoygR/7fLDyRApL1wtriyNG6FONyLwwiJbhfEO4f7y5E4r/daeJIyx352BN1OiBBSoabAZRR+3p
2Btxc4ihsPRKxLueCEAfYCnm5MxhfN8Ha+L5/XVmhbAi3NPs+lIf6C1+KdaVQwNb2VbJA6JlYJ6N
AMa88g5cok3d4nk7GbgZjs87HT/gRr66e/Hit54cFBg/rfHWPpN0TIaKQQiEZNiTw8/XY0FnvFZY
NXkdqHW2tFjkpyD041OSK55bkw1Pfiqm+CGauJac10h81fvoBcx2ni4oEnc1CKuwNY+qQGcW8x6C
c3c3rPcFO6dr7la3VMKB6qsk/0s65Spq21wm1PHseic1J27lJ3A5p+4UzwiGSuKdkjKtyHq5Qv3J
FKwDYMY9gDtVciwyOCRhuSfw4FKLhBmN5kdqJKxk23j5OwEBXg6QB3oIX99jckBH1RQ0D3L/zNEN
yVMai7ZxZ4LOugBUMGNmVplDvKG/slZjPUOqNUrKj70sC8RAarBHPmyCaLjExgmmMp6IHjgn+PB5
+fDiIzvz7ov0ZLTbeGHVnvY329SfoSCBq3T4vW/nFkBfhMh5eI0cc+u70btJ0S+2dGHc4G0EsyMc
IhH0/OJj1jJg8GBgvPw+pj0f5FZKGIgAjBbC5tTxOU37YKhkcLp5t1FisMSqoOtUrV3Kj7+uJGz1
T2QrirHeDMV5eb8F96sjUKfekdZdp3oU/n9FbdrDNn9Gw1u4vLDrmrtxBKWeR1KBIytdDF/LPhnT
SFIdqxHjpan4+N7qoWFVUtI03Wez8uXvcfIBgkRuOn2KrVci+R2o0RTKEJGa2S/jftrTJgh+GHag
xWT2sKja76SJJpfb3UPeLIbrPFsnH1ouUr/Mwl4UqAn25oPhGU7xi+ZDKIjnSP9oS+R1/NOO1UMR
3pln2lPFNKnxHN+QU9ZZOZV/Li9oSbaMzVTiyd/JNZLTRrv6nP3NvDNQppimtdkZkzChhOPZZZCM
7R6As1QbIzCaj3XdGlrtoNRSrg0hWZqDNay50LOiFrb/dPjR740qXU2J/5+g3kd2wVyYHP5PYso/
E3VqjJRGKhs54xmppdTt9FkqxSsVjPUn4iU7CuK7YBEhmlgFSBmhJ1Lis74zitSPNzyScFZcsXFm
bCuzLjRxtS/71/40R9rrHrZjOvx53480PCsnhV7t9v5bUBCZnO34bhNF+eXFVYrg1ugLh2l+gGmt
57UbWy8DDRMDshsqtmvNW9aaMjjZ02+eop22zCfnY+fdqTbb1YLeo1i+F69jWClEw4XtPVUmBHO3
hc/xpLOgEjQWOBABjBl2S2CaWExQOj8+B1cDpcJ5HkW02rNDkjuIe803ZA/OWuXA5F9dj+CmbT9l
MuO1xQE5bV3fgnnshPi0aVDeYI2pXSrKsL377ADR48sS4l03i5ITiFe5biz8UxWwyAh/KgNfGewn
IRrrlhql0XfSxP9fEHZkqCu9R13FcY4V75vtLFk4cFMGo7WTDJTgNaVz20PZWFkDvrTHodtrhn5t
52RvGH3xrkCcuqegQYvcxkGF2FlDgGsWLA2shOROEK27D+K5/6wh0/7BRTKQEUTvkuCTocCYSSjm
lW5pur/L63jXCnhyMPLIorkfNWYEQeiHAfrFKKszlk3S2H3fWuljspu0sI6CQ5lQIJwZp/HQwppp
reG0FsKL8VGLPievDD4tx97qT7L55SWvAaW8EbKi6jLwLSnlMMO5WZ3D1r5///grF5pFs9xuxk6S
3J1pCgSoDpRYTRTgSSm2D6qU5RAXmkDrgvJ8jTd8IOkO2tuc3ew3hTj2CsfWd+qlt5OM7kWRiTpY
QiFHAGI+697f901Znw26C12nzCS1EBYCcAtUSGtCqAxbqJ0Jp5w1WXPqHEuHqcm9qW5sfYqRiMPt
ZyCqq1HdrAx67jCD6aIemZpBSkjC23lYuewElUtc995Y/gR8C2eX21Ri2d+nWvnOw5e+UMgNWmaV
RamNEOfP22vIl3fJEl9LRobUDiMN1Rof427JppZuuOutqD5PV8Ztme3NNzOyrKf+mlWyA+aiu6CK
1jCWnAKQ7ICVt0f49iargaTmCvnwUVDPOCdWBy1EnI/QnVpd8+CJyUDJ5HHLXVzvPZ00XuusHZ+J
A/Lspj0cTP6pLJJmIOKZ2oXdC9PBevZURbJXfB/DgL6DN6J3RTpdFWtXD7KYkbZkb1YHrKOzu6by
Tsj9JkfpM1OIhgyEqfpfrqMq1+3g4EPxew4cp2Wl2AB2xKNJqLGg2P3rafb2tTHRZLM+tvUGBPlG
98mee8H64ZnErblgRJ2z3cxS0W7tckQey9WckS0mBShu2unbE2B/GPP7/gtmpddZKxzEugiGrsXQ
/vmfEN+p5/Zr/tMyoN6JTR7zo4+JNGTCMjD1kTBKFVfMKS6748LibCBPGqqDaUVqn3c++rqaQv6h
X/ZhSq9axhgW7f2nzFg2Gqiih5z/Ke45XNhJESf1Y7g9J3cTdrA0tmLZmV7oNKhJUr2gXxUASI4y
0z+ZRue1wZTpKuX/sTbcMmL6jJqbSjnPE0u/qLISJL8UUUTrEBdNtfte0CAOIQ1lt9/fWF7cLTbZ
XTxtjYm5lV4A22lCYF3+wY+CfrUUEcbj35O6RtjDxwDADPHjM7KdcCnUDcWN2ripX7VEXF9irIik
wFkpBNYwXoqHJNZnbkduV/5v3p7mG5PesgaOI5tzSxUXJGEpvIf25CE0Hgc5/KQ9GH7EuweCgSMZ
xWSN022onBj5zR9lUxG+tZG8lpFfECGjvNaw8B6lRGb9RIf0vpNoP60Wm1HKdeH3ODA4byDEyviE
horJD0mxx55b2q7h0OeOlm85DMb+cr3ig2QII3W1W92xw8tlsYtYgyPA4iEbOYSakFRDg8Z6go7t
wZyW6NbmEnK28Te3VQ502cVCg0fTy10RQ5Z4npfm6xFngIC/+4U9UndYiHtEupDTe/WqDc7KQ+C0
ay11AKYXiG9JYgwTFvAlgrcScSKRGmpKPd/K2rZ8j3Nu3DvKTO9q75tpZD7MUCqHq5fMTue1jw/w
MEmH2vy0ar8E9tdX1KpSn5+fwOUwa3ctx3Jm3RgCzknpGAxeG37O4xDF9aOHWylS8ThiPcdF5LLl
fkVkomwQVQbOBoI+LlIbCCiwCIxYLsZL/X9h2XiYDAt6q+HmbeWeM/alIz053bEM2/wj5lRI9udH
ZB/ugpJPTPVJKnD4k+YSMQf0qdPhAD/IRTIXnvrLT+1PQ23M07KHR1RQfTlGxY0gxE2uqifynZdF
tFDgpGscYRHJu+LsGbm/CYgL7cajDfk0tiAf5MCXUDMMGPMWSqLTOQcZZNgL9upEimtnRXQHk8ng
oldVhDQ23sBLzgCgT57obJ76apgKxNHR2/QxTnS46SH922Au03LCzbCSdSfwprydyWNcAV/dZn7G
7/4K7/zOqgyOcbEAy6wQFwhseDlzIq4aDx452IDARrSmpPWDD6eo/I0n7P9qehXqK2F9S0TwGR/X
nx9sc0R39ZSILoP6wt3adxP030fPGWvPC9IhNsCRmOKGXoeBRdeEpq/5n5W/MJ5E3S+d763/eqkg
sJqKl24n/lKHVS4Jy0XhUtxMfv+xcPrWVXUqaudRmtto+qx0hVu/Hc5OZKpltcnczL8toA18GoSU
nZKEBpr7SD4PRFAcjaYu9k76L7eS+3SYteBk9a1UrfPivLLivWi7L5ylSoGbOPxr8K0L3cuUvOvR
uG5QuwAUXrWl5TekhTsyPya5x2dSh60p7XypLkUbN1ypQMQKUYOBWBXoH41ADXb9rb1lcQ+6Wd2z
V13wBMC3UqvxpEWeuwj3V1RXSCL4vfBtFzKrB6+vwFGrKP0BbU04pPhOLRh9M5ilc7thlgpUNekA
b4uyE46l+f6TyQjQegLnsgOxXTFGLkM8Kw+KFCGbE0scww9sR1Kj2HxCieHsbyO1k4NTUG2Nro0r
kCWXKFFurA/hi4r6laOgbfJde9JylQG/0tkeLHu7ZAWXBgUlad/7gl96n8vrt5QxWw75IgwuppLx
T8cDm7rOzOSNC93g78Tb70Rmz5BJGwG9ItXZgEgurRR41n2fdfK8zDaYU/PHX5HHjxrmzFEsxoDY
e297+JDq/Ks0+IJMhR7NsxSK/mOFMzJyRbXH/8uKmQtGOgbLfkbQw/tMEmchZ8gpI1de2O6JQ9a5
AlTNseNPK/nP/DZdTY6aNmC5Pm1c0PnAXbukVncoE33SXApFVBivxowK41fJWyW6IGeVtV6uv7b7
cS5T3R3/yjcAAAiz2Ca5v5p+zUzUtzzhSTeESW18gOkOotyAJODjfbvR6HxnHfRHfOay8VbWXMpc
rRvU26Jd/VdZagKiruwnz/OCgcmyS5aaIWUY2FHP8eW8hzobyIDkCnxRZCEO8bSoCiOw8epf8lbF
X5L6fVr+2RGW1sPtmYZN5elDE8qD9UpLuuMrII1R5tTKbCmTsoKA56q5KJQIQfoowp8rUQhbKbpD
3Nf4vHDNKurcgsEVxYoORgJ8RRgq5TmwwkTYO3rCnaO8TLpeKQ5mXYZQmG+Uso7tZc4FEWphIhfK
CyNG7FmPdfUXh76XMaregtTe3MNtKT5oE248VEocDQbhUHq3eFlPJ8Mo7Yj4tpRW0W/W9P1Kx2lT
DQw++HxOfS9MR0tjqK+17uEJ2fTkXlS14Zs7GJ4mpoSowi6Ouo7kVtX48eOz5TzIhkcsbNCka8DT
osjeFzgD1Dy0gBhADGKifgBWNI8LMmKrhfLJB3CU3Kr4TxtNmG3Q1ZfT15cmGV2S9OASdDcVTEe4
OEue8vUv3d9MYqzbgsq8IHK4P0si8eojWqNhO7yzlFCqLacDcfcvvwTkn2WpxQTiT1H7WbA2kp3x
AC0Tl/4vLdQl+DS85RhHpVlVw56XGOOLU0LRjyBNhWq02qGK3O8F0SG5eP8LHlvvwGSWA1zS2YLS
sV3VkQ7ly3KEXk5BOcvIpchuYK9397dAQlxBnn/kofsr4KNJNG3WvOz7TXr2mZUGCMsSJhF0s2Qz
0EkVIzS0izzkA48kxqok/9XE9zj4BwzX263b4hN9R/mgr9J/IZRBlW0U/mgw/lQD34ys+WLRm2Sr
h0ULWzG+GAQUzKvAtgpNhG6FxsEyOdCcNnG/YzQxh8XtCgTulmdEFHxId+LqzqpfzZvxGRTnf3ot
8VdDLfLa7UoHMIfMX4CyonpWb3FkSqlqLgwrgCmp5ihdAVGTVVwImemhTR3YtzY/bweDbfy7lyIF
ZRunqtVDMaY+8jousX8iIDOBqByZRiFZZVKrs+FYX9cH1unZSEF6j/M8Ug7QKKXA3So5QTTCCm29
sTgsQWjZFztnu3Vhio5h+YfaXdK6/XAgkCA8XrS1tPjZbbd8pvbYX4gzSumDou4oLfx+FNG7U+sP
wpJ668QauX93B1FpbZujEzexqht+DJ4tvxtBQxAoOVJ32HNafZqX6lNehPOarAhH1wVI/Cp0JErx
hNHCW0oxG2BJlT6RaFCCdEA6MThs2k12XnshkrXl7dPufr2EKp5iNf54GjCPT7gByza7qMJNSc4H
57JmwkD+IChXB1OzlFy8mM5dDIMDxl4IVx5wLKze1vAJriXbN97jJVc4aup7Ac0PScyeuC2MeH5n
x3hI0I5jQgLGFP/g0lY3mCyf9HMcw+Vj23gz9I5rMPZduNxv7ag+HPI83Z1iJ9V5/HDx5H8sEGlk
fCF6p5UG8r0prHx66Orwp/qBpXGbw6h5kPKuK1P3gGoZmgbd/agkbfZ0VU8EWtbddpCbTjWOCssa
58abw3C+3UYWQNQFhWxfHFgtAT4s+lgtepmCGZUqkyEAgFt+bloeuLc/l/AHA44r0Ez/0/gFrIeS
+iIieeEV0i4r5RNtO0ga1WTL/GcLzLRDtt/eIrFGnKfKlGyjEh1rFG1Z1Nuu1gVpyOjXupom0q49
y93gWJe2EUbLyS0LDoT1twyRKl9AZ40SKgsVlF0zQxjkGSt7yOisZrIQvivS9DzzxsLOeTuiu5Km
m5RLXZWAycS0RhkKKe6XsDJMq0V1pD4swII5r+ETUvHLbDa355wSX2nL6TB9Bq/d/yi4ndsfL2/S
ffBLGqO1uOVEQTxku+D+0FlX7GV+wIy7ughw4AddDcOxWCG7D8Q+dPnfqZ4t2upKafxUoAeEEgBK
UJKH6mndq09wwyX6rhXlWun35KixDYzDdn3eh/EHf+zu8gyEsqgBAHP2bjbuBvDPMjX9R4gNfanP
J2ccjG6Cr02VlGK7NGqlyPd/7F8DiYwGZMrwG6gkPtxEwExXJlpRy7IVKeOLftOrnjLZCHV40u4V
7IRwFcMz8pFPzzshcXYKlMEnxfSAzFpYFW9pmx4GgwG8GARqerbqvU0klAxTjCGDVG8O9eKm0WBc
s+mwtBGA5xFWdHy8OJRvp7jn9q/j6WtCqbCDxtUeaajx/7jxBha9p1Ftw8k8xtrG5mweD8+LFmv1
HY56lH8B0QWqAPCLlYaDdncqr0ovxDJAFRPLwCdRrKTJRU8pOH5LCrT2MD+0jtcG8iFgRwDHLBjY
HtqBg1jiqMu36R4T434tJzyyfug0yg/TmceQpJpTqrIht0FBI42Vv0mTrKjD1AWJnnE5Uy1rs8St
uGc7glpND9AmuqYkjEe4XKTHVpb8YN+VMaucMGpvBgM7U7ygyWJjoyv+TxGoe4HHHnjz5wr5ZxyM
qJiHLeDZhnX2tv6+o+osN50Sn8eR6n3RLHQOoDizmGRsMhjHqx7ZlS05s3NWoXPuCsjrPqEivfDf
2VLCvxhbpL3+eHKZyeZzwX8dPk8OOxTWPbrM5dbx0Axvs2VyzOWRixQGkCGIxlhqdq8kF5TbBDaR
Ok/zhowTKRnYmY30Z96Pmzd1KnygHjOfjd0in/92UGcNGL73EcCpoEJTYe0zFNONzxpq3E2txXPI
lt4vBtKAZO4nFFXO2bXOikFAht0WTN30bp/k5t20YupdzMQJyK2P9b2VjvrJltJWqj94b+/5KPyu
15c41qGNykls7I5pDiUqIt9wjU3dRYx3NzI0lSnAnuxQ4m1JYr1lt5CoN+izvuWYSvurRsONLF6Z
NJUb1+kRfQxXGuPeWM11Zr9LKj/qynxPtzAh9cCzKhUCxKUEZlFxVN1nE9E93ltqZPfsnp1qZVIx
okfXgd6s2cQL6eiXPJ3wS7hyqpPYe/eEitoPyl1LwBCgwNQhPxaN8cpoT17dWa8cMKbxv9foYfk9
Dw4wKY32OqRkTIvEBPePnlZrFWwPPoMm64526ze1dXZ6wAV0IAmCzAOCFSkl6K+zOfbD+x6K8jHf
LGJ+sVPLJNASyr2q+0+TJf0dkHgzu5an90ABscpKEGkTonbDkaH2OoipCM8nJUv8JHU9WPsmW9Cb
F1VNgPd3y2kGr5bidtig6BPXCixd6aVF17AShaXVVjwKKswsNycB2KOOguFqE+EvIN+OzdM/Z4OL
N8YAiAd8jkM6/DbnvsU2Hfc14abhwjMpWY7LyrqhloSCa1vBr6kJrFrj2QA2uT1N6mrs8lywv8+j
XURRWaJs4Pg2ZrgceqRSLAtccbRlhRsjLu425On2yAsZHo80D7dWbISngdbXM0FJDPgsHFS2YuwN
pUr+34WIVuVhjCw+LJm1Fx9mgQisIblpvuUJ/V0MqzToG4tnObpZrIrNFCKP+4k2J1ITrhxv1rGc
PioGc0YHQI0CuyS7tbnfMhYtDMtIZzi6h4gr2T7KDjEBhCEM05GObX/PQLBR2VAXZBjbliXY0qwJ
njy46/QYYnUmKWnbMutw7VBCWIw/AGyuS9g+LEqrjdfBzJHakmz2VotinjJYF+u4Cn1Ug6vz2kYa
FVXN5E2KjCXfdhxyYj9ZYrjmSYuBbOlWY/y01Xior9+9CtbgHiVlO65cj75qyminjgFe+QAiRSmy
FdsGhzd3uqudeRWApVrygcpErIbe0HcISHG0e1cUM/lxWHgZybuMszBTA7sUJ5yjlcTEH9PgXo4u
l7YjGX/556yCPbJmS4XnKxmH+IqPs48WvJQUDWr6ch+ur0Ty+5NJjrTd+JigRntYvZoWkPohVNsA
qHehXGiDopXf501jaOwGwFvhfJxx06BWE2BPPIddHZ+jnwKPnGc7Fo1nZ3Slc62ra2SmoaZ7gcYJ
qhYnR+E3sYjUemwoNVYokVkJBQqV4NBakX7NneFDquIms/tMiIzY6kZ2GaHzo4Ra2rpCM/9mvL4o
OT1dt9ecObWA+nZl4NgEGlCoxQZ7yxTjH72o/5YNcZ0M+e1eDS59gR8TYeY7lxPBjZilLwNdLwUC
pe6l7uODvKOU1cMsUOoCuTHaReN64dpCnNG/sGhLP//dI/YHap8HrO4RnSkz5eLB+zQXHQpCKFTu
VQtCG5M/2RX3+UR5HafcJYY4OG6d1a/YICpBAbVBx9xi0SXZXFwJMoFBt1OpZMq7+9H6IWWxldF8
wHHgYNMopap5DQZnIY7Z8IsAg11ppxFDAsozZhjavVigHzvTk4uuK27HxE0cYH3LXNHJczbZdXSt
p3kHKznuDzXnWGmw1Le3v8Crs0GU8FPTh8GbziNwiqBCMclHrUXthQGbHtTL9ajc9m0SzA7TC0Oq
IVgkdO0SnBdmb78KYlOIuAsamvMjDwQGAvyuetbLk3pFrCCUGdiX1RGE91o5N0vs4QOcu3RJsbaM
EaySxf6LSMHq57EKgoLhUS5Hker9Z+FDnDCqE7LnhxAadkfHWgpMwFYv4AFqBZQBxBt9sZS4WlOH
0LsSA711MLIes7IVi1ddTnI2wO1p0fuUD2u5giG0/XTiZ/annrCaHUtfsjQ/nsjbf0vMeeD7x4D0
wPL48nB+XK/RrP3bQFFd6oC+iBvgkDvTLzx01hculhBGDG0tivBU9mjGtswlD3ES+/tl6WD1GHxq
9pfb+zu7CEULt4+8axMICD795MhkB+7Y3og6KvT4bKB+x0i1WGW6WCc+GOQufXXtFkQIixH6zDRC
ExWhC2Ao23IRav9UOuQdMQB8DOmmEUi5Chi5PwiHfDJ0shT1P/U/dpEBjxlrnzNG0PMDjJ9TMG9d
TnSW1SxO2nq8AxWX4dGjhl/nl2umILT4WwFDOuD/Np8wh4P92j4O+ff6OV0fAy36l1q9fUZDdHA/
D1kUzVgQ+7f3sSlTvMMczjVgGCD7MwMAu6xupThOhzzPQzyqOup0Kiyn3esoSJgC2DPro6v5J9K0
TZqjdPm0eH8LP6Ume2YDA9I4lwdK0UQEZS4fz++4MupVJCNiO1YroF03jAd0YfNSecUkFwoVrPV/
12nvkYK28gI5qqqhLTcxasfT4P8BkLzbsDq8SzpIxUiVFXHVMXPe3MHvpS4nQMwJPuaDC3BfeZhT
S12UqjJ+Vr9ho41n8EjisbDRYdf3Jp/dv792p/QYG3r753NROwm11xSFpH0iJKPg+dhNcu5CO0Am
Hz3gqwE0eH1v1C5bP0FJSu9/KvvWvy2S+Z7G3K2TYyVgd/Yr8/iuTBjDU1sI4Jczuv76xTL9RQ4O
WoitpNHuOw3VvYbTSurttGi//OHnHreL/E15bUtYnJPn4s8Wxh0yuVWP1P9EVVyDizar+zhnQ0Iz
w03RKsi/VJ18ZgKPMSPij10vFSApO5XN/J9C1Rn6wCj6fCbsCUdVuhLRUOEE2t8zLz1Pw1sqcH57
gj8WvC0W+q6wGzJZNmD0E855vFRkGqntU9Pxh09GRnZ9MjMZqCchTVyWJX1387eKBIe/8OLQiH7y
DW2TJnd8wjQ00BsXyopnntUSi9CGbbHwsFrC+9NZ06vcBqrN/7HnQCopI6t1rQDY0vVVw72l3WpY
3YPmHmZ8O6OXoGbaHTtGNyYuDqGbDnyFFhy3QjcBMHpHlLcpW2UosefZnVley4FQFMO3v5iJX/Vc
hMGWExIQ3pikcph2R/1DBfXiu1Ri8gFmDk7de2UyupMGHjWopkcsWRncpeNIawabXhbkJN4WQB+r
ENm1LDuCqa5GFMiuLtKq5OGXfwI/tf8Fc8AoTL/2dhJ7sN6xMWjt6iGxeGjBYm9hF0WNUTvvHe8t
28rUwXIf+Dy27KlyGYcJgOasXfGft4J70UjFSzAxtmvK/jLZFyFvee9MHHcft4beBDTXUufy84iS
QdiHBoFZo26kpryIWX3EeCVKNd08Rqhvoq8QVXg/AxHosmuyPlmNQqd9Qvw+ACBkf1JvDCXznai+
OeanFRW4JB/zr00pgGLvOHeZJyAdBgiPyoSgZSl3RjDD0x8bgl5ijKRYCHwIwAnxQTz379iqhZdP
kLtmI8UgiXKp07yu2x6398AIm2sTaHj+JkQSUPt0OXMxnk0o5J0Ao5Nuwd3BXMuKFKyRY7hNeXub
tB/6+XzNlzp0pIFtCmcHOxalYW1NsPJlXv/OvIaeo9o3/PUEFQ81V4xxlWy6Y6BeCX+i0HWkBFrL
NG3G7LQRGuOFqYAGLS6/SZnbm2VmQKYBaiv88Dr+zE6Ex8D97NC1gIerCyPP/mo+2rwt/mQaK4rZ
ZtTl82b1GfsSCmu3AbtXYqIbCrWvv3mCL5EQxWriaQCk1Y8QSi8EoXhkhTrAxSxWrhn8Vuj283VU
6nA3P17jCVvrsVk5Hjgovy8V8+5b/7JJMz7PdTDnyu77kD39wYxVWCbpqWc98JS2q6PeehDiM3XW
dV5OxF1+xmlnp7zqRT01WfRoiOUrhEHSM6c0nXL1s7Fu6AB/JVrIMaiLLWiexo7G8DV4Hf2R6BZJ
Y5YkOglB/n6TiWwQIr/l/Pj8UuMy4yesTvDoz5w5VJXvZj9GPc/q8fbrHbV2+HFao8lQCvFgOQsM
qEYM5nvfPEAUjSos/aplwX8wSzJHGyCMASBfQtiW6scZOp3jNW2LeP5Wm67EIR3ESG7RSWPTStUq
wj0cf7rgHNUkxWbK77H8JYD2Va0Oj9qcyn0aONPnjf4xZ3KAlBrvz4owP1PNALjm5GSI6euikk4p
7I37N9tMkWQwv4BkAo209NfMu3mZgnUUmJrkvJh0zzBxUWW+j18XIAP3Z/BXJdUlYXUaSarYPSrR
0VcPlLhrHZNafUGlrB6d+9GiO7TZKKsOmoxh9fXW5oQI1DrhPGFFctWLsHmvlx3AuhHKseMFB/72
3ykSSKQTahPnfp+7jXZvGlPALPCgl7YzC+Pm7461zUwkn+trFo88QrFGYqIi16XS9whuvynUSQ62
P8oTwslgifupQtisF8qvKkpgDqXOLSpq5AGioT7wWDd0hLOK3fbdieFkZJvL/Fl9EBhbBrf+AvNi
fMbR7xyo8p2L3Fl2Y2qz4CoeXfsBHX4LZHeBdzJApioR3KmFgRUMeadZIQWl0mf0AZPtLpnFqJLu
HJ+eLexSDkvFnSI9Y6jFaVilX1ahw4vKk50cAyTdzSwvM6220V6Q4/YrKTa0SIbpGnDt4vqKoZwa
gbMw7xBV0nW6jIGJHXMys2wd0bQUZ1fJnSbVcBL0EozttPQHtgJxDUsA/iqqMq4XclibeRUoGppu
Os9i5VgivPb8ll6EyEoJpvNJcjGXCprQm7WRlbJRNYaM1i/+M/B3fXT0WFob0/SGzNHQbeftEg9W
WI2jAqCGNHiAP+kO3ymPLRn7BshBGESeO6KX/CU82igMcy1TP/Xj/MFzuVDOLrTyrR5hLIw6wuCN
vaF7UYhjqE0GibiSwX7Acq663YbEWxLWppxBtlFF+ot+K9LEUL2XgVv4aaQU/N1C4s1NwB3H3P+H
M447D81A0xIcQSA5wTomFWTqC+DDEPT0Qm3Yk3U74IQjh/5hJqwQUiFlDST3BPh9v7usI3UfcJQY
8Rd8tDgo7qSoft+5NXU+AO61GQK6p7zKOX6aguN/EGVMwoX+SSeljoM7u4Ha+IT1ZdP7zAGcUp1W
MJK57pzkNqZygOeULypuLQbovVdOh31EEw9oW/CovpBwhtS9owVQfmJMQ5Xnsm3rcS9yv5tZd/d4
eQg1q0OX6GLQTN9+n6RHPgZ6VJBpmzf6la4VI/bzqYvMnmRQLa8vSxlvFoOx1ZfnISAC/ZyuiUXD
Xelmt8XtaVx8HXe89OMeq4n4LZ6zxQ9D6bDLer15FjTwgjtXG/2QbxDVn6MYY0ijSbriEd8Bhlbv
tZVVjZ0BPyxfJwYA2SScWV5fyohSI1OoCdLdodQC7J6NWMbTTkk8babBQShPgyFXsu6UUTEr4fWE
WfJuqU+miuu6NNjacdWDMHcjYOhmb+7CMo70QB9Rxpje9d5hpD0yGXGiaTj3cX16g+GVShXhsAnB
ZfMAXFDvA1nOt54N6g0s/qNIHMe0ZJ+f4JSi0A7DSmTfj3CUg55a9ao74sdgFbbhnYCnGnBaZpCx
iBchM2d9yLNyD/ExXcO7JL35Wq7QcqNsYED0dWsmDrfmJMOGXa2F2NCcVePhcbm6N1e3iWwLM7n+
Jjqqn80IJQHNfj8QHAZBriIqTtzpCcJB0xWM7Gz0X9suICuyjNNITq2O+3C48O9DwEjEONwHkvwq
I7INbL53LmeK14UThMHDIKIkY/7U4DZvufb3Fu86fcjd1M+nDGKxib4/gqpWRkmDBkFwg7e6QYeZ
6qT0BzpgjTr/H44KqDqIKWw2d3MgsID+sE06Cgg1E2riMnLpr8aeMLxhmgsehxmhICiMPOJLAY6G
cSYPqgJryuuO8qROGYgLCfm7sZMnhW3HEzIqW7NjmEMOyIm5+6XdXcMVlyQvlvfSZz+rZwoD0cjk
4n9yw4zx9cBpkml28Fg8pjaqLa3LFfg/OBTaAvebEBQKOM7o43n+u4ObZbATnSENiWmXbSa57bHT
Z4cUBBLAt8LK3LgUT8o3Gq1+32RQjw1poZwKxjcpZQLLne2NoOrj7/YAUgH5noLvAhrHb87iUbLE
emcSNddj9373RrzaEt9Ebs9f/y37XCkAFtIG/++65kL8tJrOhClnq/hJG0/a3AIGRyo1IAWlYjz7
mnBrQ851Jwznp6n1+Iba9zf5FJ3+pqtohXVcwpQ+mB9UHfSNogUVSJlpUVzBWKHL+geKUQZ3TUAa
Bay4JNfgJ98JENmwdQOt+IXF0uUaK6RNzYk4OwOjub9bgJbA5fr4TtE0zeUU6EoaKxq7+d7Yq0BP
PjojbwMfpjYFJESmzyiOIEw2aH/FwlMcCyenZjBmXKiakpSZEcm9yNk+WzOOhWExGc8x+SQh8Qsu
uJUUpfb8mbyVt4hfFPA5E2Gozu+a88P2DuVlNQbVKUp2laEW+9CsN0x5WXuQL7rYzyS7FsFT+e8x
Ro3f9gXVA9VdGCdTLEg4bh35tINT9EqUMYceTv7NM0QIS4Q1FVCKc34Ny6ZJaK3PbRLhl7uo8JiQ
im49cs0+XV29iO8UBVkZ1M0kFQu90hxbSLSnJ74VKCsxmNbTLYn+5UD2xs8hr3f3AYMWS9KtUGq6
/tcjco+/2bEa4jj5c4tTxuJJzuS9gB37qCaxQYZVbpL3n3QGwKShrNwfAGJsZqqcxC/3wxqzH37L
71NTJmaorpNdrgwMkk2T3cGMeVyawu2d8ubVuV5ZNI1ue0bpEoddl60rjVLni7iXNTfq79s3mDXu
B63EBH1tsF2e+4SQozwJlH57vhB03qOlHBN9VKFyIYFTMKzfoeYHokfSLc7EIMEr70XMwdq2FBFK
Z5cqnjcEqJyB6FWUp/PgwWFpMTFkl1gVMiYt7F/rBc4Vc4QU2vnVi12AhclYkis3iNwwc2vYkVKb
fU5oGtWI3GSHMtU6ZNB4F7te1BoEhXzRtW8VUURiH5//vdLU2IOMNbuOwtYYzJDAfe3WdzeE6IS0
l+T0fxbKJvuxtFiIMGv/fOhjrlNcFR2QJqNNjNg3K6MdggulhnzFcoeaZC8ZqUmlluFlDumXIOYw
lFnHrNmZXjxTcnXLpGdi2EPfnB7RuALV/UNz9kOfD0Z2LW5MRpbPwJ7RMp6wu3Zskz3S0QZEdIPG
JcxRxg+2EMEm2Pk2HQJGEoBVPAso9ku/zKCRhey3TfGRDJGGilCuCCtNhU4pOW319PgNpAhI0eR2
WsvhmOfbGgcs2ymRlU0jbjiFSOKZkByQ4OiOHqodoWWnkI1PD4oo1qB3n85kQZQOSOinodsTgF1r
GTkFo5MnBtXPRMruNny4GYPeG18RoX9ZjzyIULZffRY6eTMVes7aGnwLTcgt8V4kZfpAOqnKaSDP
6MjN9qsSo4Nr8R4fMHqpB0+3eeb7vLD2hUj2OJVEzucPfdXBMHsZTUhxhkV4tYxVPnNtNADmuETb
sdHY9E0LKPCyhv8xlGhasoXY4MqHegH8Hc40VTxrujGMz0drPgqbTKy2NRibFZyRJON870ugFYrC
aAORXsq1ODdk949zcN2ex5TT6PEPTXcb3C97x9kjZ2TttxGsK1SyJ60F+ObFgOs0q3L9k02TPOQV
wWXrwf9e4CIuSUPofqMs5J29E5EtU5vmaBAYue4aFPbJxN78Z87sed+fm45lL4+GUCjJ+tszs5Zh
gJicHpYJJ02qVgm8S5+/UFmkNG3VmAJF8oXnsJp7T0ularYyDRmqL9UlT2f4CHZR+yIzoE/syXRq
nr4svUNkGRUX2HVlqfdfBAcH2U6nh1R8y7CSAlqINKlxO2rJbxiFVdcs3KN/b7H/R7cxfPKVbND5
aeKh40q4LlaM7Qday1/U89Ws85xpaF3RnBslGWMiZ3vXDX5ABA1DMEsRf5ZpdjXmF8481ricce6D
ae/1h0Hb2+bH8Rk7u0pcwysV1DZ6qywAe5SMyr38cTUn19tzKSmoGeDm4j0FkdkaepP/89ZxGTCg
5TmvJTA8V1Ap9zEn8EtS03osEvN0QZjSYNLyJacbT2TP61gn3NKUIm6jFmScNCTfDHwAjNZDxuV0
0TuXVUTv1q49nCeuLcnFyzT4DhWJLmBfRiahbMLY+EttNdTVgq3QGuCb+rhZiFGkeblqIOobL/E0
PH/pRYYPcq5Zta+hYedfTwHIErbXYO1M/fDMk8dFTtzG2VK5XETEGbArr8wKEm4XVHgB5AH2wSu+
pzba034bgeeRP9ffWOt7iNQW8rKO+9YS1KBfeQgwVTWf/4a6EUZe2SQXAQ+VESQjQ0XmfAa9NX8W
qsCtCNlzYk5ekIxz5wUbnurlSFY9XndZdOEwSfxf5PTxHUc2qUUuTyhM0pdG+iiVvbZuA04ZjHhV
pnLycpHas8Lh+cqduvKwQ//Il4AyognFj/udW0mcZOy1v+lnqlypXd2OrwyuOTovgYy98IFs8aZW
sPo9U6wO9ue6Anr8czBjWNqcW7dHmiFuauDP8U/T/+SydOAFUxg3FDCYt08mgIWNHZ5soth3gJBB
b7ZerQExeWvHJcWDGbhxC6sX7OCmipXfQSXVNS8MwxHz39wITi2xDUB37COE9LrOKiFi+6RrzLXv
7NW/wY0JOWnsEB9cOjZNr+qW0Tw/uaQFOATmUpv7tM8FyYMiw918puA+f+iEzVTpNTI9lEaZrGZc
rzSqF0notIgooLXySfCrqpPck8W0ABBex5r9rRdO13xqV/cyd4xYo9AMkrB7Bx5lmIQpb6CypKNm
8FC0NQkB4AI3lAkv8cT0ZIBPODjbMYFwcl2eGZQhqdIi8wqFtD4cPoB6ImSW+LdGzl/zT5uSj6+H
5gm6UhmLGLe7ML3z24/d/AIcMnWfPMMnwHETZVSX1+5sV4D7ERg5yAfVIwinx8JGt81DSvtC+P55
rC/2DKXCKame7gbAFOw3MiSH/UDPifmVdlk/LGPe/jVokP1XXeZYD2E4n48APhbmlilNV5j2KhJ1
q2VwZTGXZyVpev1KqIbwcmZTcIaRWEL9kYeIJh/a/AJEU8OtP1wWjrjOpKSxEUj2tgVBWUCC3Gas
Cq+tbhUN9ftXwXOzbO9KgYWOF2phlqVWJ9JjZITFrBTvB1kVrCD0zPYjMIB8SZ0L1pZb3GGSUqZV
9M8FgY62GXHk6WzydWDviBjqteUsYmD9FmvM8KSaep4gCCk8khX1J3IzvTPT/H1/bDxCpQZIfW8K
jBG2+OEM71hLtdy/w4F94BzD2WUUqDLL/33aZJ0ic1JUWMlhHg18Sdi6TeoByx6nyClZaBc+DsJ6
27BGQIktAPys6/UOwvq2qgIRO6LCtER+h76UaId1+bBwzXnqpYpEgR9brPHBs/bBOfV9GBqIUsYs
XvRBwadv3G+xjYfPz89N82GAj8IGtY69O5sO1zhMUOg5qWbA5NjMZ383UKTh+UnBythGWZagxbaG
P4QgOQQsi6Ki+fcH9Z5g+7m2LZXplDnhwzsDMzg4SvjIqrkYdMxN92REmOfYsO5NAybf1gMmG+64
cUx/g/wQoktyk1wemn26rTQZmbuvDSRlk66EEQNOag03eItBWCPE6tA6O7jdjux3IJhg8eTDeHLD
psbkn8c0szhkdmUyv4GWE6Nge2CgxLRxYN+gtm3MbL/k15wWQCtTKSsz/atJlcuViMGiiz7/YDD1
0P/oKsi+RNSfx9d1822PvAepY+e8zmcn6SX6FKVQoPQLbJMgKNliE4Zsv3OaYIPPoKll5Lu45ijq
pfC8ChzGM2ur/52xiLeLLstyDUAjjtrVROdU8FcGyJR02FoFXlW5N9XpHrhXQIr/ctfiPTgifkPq
IGftTzPAf45VqGD5r35WHELc85exLkh73qY7i+MfKbDBly29W1+rvVvmXZ4qxJu0fmtyemShvSAM
QQ7WcHVBMo3QB7sD6XXzILtMHFiyKXod7wNpChKRVqvhcbIbkvVRcUCInhmC5QIHjj+bQMrjYuTp
ya7aCmluXDzl7YS3pv/QzXahMdSuqtTvSuXHoZXy2HoiZPc8Q44PlZYqBsrdPoc8uUOrWbwOTtPg
WnbdfaGXHvz1IzS+hBahDxSqj5UXCD74V6sOd9H02W7cIKOlOW2JbyYFKYX8sUN16Y0nIiSxccuZ
tMpKk+R67eQDyJEoh0fkduZjOfPP0fzSzS/kVB9spnez7ytsIKVJ/NwnV27dC8MeTvbFW7jKz2B7
zP/h5iRsDfjviAr/tCgViDBg8OkHyvEt/oblFNhfz4eRvxvHMYIzo5aRIpp5Toa6AVRQsKDq5LdC
1DOC91XL0hZOTC8T0o5DEzUph1zJZy08ijjDaq359s9d+RufNVoenc6RXKS0o5SBWt4ueH+zmEwU
cAeHQ3s9DwxDh2zQ0PjRMdflSBhd+iAuOTsaYb3x+6CVD18qwN/lzyTe6fgMEXXvju8Q8BpDEzBE
mwNqTPdDjD828M9jj6gaRC71lIRCZEXV6Of7aV5LnpNJg77oZ1igxOzNzqPsd3WMn3I/WdExn+Ow
4HKEfwFmWzGrX4L1pv37Vpxw33bo3dpRjF+7TxQCMJoFmxweLsOGhBrUM72xMlQ2sqlYpLtkGGWI
dETKD8wo66heHRRa4KC0ZX6HrRHI0/4Mcwnt02C4S6RhWMktsGAQdOMvsvMw1PYee8UyHz/DUWsz
tcASEqSXNEVd12AUsKLd9rwPy2yBmvxohc/KG0EVOfx4urX70MfEmdDLYkR51ko1FXdJ246XVzhg
A9I32KJF/FRJizvQ6H2KWWYS/Ln+KV4zt6a+5qUONclmWZqIBpVTXT3leYxZJ2mIYsEsovFeM1lB
7RVFQ4hD+lSNA7Wqx+Tp2XcVHJSoG5TkRT5nm82esMFKrt5ZrjxmssK6HiN2pWYz7hF+lEcw7Si0
MOC97NTByhj9qAo4ZDCblQF2/uyX+tHbg4fiFcgkD8u8bdHZXsT//SF5e+y+AD+jMsr4Vd+n6lXp
Iw9Xcpwp+1WfwlSiVgdkLmeQ6qMzJUd9XrmPprW8fnt2okvjOXrhussv3aj/43gtxliU3Zsn74jK
X3VMMMRQuR/S+YFfnyO1IMgFMYLN1ukn4cd+yk75avJDWgR3fUuuP/jZv8p9eDIauG3mNCkJxlVy
vDp9XGuY8jT2dwQg0Vfqv5IWE0744NUIpFNyuI4oc/UjLUS6rMr8AsdOUwiA+yXEEKjtnjcJ4mxE
BVUABTwt0nmdw1x6ePCqvX9ZMfLsv6ova1GWcehT9QcPuFOCbLys7UuEGjz/IpvhdNcFMvwMSSVd
v9TwQdLW4pgWJx9JhUfTCvck30YyHYRmWv4/xQtOG/5FU4klOgUZIp2bC1T4O87kSFrC6zGuL+C8
R9IBQeoPkVXEOMBZ9DkJyMi9M4lV7rl7WeC7QHhZSmQOTtWkZ6PbbJshzT9IRO+ioqlegBMlCGLK
pq8Zl9cvbO/7BjQ674lN9PxOY2uY9+e0NgzDnjun8500t9kBHpQGIDYYuE/UB5USJP8sazV5azOv
U3qkDIYF2p7ZRBcwOcyGLdRveVZgYtGIdCojkHiFAMOHEy6SrY9m3iMpqVVHfpaubfiLC7hMOLz3
EmmsgaO+9Fgyp45Nz3OAaQ40/l5EgykyGmCp1/0zQqxxJPp+e45nZDGMmRD1O9iSYy+2sT2J5Jjj
JpScH4P0ocnwiWE2+oclN0Z5ctEhe+17SQ48pKMo+SaA0/sqkNHLyFe2J7hYKmC2asYcKFJ2D4E0
jrrAUTjxBZZh4eM7Sqi0BY4ObcKhDBQtX3RVsi/iKHz7ORReclwSds3DK5PFaM1NGjeXZdHTUQoZ
0Q52wSOWaYXJcjXVC/yXZYyEIPkT9q4tc9q///PDimsh7aR3Ap8YQXqzcWJL/Tjzwun+AOb3MpPK
xEfW9lDAJjd503P42agzgzX52hzDmV//9aDJK055r/tSGHGisruLUOSqpV02APZO7TFYGTWpk+Wg
ZU9o4DyQJI5btRhWhAw0XFW0mIf2Qo0D9yB+Ds84YP0z0y0KFEt6pldngLAcKsbQ8O/O6rNz51H7
sM9jKjyNPdaIBxb992CtqwXprXDxxmW90MNJlp4eSkxV5Ls4ugC2Hxs7XyEGQi7zIkqXN+LhXVzX
EOPiMWBRSVG42gwEyHpBSZKMVSlkKiNwMXRjyBSZxiG1ucpYpYg2eqXWhEBd//QXFvG71RZHVcoQ
zCJaFG3S+ezv4pCWyHk9+eTci+R978bJa6f20o/iW5N23lJzne9zpXr7y3r4OaW2j398F/7cpgAT
FyjZcyqICr6wmz1wAeBE8POAvyQvwvx/eirKaicYquYkfBYx1UZQDJibMRFkSlfuocLOcrDwjQbC
w25HI9You23kTOx8HJ3AtQXh66EzONqHrhvdP94V/71Z4k71hHz+7QUp+8ygz34hX0eC9Q3sYmDK
HucL8hC8DNv8O45Lg9lGJszoKBl/EcSuSx7INI360svkaZsKWoyKICwVCmZ3Wzg3kpz5NTU3B2ge
F8Xo25WERk1jgfBSp5wAcMtIhtXDkvB708QEaWZaRbQhi37B9tPTebPul48BjTALCARzAk5s/TBE
g6gpaznRyw/Qw59P3WASoN8STHMyzQyninoRumykfVJuzBO6w5WNbCCtT5xreFim9ULRVjvdplrY
nY/qkzp9WmzvfxoQPuobnJjB8H1nXnlhUJmdI9gYDHZyO/3PJwYepGAZkGG6iMj0ehugmN0TUWqG
YsoTFYKgIZhc2VK/ZfWV/xpd5DednlfH08la8IbLeSCisNfNEH7O7YJ6qae8Ew3n6wUKSenb9zI/
PPJYRREZ7Wxgrk5Z16129cazLB2kXb7ExUYKrACaZLYybljaWObKr3h822ibmZjpREa2Fs2dMK1Y
3b6UPiv743WwupaEiALLp/epMWucWBQiA341e0S8Adn4BaaFd6nWNzJdrBmNpfBwItbwlyuhmR6r
+C1W8BLVFWB0Z0FtaL9g8j+3466xlmlyhc0ji5p5Hb5Y/LRZfUAqDZuuVPz4asmSgzWGf0IwlC9O
CUou1n2yWs7wKHKB9g9X6HCLdfnmvELt3dUPSrSelcSO1yG52YXRzQx2WgQMpfVNCz14H8jP9ORd
ajMGEOsQAwQUstV6S68iZaF3Gy4bHWy9BOVvmOpHj92Y+EXCjc0TWIei0eyK8Jb9yJCtgcoJMLXZ
yYVV7GwkbrSQk7yNsp0+RLtU5VgU45hiYP+tiZsbsjGoMS24jDXJY52QcQdSrLe/7WFad6i68C/1
O+wOL11/x35hxxcQHU97tWCpbn8epTOUFnFvebuUm8E8MN3I8k74DqKwk021CgvCR1rXz7Ode2Vw
T4O4BlUOpQ75h9Mlm3cCp80sBGtRIZE/myQWa4aAGH5v/W90v5lSQd35M463tf3LhOvNzQdtzqGl
d8RdRD/iKdWPUWAo+7ylBGVfp1YdgkiopPhCg11W8cwVAx0KCNQvBJs9GgVvj0LwW00YHAcNrw+0
Dxc92YFwJJEfsnMzVBK0mE3t7XiyF+6eXXbZ80N1pVh+aWs5MnUIwOq4PoFCIbkwok8tqp2GrheX
fMkFTYbX8U1ni0NIUIO++kJrx232qJoYdGmnlPGYaIW21UjERfDh9CI+QgMfsTB26NdFxkTXDS+Y
qGCBYPBTMGLlV8m/XpmrmQ+AZBz1O9b4ocQAH4aApbqHRqtdLywtL3KsEk+RYbz7SYwu9yXDMdsC
/qxg7wsMODOr9aedCYzkgC332XWBuo38dKMsEUCWxXVUDeofgc82t11QLfGu0EjwA1wDGCmMGkKg
J0BVpXMAu3htxf4w3eeKx5HfR+hmBDiWvYeGMh9X7ZsaZUJuIKUPBYLiovX0nrYqWOCGcB4iwHEe
CQblyeQ6cXBx8PMCiU10oigx03q9bhQQruvDtEfGazGiCKiR1EiGDpFBF2V7mmGRW6d/EZXDicAy
Qr0+qEV0KbCwP5cNgvkwtFM8V8t4U5ja5mt/LVybT47q/pB7zK+FtY77ip5KzlhLvfVhZRIqxUlr
Zv2Etzk3vs8o1YCIkzATLBLmBB2bNN2t/9wcyI8xe/9fZkFMi8Pa4dQI6fVeAnQY3cXiwWVpsGjf
OCrJ3609288fr4YbKbG4i6SlvqgAtxVKiCLdwApW2w+CEgR+UUEQ9Gkr3IBe3Xe6kfS7c1vkGOBs
dhDLR3n3+oOY4JzE7SWNvXPnj8ajXhAolkJjZRcsFgKR6JiKJdhvNU9X2NBKSTv9dDedsTv/WhwT
/4fOwrbOj/qd6gq9tKWwUGztS57kUBJDi1pXwog1PFcpIRgs4Y8++jku/YcmTgTq5Kmjtt+iiHbf
DC3MzjeIOr7jQKY3XuzJ+KJictlIWRj5wswjIv4vAoDjxfE2f/r7jG9Tv61WSqltmw4qZX+2USW/
EoyO5bdi07r4WUN2bNdi5TO87NS9QStjBm9F37r1AxfpJ2V1uQkzIi6QFa7BCCIkhZL3xITIpADK
EtGOXkSIU8Z/mZyvRifRSSmx4cX61zX986Irm6mGiycyfxHUC8+4Ln2XgTpGELiOcuXiMnEY5663
XrDHZcCWDNH6fvWaTs0TFypnMoxGqjmSTv/auUN16tlY4iE7eGjNVj0BzTLM4MY5dzrO4cRN0uvB
8a0mwAiOhDDvUuHsUV0EATyP+Rx0vXuhKSdpyFzZwNktJamVmKT0ppNTOFNmC7d41V6LgunC9kSU
2anoqXPkefa67dCUkrOQoCxTqniPTlHTsMJxYRyBwhf9Ed2dcL43AZHohfreLzlTLLLvrb7QcD3H
QW2UtgabZvy6eZctsMkhgfnZCBaWcVSM7fop6E0pGIo1kknWeZT2ZNloal8XuNs/IIegMgb+TN08
kh957ujlhEiigNn7noqEOzeEkKbUtkNnNqRN2xdVXBJ2oBHLI1TpqyKbN36/ExSgOQwB/UyjEZ5C
upJGe9Y+kK1BC1szW969AbYK7CN2Si5Wq6HpLZcj6FOACUviXNZdwrqlRN+1jK/+z/BZXlYZcCgN
CxdUwsozWO6IO1MxtXGphh7bLmGF31jNixrXzXdGOqnaHitlV1Th9XjQffGcmYny9aUmfTAv48kJ
i1I0Tn00pVjPYxWbbFg0GJIuvOfm0dg3/5LSf6bRYJcrkepm+86QP399dp98gCmYVK2ilYOs973r
pdzCnPPFu53q3+5306r6QSUeTWfzMjaTCAA2YJgCa0iYkF4RwupkSVvoxec4p+omch3Mg0POUUkz
obab4EI9eS6atK2pPx0vGJAkT3Feest3z+mKEf1jKyHPH5YPbFZ852T5P1M889ZkK97xbi64dsJ3
g/nE8JclIGs3aygur7rQzRi/kTCR4H7+3duW4dArapYwLErtMFXl03qkV/SCwMUEu2tHWHCRUarQ
4YG+SQ0Iq6Nqekz+LIllS3fsChuUg2I0CNI6tKEGAjMAdLLPYS+CPLOypLj+QUbPqFGStNETiBKg
WAgoVRczhzYCI+xeXKQg7Ks39Y1f81xqdVMr/GVq8wqm84OwW5hDvV9BzV53QX6zjBRrzFelEXRy
vA6O4TfUdGBqQ7MO+Y607P2i1GSm3n++2yMFU/uedJBF5T2Ia7HhZashK3/ne3V93L8RI4fJ4sJh
YWQU9+LJBGuPmm8Ja+u8rWRh25hhAqbRi32KuzSSkRCFihS05q9iNNSJGhdurppagtt0FhpBZCYn
ZpA44Y16EjT1eNqSenxfJpFb+Joy1twu93RW1zQ3x0i+Z7QdeeTC482xTTwmr/XuNzadZBJfDB1a
wJHZb3TP+/kF/vJ2UqcTePwtdzGVMgNSLm7ARz7vOxYVyzrbFXPKGGqw+4CF2cqLvCme8NgtRMYB
CeekcQn7cN5GS2aS9m3E3lUEve6Y1IhT6JFO2CxGoUDY3jaNfqgUW6bhFcyGuErHXP1PFb7CyqSk
KCay8YO+3hGvr+VIS7RX/668FgiVAc9htWuLR/OXQuA8wt5QvCEK/1n0RLMFfCDUCWUE+nOXzHA+
RMbTsnH9XdtnheeiQMVPE+oo1MEk7IdgyRJZribzrDeWgGZNWcJgYsrNUj6Hdjb9wUwMF529olCB
1CJUkx8alriYD4XtIYcDIKROuYHjySkdB+lTiPdhDKPcDN4ITF00sFamfgshHENG4HU4xKvP+IB3
dD7Oi13R8v789zGngbOlTTEajtQfydOX7E+MmoCNjp9mqqgAP/aCRBjvKUlM8nc2NTJhghDbVyno
bFc2uYwWHc8ZsPxqRtbnhtE35XASg98AyHC4/IJ0WXRILxoc+GA3n17L68ot5xlrw/SLuAEl7Fcu
wAtvM+pC2w2TNjgCpFIzWsmBTioNZv0Y+Ix+zR88k1eNPnY/i9rIU1oK5lkrwJOtuOhmn3GSfUYz
GWwJILjHJH1AT+mbmzWRkDGmJhFbsKVVrwRBP3stF+5/+hVvVbhdKA/acq7GmGTXi9/o7ExcqOrP
8wLgtRpAmkL0G7xlZ1fBFeU4Uo6R2IA3VBfY33MarpXuOR1nJu1PsUBp9iu8peZlSyrFNLlQA3TD
S0VPl5SrtqDETfMWmsoJdkrzpP5A4W/D81kTf30t7hF+V5OdtYN3NvnoF/PNcWNHBgRgAwuL7Y0e
vkJxfxhXBG049S5Kn292lXQ7vSVPQbjAOMUCWFdhmRGiW9AnSTsetx0KAj3hY7WHbwnbsEFDMZLe
fUQ/gQcTYnfiEoSyn+RpULXZFDp163Mw/42mKwnHqL3gB++uvbuIkF0Wj7JFKBsSQHfi84l6Jxtj
tST1W48ucgQSLv+e/5yIJLLrr9k1py8vDezddGrS7KzNoHWPiWHI7MM+uEspkkFJlyShAuepNuee
G+esGib96UlPNFUJDLJhk9pC5b0eEa/f2RpsPw8WNUQP40jqz6kPM/RVnLCrofebQR5B5KYI2SDG
lYCSW5RitjSYBkaNpxB86s4aZYqlVbfs6vHYLILGVeg2nrpQ/gWEtQHYhV8KwYfjoZczJw8IPGCc
GCUmFXsKiX4s4F8ZVEdsZoTSRUPe9SorhvgsZ+deMj9AhenA5Wu0Tm3vx/4CgbRfMJ5PVNX6SZNe
YtNfVVQnvpO/m0y8vHeIWZrYTHn2Da9vHGrI9B/a3OOvICjV+bkUWYjh/c1sPEIRVG4Ekp1dFAB/
Libq3S8k4HWk99fIEzXroxmJg+L99WZW5SX7yHcrpGZJIBQ0yuKAmytDGKy+VSAgZrkCh2CcQPex
CtknCZaadgm+GlYx/dKF/5BEr3bh9i1cTfmJaMsSs9ruDTI9G4sL/DcQtZWaE4R4FWmk3OzO634v
jFDy3fS1z9exkmJp3Rtwt8hLrqvuOfw6oAPPclFCw9uC+/o9x7e/MS4sI1gPJol4cW7luoZ4Mx2g
EAu79CwyaH9ejaYK0ynUM0Lw7tWHcov6ro841K01RoHDPwOaS+tAHaQzwrVu86uqCiAUtMJlkyug
/uAwdE+tJmpXdckaGAcfueRMgtsQ5/0KH+ff3vaJniUtFAYrnpaS7w3j/6blXtMDbdpA298Vr7WR
W69eIISqEdrGY0Wkalq4cMl2fXKatxzJ+CDNIYFas8Q9K0/+Hfw4/wcLHF+SHzQ6xYFNNVPOFfvN
miaCWFW6O4V+bXfdMVok/E4awI5iB1QthyJFFAl0wYYSwtp6Xe8Pw07nvpp/fSDaZWdbnT88uU5N
MC6EsgtpVJXPh/uk7oUQpiYlXH1oYxGeqZTrx+/GZfaEn9Xqc7HOqjy5WGDIgNdmRIvH6oH6XITY
R652TMSQQxa5sXo9fqRd2u8YSGSCOFS3Y51T01iV+utV9tKQiJENHDo5rw5+urdvu/Sh4IYMd223
H4jCCbi/MZEU+qC8oHy0gvXEHPRgNioOWmIwn738eRY3J41erBRiy6rGPizQ3ArYf90xqBfM4p8E
mIUfoIsHRMh2W65tq3GUWmrSgSrtbwH45IIInb3HhiXoGz/bFrI33SM5wVphnanOBt2ylBfruTK3
JYL4qwSeuoWN9qTMlH4qRglH8MrOtI0YSqIwKVEGWrdox3uvK2mezkcyxdv69XMFCNZTyeYZiLnt
TJMUNtB1VhMJF+gBvDs0fWTHyVu/Sx/kmPjLUeMXvh+8iulAxyHE5nFfXJtycpEipe2CWQaH2A8+
xxBtkINolpme4WHFw4pdUR3cTgeNarPk5oD7seCNbk7p4pQ6tieOWk8HStGS3TvOEVhoaqSRz+gB
fpTOSGckVpdxB6YihLkMgjWqcdXWevzDq6mGy4sHVjeK0D9GkkS75rVLZG5E7QaOCX9s+3IrCjeQ
q8qyiILsfpQLQW+kaIan42llgzS0Jlq7AdnFHHI4XkoBvYIB+jBdrqY0j0sYAQnxPo7QrW9P0WHG
OU2Br73fyJhHaBy81mNJjI4cmpmnv/irU8q/HqT8aJjVkmj3N8g2wCgc4SstwiYaCYa2w///A/zh
3dCFzZFJn7+RAdJc4lUKnOEwVChg9GYmaNBvRNuKw3cjM1xCjvksbySx0BIgVXoeX3T2wUgb87VI
AXSdd188wwhSDRH/pr6EkLsuXVeFc4KK6TtuiH6Iu/eNecnC3IvmDCXvJciDz7PuLXUSBBhFp8Ps
QuCPbKVceqU0rebN9mQWsh+fpO5gZ2ArjWyPq4DBpL6cnSENOXHwwn0itQtrJuoaY9LHvA5oPYKi
ZmHfEzmJnBuwR5NqVq0Ed2HPJ+SZg0dLhjbzZ/HI9c830050yq1+8xUGt+bOfHimEJL/CMzpmWnn
V2XCrzmN/nme7GIau7jyBMCCUxp+9rngXWH/iqMnvgGngd6bDte5ydESUGiebRd4f5e+8aTd4gHg
p2ENxYDOT52R4GPQHqIvtIH/aV/k18UvoRcaeFDEq26Ga0GK5hQOxGo50PKlFntOUcPGtln1ZeDD
Nak17YsPVkLmSa+PNLxVFCWkwZuG2i2cSnz082fb+doXts1mFerPUHWwd1ssRxKiabX/9kcheiuU
03HuttN/P/XHxOUQSQuJfLCh61IilmlUXJmaxWpSCFUoG8CkucHuDuBkUQ6pp7NbQGPDS8IIjbVU
WcC+choSkCZCBYs/n9W1P6pdzXfpcfK0w8JH/IY+bxthIKPY8ZbPd62Byqf4LL2ofs0afDLXkRRI
Kn+LbmPTyKnRRnSYDRzr+lUNp0hdbg4CfzVXRiGZ6VGEudnhcH8g3NeCdPUgXSmXZh2QcrhbW/i2
gRyy9HKElFqNZu8f8yLdG1QWg0n3o0uYLEevtEW6xeLX2WepUKjuHiN/kjKJBIGLH+kaqXk5ETL/
CeDf8eTRe5/Lk+hrM5wNvMXRNoyMNC8hI7O1I5egfHfOrF0X634IXRGugesDt1OCPvYlacOmRn7h
GlygG8qnktkxHJvWm1B05Q9ysRuk7E6GBvOzi00oILjBn4g068vuy9cBxU3UBFR1ilgB9qPIwcVm
kVZJezeEThH5dMeut5V6r9oRa5kFjcmNdvfzsJ3HNjllV3O0pQwVea19lya1mZ+B5DcktJQ0cNve
dily0IRYTFckttlr1pJn+14kn95uMNRf7m771doCx7ALOHzBeGeKSk4jcsRtcxfzbtdUyDb4Z54u
EQbFSJpNjBq1+G603zyhDMXrZV0llkLunuWUsr872grTgEeEPCEopfv2ybXw6RyADBTb9RgMbLHA
oeTbuNfm/MElMJf0B3q6LcdX9v7j0fWrwcTO1iQh85Buee0tjVzVmD+WKwbg809KhAVSrHkCi6Tq
/mLX6UQzID9sKIl1Iyc0OiAu39kW3xYMmpnqg8et57DqNLUWPSL1JBC+WYGzRRqdJtvSvtzr50fZ
ZLRBPYhzP0N4r5mJCoxndIExMAz7Q1n0m2dahyE6c3PoHv92pPOHDHoPyQYg96PPn+hhVTMTDpUw
THkL+Ub402DQyjojuRbIlz8DZ7c8/bEsyJWoiti13D0CijtxUwVZW0NWtlqL1WKwmcvCbZk3z9OX
B1xo+QUM70ZBQvyt1R9cw9T83zq4lb3i5SyzUAT/DuxQ19fV58LLnbU3SgBOMf9zmujKfZzkdC4n
hEmoZ+tFfvnuG+bTzXayBYXZuZBTrR8u79BPgLkJzDwosHqm2wyHMnBJ8Te40c8BtR6yo8JpiPA2
odvVkVc+VQ2547cSk6iV4jQoplWpfKJFuNYARuigGx16u9XuVo28xJgEtZ6MO66iVh3pEuS2LWKI
T67j5cEnoqITz2XBBy77z6Ee9LdozFX9VmWt+M9u/D6o4UTxdKRhV1KIQh7eWee8o76cFoW68AVD
NCfvynGZCtjS26IEBSlLGGSdLQw3Gdy24J8xA2msz6ZdLQLOV1icMIgYz71b/aYKrjbTcL2/ca5/
V2VXHxnq80ze+E8w+lKGh95pOaUAjBmHDanbUb+UWq+YxfzB1bbc5CrVS9h1VP08Af0tHCgxLOMg
rY36gBsyHwgnfrU2FXypX94c51IqezUIRKDwm0WIIImMnPYbVbRZCgMCfaBKZY5XHcw+k2qW25Uh
79KApH1ZUwIwK9qhWutx6q1ltrTjvvOQJnFFmWkppzY7ALUfQTHW2HK8Tec9bZft0pOr/DoriXOQ
xtsMwTBPR5UwlXrE0t8NLwxmAf4CFQ4StURxb4m70CaFkQOacScd7hbG3yzvZW4l2+32AlNdkC7t
ccbao9A2e+djCiA21ZdleY0vu0u5VYTUAKzALrSyRNmvryi8gZDz9GZrsy5AhZgFFDJL08QEMIWV
PVWWUEFDG53V1rc0O+eCYfSwP5yEMkCKkPqXNgAgYhU6xZ1hjvkE8gxNvHHx7/ysZmI9SBk8CYS4
kPQn7Gw/zTZYlazkjFs0Pu8fZlO+ZHZmwlC1IhdCeEoWJoc1tlKkgWbJvywX3F2ttlC4RpDJ9d5D
IQHhWbsE8a9fMxQ3kmEGcDcjQ62dh4yRfTQ38KkBlCxf9/ijtFzLWJkGsxOqAOc7VRQCYrzRbjAy
ME9h6w4QmNCfM3QrPpVpezkuABK00GiH6BSt8P1VJP68zqBWy20kKEfTFDy5aKLoJcwvcvbBr2x9
yOkLgXPZMNUzyI8Xke24WrygK2FXqTlDQIql5wBDcKAvPKlRVQnEb2IhKqs3BP+0LtMRLuQ7kSFt
Nl0BPws2Kmmv+SuhpoJHt8bHqYRfhtoyBcW37zl/k+AxhjYTt55eLUSn0t/AIwXpP38PugKKBp2J
a44zI1hR1uf6mlhb/dnpBsD/BaO8062od5Qsa9s349of6KEZZ+1j6VCL3nyeeTjG2WQg3Rih7Qf1
0f0UiAVCscbBdJFD2f8+QJ9q4S8xXxz5p55LaI/TvkY07pX4fj2phvoBLf8XEzvrgXWRnLbIvCM4
TFxtek8/sh+QsmEMjPJa9wapN67DQGz6Tp+GFpu5qVIHmTpgLQK2NwFEVyyl3IkYy/GO3N+YNN/n
UfFc9F73lN6lvax53kkCiy3VqhNKVIR2Nqdc1Gk0dUEuxPQbdFw2PmE/OmIigvRrtcpdGOF7RYte
vI5hD5quVh/SeYOQ++9mduXtDLC6nNhh5Hj3E0ECdAqYKhtRi0ovzCXsKOXzhlWf+Qvq3eGZPPK3
S9gNhankf2OuzSvro7115VsJVtXN1vT6ueStwN0Ex+P4vPtXhgam32Sn8cBFtlFDgipfpg1NQ8RE
0zDgGvDB1IaJ8zOPSdsUinYLgkgBp6Ic659YMgNCHRrOWP/C8A5DNCkkKayHhGlvoPmYeCDJg60o
mzBT5MsPZovrwdm5PO7fC+UkjYuqoG+0mxiM0XwbRYtVDuZPtn5NRSylfCpe6Uu/mxLwuWfLPrcI
k88RtEmO7AKDOi3FI6mW2SrQawseGTfKI22hsaJZrmoJHwWBY8A9BbcPezzKSLgpfXhnW0YEn/AC
ZcAL5gBU1ZJkNihiaDTbYfdC+LXskZ3By746UUi4tBM0AFxBKR+6Nqhl9Enf8KfvdQ5OIA1UBepB
TqBkv9rIDbirMlGow80T3A7OFViIiSmuGS673ICSZ1v3wK8xZdRQYiqXe3mrd64ZoAiGmkFmualu
MHWuR5Fzx2aa+dqv6bRew/QapNMrcFeOhqEsj+3anjSY4cFVaiNYXgTPX/gN+wzKz0hisXYwL3Vh
X1famTjKSxYDuQI5lbKDhMSyhli9fmPNsgPqJblva0/nUHIAcyQuaS1bimB55Y8PO9sUZnX0CMct
R6pE5qfhiIaCjt7XvAwq1SZ3EQOoO/ie+jmkuccM2gPM90OCP2NqnUwJA8zePDUXHXl3RwG5GtN4
pbpRLY1pWwYjfxmpatbQIv7ppmu0cG5ughwzEtViSogxn5ufSLvQPWpPbNQAdtqPrzh7NcXSF31Y
MaWtELk8NVsd3t2uZ0OkBG/Z/CgjrrDw2C0Ey/Uw43WNp0BA+NRtm78h+5tHq1Ci5fX2vJgDGvyg
PHOpHoPhyp1V0JNXfspTV71pwjlRDn/q6ZCaO0TLbWh+h4fmLwNEufdocP7XHFL7uYfF0r5XC+2R
MKFHuleHAFHQLTvQeamF1UXuEIuTKmb/z6PZuOlSxSZfMCDbw/pgxClRbFA6U+Na+kvOgO196OIX
HV4Os69rfRD3gODi22TWUaq9by1kTW1YxmFqPg+geoyLQIg0cQ78jMKbWMvrynjpaM+QIjh19egW
J2BBqyWIY8cGs5knk5ejIAabiQCu1pk/flueCBPAAk0kTJR0J3R/p8yRfIJHX9l8/gXfp+xvSx5Y
ryH4tNLQu6RL2GH4zzo6Qh9FWKTaNy6EzonezXy2TsozqdlrMZJ/Th7O5thNU+5aFdeSFWiBJS6W
0tPzmiolqhP1Qz51/QaevBodY8BTO4AxvVJ+KyMoLMDlJQfGNVSPktmZY2nXp4LdXyzOLCxrK5nR
+OJLtUuG44rQU3mulRz/D+K7x3OuaoBhor0zW7M6wSjnu5BwfzT720Fk0TxRqwjiQHBXuKLnVF70
yXh36FtNFJtf83OsWaMeTOkqTDTj8ACAgYTc5Qi7nLR6QldO2vuOQUjHL+VR0e0/VQrsHOiJCwPT
EcrjWiv2Fg8U0yWv0Iuosun7ANVvimTIzhavz0UAfzr72xRHmzXUP7aJTBC+dZUp1AlIb5hkmcCA
0hxjr11qx0/yznrGwo2yN/y+kUhhHI5eSFutA5utQip9RE6HKvHYo2XS1cXnCCV7FRlzw+hJgCcd
acHXZI1I8AZBWpr+kCGdsXnRHlfui5/T3qBMwCD8AzOuykZCKdf0cNQGSJiH4pzKFUomAM8P/965
H1CQwXq+u7ELM/FJ2pOw4ATG5tkGU6dwW4J7WJyJe9GHCvK9hH4moEXO9iatAuVRUCsFV2Icn7np
vOp4s+1hsWEXxVqvCQYO0VBZE82s1CkdKBmvsgjYCZvo4uOG9JMwc8m+VfY1EiOEKeGJukNU2+bf
CqcEFufa6yYth838iMg2UYKoU7O0hhjv2rCAyk3h4ACYPmPx7ShUmzC5NH9q78JW6rOTs5nKFdMp
hIVaLOfMAJEcOCD+c4YQxJNa3YELhmZzCBn7z2YfFDFAqJ+N57J2TpzFbCYqNzbywx70cHpc+0M0
KOMVlvnVk9zSGJoj8swGduo2iU+D3NUXyT9AYUlbUwRHCnN+WLwkzehiBAVj045o8vDvp7aDUU2e
sQNrBYSn5/Do7RbiEciGMCkfMPHB0Ymu/SGBxXsVdOYu+42pWISorEzvQofBrlMJw95wWVLdTlw2
KmQNsBKgBboj91qiZHUZfWePFZD1PiTnh4NJZxhHGg0sWybWwtKrvzg+NOkwtb7FAnZYyrGdGueP
xZ/25Fc+JaIfUZobLsU1Uo2G9II/wJ6IBLJBIk+EPL32BHrb2f4IjHB/Qrk0eSsevLiDVDOxIHfm
M/ER226AolR/ewv05JnsgwtloWVbovUXXSrlKmFIHeeuO2t1f+AoqlF0xqX6yJ1+eymqIjCbxafc
DU4dE/+bhYRn6qOygfmFGtroDsNzv2mWBix7mFeB0NjDExQbu3K/CsBmctVYvZ7slfx2xVnq8TNc
Wkzx5SdDHKL8ZHWYkJ4iOnZcZBtwafjq9kG7TY2Xf8FRdFtIe3dVRcuCPYBlkD4e+w/lqLtLTf+a
LHOJ7EdCIkM5kUprF41gwCYcsMmaJJpAWwS2VPqBju649t3oEgfUHlXsSSzneF6uFsJhCbrPJG42
cYrbr7Uj5q78WjZdmw9qCy44LezMDqxF3AJZsehpWgTk0f0Op0dLfPbMtf9m+ryg2wqUrdmWIR8Q
aL0Y3V0uBUzpXYGkwrkwPl90pJkH1cZ4jPsl2uXdo+la8y4pt157CXtkV133mAcgK9zGZC4EClCk
dJ3TqD/Y9PkkSKFzEBzWU3sk7F00mvI3EpG8tw8WI6s3BofNFIDRd+Q/WYf0DT5vkdClYyXiwKyE
l+/c0QusN6awFDrhbVnl57edPMSBKZNybrcWkAGn3A5TGSXFKjy+4zTptkHNhgsq4yYqa+bZrXUP
+CdQuttqiNI3c6sWlMRdmYt2gj+GOO87kaoZFS9TGHlORBVTiX6AX92oRuLM3p+fa/rPyfnJY0CI
kByywkMsLZal1fgLmwuD4pMltPAMaZY+c5BDZBE8tLP5jA109xcDc2H8poWkdzy/CA9tMkcdtUNO
wFd9/vh4yPdfORgrdelx5cV6XKxP7Q18N+HoC+qNH8C4gU+zBdrMm+VLfNLO1ZrEApEQit7S0H0R
muAS0NHJePt5ulvS06tBUutGfCerqlKYKUivPKYVtWlNc3Wv+qO4dFbEWhHHC1YWZYSqEdT6rjZ0
TicDj9n8wzkvd1++O07VMSh/z/Mm627SE2cnXyL+Wet0cFNe1rImnPrC99giG996Y/JdZNrCsH+o
Zj7/zEjdw42KpkX5SnfV//cWM3fm6dPJt/bkxBTsvMo9DtnaZsomTWcGU+TCY++4AsPJ04zjP5ge
T80KdHYG11m9BcoJXACx2BchODcl7Yd4w4Z4OtWhzD2YWzAk1YLCMrFKGZeYcZW8szIOhAjN74HN
G9OUIqCzY8oi5M9/P1bLoTLl7zV9wJGltsLEcuD9h7zoBXqemotskBeUXyAj86XJb2hfuknzoZk7
hd1sSa7yDKvmHX67dgjNiqeF0a0G4oqADJZ9E+Rq2dkfiAFcRWZPaLKxsI9m+XlUKg4StSwwDjRL
royBzrLg7B+UIxg6Q/Nhu2nruptvAGsAOTYa8OeE/MVkmpwGvu+Py+NtmOdXndk8WR94/Ru/ScFa
YOdjk6JfPKN0Yksjoig1nb9uKJTesM1ZjjZZuB8EGxdL6W+s+U6uY+9HPd+t15vC/1sEHr+m743Z
8W0gojhwDMdzRruQ67C9O8Eqy6ZoavQAF61kHWwopVY1Y00ocCq5Zb/b6A22FgbHE8rt68R6Z/i3
fuWeE1s12gk7/CzSSUfqoCOy7c5x5ctnmVcgXQ2LmsLNJVHqKY+jlUGxEZIezDD87A2xLSJzc+g2
9MoKkUCJNxWYp5LPAKhQ+NAao7Tv3V4oRtAchf58xb4l9TjWWGOVqJLOU0hLhJwqOI0SM27N5Vb6
NU0GiqEnUcT2ZgduiezQ8KrJXhr9Fd+VSid6kBqhBRNddp1ogAKw6E5khsqJWxdmAn84tcpfdt4b
KpErhvRn3aIH5NfA4PBJloBEiWpM+ZsF1BwIX4pHwciiI19GbRo/oGMFkuxVMUOJvdElXbctInVL
8tEEFTjZqo//SPqSF94xY88baYZfm/Ne8qvU0xgohIqzSsRDJFFkHI/7jq0HB/blnpmdK49zBSwL
gmtseIl2MZdqBG4SW+rYSAQOPm768WgRKNzMOYNkzYAzeOJNzlgirPYemOq6bil4f2grNUOKqNTl
J/AcfaKZaisx45b9NBM6Yzh+TtmqQaCMrPq+SIgJUvG0omYt7AOWRZL/1NGcaH2/49ypxZUU9yFF
Yo+fetW93SsjKSswQm+RQyA7MPP+i6bpAo0mGDsNuDrOva5AT/wprn6/GFfl6B3Hjmip7DtYRdlD
FcXmQ/OHb35km2B4mi3it10yNlM8I2T6Cp5WRWLb5M3V/m0XZZ2xFFuE+h0iDZwQfM4ya6DekrCP
h1fuf+EyNRe4cMDjzqVFrVXyw4w3WuEtR0ImuebLBn0mosJH2x7G/MWjiZOwr7Vx5+/Rd25czp1u
GNQjmSOz5L13CN++9O01SAMdHzUj5rYBVBuBViRxf8LW0PRpE3z5VR6div5V+zVJ76DgICHzfEp2
e4QO10mpnnXQEwM43ZDUPK50bGCRes5aQm2PgRrhfNeuvqTJ4Fm3v+dvtci9wf6vBKL+0OP2XlTk
X6bskgPG4Jt4Pcppub/Y3F66cdSf0FWdbK5I5Scfn33X3NpBm2UTWWN4fPxIn6PyCHIEKDEbT3+W
IMvfYb8v0goKRNbM99KYj7c/pCEaAMO04t5L/Cr83EFmjVaPrJbO+1jT3/v5HoUHKv3c1ZycnG2P
qArtU3KqafaQpu5Cx1Sx+Bl+2Jmm8kYfHKEmnIfORr/v9h8Wyf8f7AJKHkVq3hxlAGSwlHG6BEPi
ii0oDYHLuKHuKmR7dAS8PnwqRGqq3vHcTGA5aNi8B2vhCXqZZjMn2oR1hJWqQMNs3TUdCpt1lGQz
WhiY7PSHGg9ur81aqBsL9jB3lz32/Y/W2Eo+e4V2ApwfVoRcHpKKEmuGG8AelGz8AUK2wyhMR2MH
B7/TgOc8JuySTvPjmNaOra9Qys4eFs1+Byp0/mg8/ro+LW/Rc/ChOzsfxtRMFXaUpjgp0oaPcFSO
7TqVVjvs1kQOvsJpyJQnMysT546Hv7ozJitcY3Cwql4xJHdwXMZucqRn7bGOuz5T4p4a9FdNrt8Y
ipmYG9wcYzkHQj1AONXezfmuG9gH614y/kzO8hZG0Q6OV37+cMa4/oGPEP+55bdQAo6JkLdlpmFH
j1zXYcdGvgnmRm2fKzkXOnHqEWHCKVRS8xLGWdSdKgFCA2H5NEh6ZbtAFdtTFlbBd26nr+DeHtJz
4SpHVaKfYZxCQcPg7o1XESQWKp4rB7v/96XRmL4nm8zH+z3mT5eIcXsAuKQPZyGinyhJ7p02DaE3
FaSXC9Ar9CceDnC7Qz68ImHtWOYvbBPvavTaAuKcudqdqKwPeL+zHO8oncLN7y18r4rFFis+xoLU
CoqdJbNBAsSGaQMKH6EHjNZ5r4Mhz+e81Y0VBw/vCPJLyqJr4WiCaqdUyTHR5/P4rDZLJiVZHfPg
LR+o6YToCJrPiCdTZ9MfSlr7WGK34+Hxlb6reZEbVEHbljNAEMCqSONeYZWC0WqURJqWN12FbKMY
A89dBwz33AtZ92M7ZfJwQIH4qTWPcoMo+gNsVxDkRhEnRANSgezPAuNAXn3M5TrHn/m1PwcRmGOa
30Q0TFxdr8ykwvLJyT/+u7kD6Jr2YWUVG5HHI6zO8+9yz5aP5KhKuYYV32Dy17KglsWrpCs+03Yx
6qe96fRRAMMm8xf1BKD6tC3MG0euSbvhEv3Vj9E+rGhG3Gj1rEcPUAtPkVS5zTBDrtmEZNdGkqAl
UDrfrbEAbUzf6V/FMBaJqX3VevF/F5eV4kn4gS5dwr6o5iL+hb8pe1OuNGMbgUF4ZN1+RbFUm7XL
2izRNUWbiEK/xslkCYyrqKNVSyIHK80Rc8qzH1IfqtnWdzDTc/QT0hxu7mp+D02kXMcUMiRzwkdt
zZbf88KJe1DlK6f9EemQvfKnjQlB+IrZG1d5cbLV4jIxb++7MTl9n4luOLci+jnV0hlxS+J6tM3C
1QkZTeAbDMUG619GR88TJmNJde/U44MJl0mx1Ap1QXWkGf/5SNMSgqwTUmMkNdaotnF7GcEcain6
CLq4UxJe+kWovXA+e90GN2XjbE4VzLfBp32ymqPfOqXFT1ZsgDBjUWnfM0H+5Ty8y1JjuodFTezI
cp3ODwjBtHbe1gEriZaj2rUI+/mDV7H47QRZXE87UyqmP+HMd+QnZ/KZsIH2YcZR9j12P+leB50b
JB6O4Izbo49ykmmgrnROP8LILnM+Qdr20mL2Tpr+lwL/S8J2nDbb2QyZLFL/qxN4vNd1hz/GCsUU
xvrnHaut4XaUgAkUe9nXmfru9NZynovfHbTMdk8ancd0KFgsUMctiPLYwUeT8Idtqy7hjoMEPZ6+
UCMm9Q2p9gbfFuL+u9Ve742OWejl2jwZ9LcTz3Vpuv+sPLRyqMGW0JryhKp2AsxI9q2koE7DxtvI
VpW0Z547HTnp+lXzBifaOQYlW+XEbWA+z/pnvqmxML0YoCneM2fktR4KwAp27O+RKfjxhshqNwjp
tRAG720dc5+ArqjZR+ouk+a/2Yxr2pHy/R1RjiaKPJjQQA2aIfXHeo0S+JBhhgwI5dBZYJjdOjH2
nd7SiOUGdH+hp1Y5K4ErGt86tvl22okfVe4nROaXsHqLIjkIG1E171DkWnYqBC2zs+WUPRcQEYMD
s/CFK5JcXnfl9soQpvmVajgOCpZxCx6CtkIoMyiikhayZh+hnjzxWXVxFrZkhIRPYjFFyr5ppcvb
cIccyJiBHQWvtBbG6OOkmeit/7pSWZACXlINMLNiiPYFdGqGJo0MY9XSfqrMGt8wwPOPVAa7DowE
+NLPU7ajWflIUtjs02GQAgPJe7KY5bgnDWNYGi+L7Q7NrLg0Pg5p+8mA/TklfN2M/UnVRXQ/sXUJ
CaoUqSOILgBpz2KlvbKNGG8I90bzGmuZVtj7NvJFLJk8UzYeLicc2x7gtZJxDxEvSJDsrC2dgWzf
UD1r1Ex+D0mn/omDZzHuoMmJaN0qSggehgZlT6iBJ5MwfF4WctwyKAnOZhpQn06IIwnfrY2uuNFg
HrgTudcP29f+wcwd2+rWvRDhkZ5dBxfAGyIg05F/Vd7Qd54a7ny94nJ4Zq9wfvS3QfRBiK37OOSF
YSkOu7fOcu5qQGA3Suydqi78/9IATxqCyA0olOb6lIW9/SiwWcDmGbiMMiK3OwjwRqAXzJIQM51R
fuw2HcaWi0sZQGKjJIJtLjOoVCIUXMX8DsVT4QjHFMJTDZCx1Hs7GMJxOIUtlZpIBHu8JWbP0CGO
OOFN7V6HhKLKm8sdcElym3N6aLchYUPUM8agKv3jhp82c2SRZONvsWdm2Y2G3kRIWQoy8ogmnjhi
v7bw8L4EYhvpuAe71lQpxK8SYUXoLfNJT0aSVoRXMHQmQg1H4LWRBFu85vcgcc1AVNHUDJXRacuB
YKuabdaSe/zYJLW51CVct7EXqhqrrTZSVfE78BWZs03tIVPyllPTfcd/U+/YUTvNHiL9N98xiMZO
kjmwfkE2eoBubAMbhgthNnmYQtYqDls/pDzRRYKblQnJakyXZ7RnAXcSc5bVTS1icVsLZuxZxEH3
sSEpmI9oXpRmXjHNDvCuTMDL8OuK1uIfcBNVKvPeAQ0rJt9GGTb489YqN1ixnBS4OSfVHU4I8rLo
OEetJ0qGZ8N2UtrhcbmpAV+bTBsHCceGteDYQIzvrIsvAKa/Ai7sCNkyTsxyZN1kvYHcBRnZwOGd
uS3T0hL8B2IWYi6Dor/TvINqAp1elRpiP3zyIClzxMMi74Ni2mKW1dkzZnL2B54SHiN9u3OsPV1Z
5nmL21slyhLAdilo6yLc2VG+lQ++VgYuYOVfpHlUqCLbJsl/GjnCIIV7qEN5d89+qqTaTsfM5Kvm
kKsE8x0/uxTQx2TZS110+up9eIL2OjDAUxE/xxrn0eWhByig1YCX+18WHiU6EiQXbdLZaMqDFeoV
0GWw0GP7wZSoc1+j+Wu6ACMvGSYarglR/MHbYdfCQ2HOZO68tNoMUP1zJpixWw58fkFrPehyg0mN
Me+gTTLBhbZK/Lf/w5QDB8lMq4Cw6WWIH+LSj2uEpWw6D07R8L9HEcGqZ7p1n8Yao63ZDxkxrn1A
IM+8veFvLeiN1ih0e30jAh2yrpNutwBRXWsMv/P5FrjgrOdpkimtb5iNnxzsJnPZ2HyksrU6+KNP
bhQhuXBxOdOvGKkM+k0PEq2iKEyDefcigWC2a9q8iuZ2rXFPlpZBtO1t4cLRtoWZ1ctN0dTK89aq
TDf1ZaqXRUSUASPX3KVSUCEUxSx8dUQKXJIOBmxHx7rDx3lU+xckBz3fIi+oIgNSzMH0Jc9u6cdw
K5v6GLsf7XsNqpy2IVOmpS4cOW2sOieHn+Bdn9pYp3yNSNSjBVJ33D0WTUpCcZ2qGU2f2JlxXXPk
FR4SDNZxviRyAxezobO0t3cZJatl+wl5MWifABg9Qu1+4MvyHoFUu21ULzov3pmVcbJt8MrajHU7
a0YDSg9wQpTFgPRl//GBn6kUWZtiR/Ww5rG3wiwSGfxzaiVysBgdZlch0ZuwsKiMRC5EfRMFLGEe
ybNaK7z/b1vQVQwpC7Mpd81ck4QM3CGNmheB1N2VroF93XaQ758fKldtBE/u0ElezfScS5SrHoZx
WMLJIb6jCYUrAD4JUn2RwLg2dn2tbbK8Ae9ged+A6aOc41EwfCCL7qS8LXdu6KmrsWqSsdOb331h
xQJHWkGnLopMwoM+4HM5i6HkXFhhVXjsMJzLrhnEZG7yiyFpBuA1uhKyteRIk6wpQXsztlcwjeRY
ZRx0swNp/NrdDagbflgotRxpy5SP4sls/rp1JyieyylnFNbblYEujPGRDfebxaP++bg5RFu3DXdq
akmrDFKKJJr25ZZ6Y+NPIHPLVEV2zfyGuXCkDAZIVvxC6d0wmd+zEpaFTzysBtRIS4FgwoJiaq7g
WGh1D8U57CGiYBGiDwZ7FFkHqhyuZIV8cvvu79kfjoMrJ8RAkVKyUssW3NNr/0RExnRmSv4HfbfA
B4tY0W6muS4ZOYqIfMdnBjuT3qmnjgFNMy+QF2Pr97/ZbpGDpfzcBjuXcxmNfVPVDvZntaJpiZNN
Yshsc+UvaXnoc5539uWaaTdq1vih8VKfFA/HSyFVkhh/AFx4hX1Mo5b45oEthXxbdJClXWMwX+qo
Puuhx0YYYEqBfLJ+9dJtqn0vXYo7WkonM0YjGEh8/sEkqRRbz1VwEsw0Z7rK+NDaBwG6hJqovWiB
0D46fTSq7b/6JqE3dF6FIGTcMnRNbx/IfJUdDUvDctF6D7lIRsdOP+DvmWtAqGhPcDj8/oZoCZTp
npQ3XqCbkSjjQcT+0bkc2BenPDATnIU9+hLVovgQvfK6kk7ttMKdoXq/SkGXSvLfke7TP9cSdmcL
XBskYl9l9QpXD7M/cUeT4lcMIFaOGjF1tpH5fO3ychVp/cJ3nEu0ALsn3G4a59iPwmOl4G1r4zBi
p8ZEA5UNXTii00lO/13gaaySyLHAkg+qgc0kGe50F5c8dA5LmeJqT4PSSZI2fH6QOBwD3OB+SBJE
FU8iwLlhlw5YkUWvJVS3F2fbBoSSJLstqyrfBCQENDU56a9BLKZIY60BhZJXpWxMgQirhIZexOZ1
bfG8ZlJiyWoxG9hUT5akb19i+BWED9hvmzF5L382lup5J8aBF0qqvc4YJFpeGcgR9+CUNN5MOPSz
rocTnHjqNzd6p4V+N6dHl16DTjVlOX5UOdIU228c4GiXCJToWh5M4BQ6ph/Re6hgsHt6G72/G8Qt
+Z7kE9Q/XvS3snz3WZN85AN4BsOyU+j0naIvau+2cxqT/7pJbUokmdjxs2+EYOS6vCfmDZxX7Mcj
veFCe+fzdF+LzprnZ8O+FzWes2mTbGh4F8kHyXvSPBhlKpqFw693YyCrx/QxuSAIGKvWd8E7BRgA
7f+8DaVvkmkn1MGboom874rFIfQ5L//A1l/SBS6cuZE1gculL4b8wiQY1dNlI8cXHkxGJEUpStxI
xY+ousNZ+gr8GDrHYD+6h2i59Bz2xCo13S8yYqeK0Y72A5VV/3AnNg+ApIIrfSaTR9cidzmPcqD7
M+6ky7/iny/dXtHb+ZKfUlp8eU3W6LbdKDnAS5hm5uvMseC0PGzPyjcrnWsmtkF4kxc7ZCHGPD4v
R+1gInBzX63BDlLtzF/ZVAG/v3fOd7xozxWCLAS3QaZCXDMDhsAOWoaw/TOposbdk6YcPij/NPkC
cUWvLH5RuHwO7Z0HnXdT7QTyyzkrIl3qW4diAfmR2eedDelTlaqOUAhQRoq1YjnzYtB8qIRsLjjg
Kmuvcuie/LIn+z92zLikvdREcnmTinbULHbAr5e3XjfezEkQH/6jWeuo/AG8S9pzr8d6+WIHpK6F
4XJOQ6Woagst/KyiV+OON3RvzYXPndF9CeW70TFpIXkoOpAhewEbDBvC6N+1TBkgCInaZ/np1bpd
cnhm8MtxGayl9ZWROJ31olClZRCeo4neZrfQq7Zhr00/yFy+vrFCI5BcH59DIx06SzVD6mwRiCPY
1PGPRtllHYxqm3qhvN4RTZ+AgShgyQCsg0zkLedcW1M8Zr5be1eq0orXqM5MyFfVAm5DcaYOcRaI
65EEhYUKEsNRuSCy7x23ON6U9Y/VZY2Jd+LmPlpzP2g1RaaHJskB4Oo9Xcfi4KD8VghGlaB2oXSk
5fxZ3KK4kjEQulC8gOaCSkKHStlGRAzvGUZ7xWnFNI4+2YbjQlciK5w33FVDtHtuyrzL57YZtaGv
+qsLVXR/pWnfYzLFuJwPsW526F02v5NlhTCo/lczkfDw5ARH8Yj80d4JgnVMP34udemNGnU2RAVC
3weSgwdFsOLsi+wxo3rAoKiCQMWEaRjhog0PlJhZ+YlcONgPfY/ap2c45DSZznt1eqoZUYmVbbJG
FB+//PiQSOQ+ivM0IZFD3V7/tKnV4yrNTqOsukNgORlrq498y7OGCjPVmTgc2hMnoTuWLRsMMpxQ
dB7haYZszECMMqcTLKC0Pd/O76iOJkO6zH8UZNi0/kyFDYA/dg1K5uxrlTUXPnMzK9MdwczwI7AC
cvvQiqglSjPQTsmBtQVucVMr+bIxQyQADrCSWmjltjp6sjgXvqdq8+e8VCDMkG1FAgOfBbZnIaHj
2LNQG+S0KvVMd1OmqTlup69B+ZqMms+ogLvj46a2X2kUQ0fTC75SA3Q+tppobUaFz51aUP4Yc6Nk
FX3sNnPhuhqYPea6+uhaghCupDiFPWBybUfXL1NPPWMo2hV/d3nbEupO0z4MnJ1XGYbLLjWXACcJ
Vcv6YkPohCkzPixMkxjV5SCdxYsfGh0g7s+rSIJLE1TTpkuqtjwOPJdOrAb0D/ZoJHK+t64DJllZ
cSQa4rBykW/cJcsC7GW5NUOWXCRRXyrENPIVpFm8XIrLewEmMcVTz7i4N97Wm/y9qYV4sPDXGkQj
RPb1UNJKGGTXq1V+OHGmuRD8pnU53SKmepSlwBC1DMT8q+H1J8s5itWBkCJvM4MdKRx19QfZK1m3
vz8E7Xzr9Tdv0Ks1KcTXl9XxiUt+CKknIc7lyIZqvy3n6GT22hGaRTQyzZF+JBKFsONnjJ6e+uYR
20J0fjs+4Ti2Cy3Y+SDUgVJPCi1s5VHMwZuod/Uf4QOGzxB5QVaPbiTXWkOLlDYaUNl8ZfPEdC0A
IhJ26alxr96LKfxwUWyWWlTTJzvt1nCDkHtus2aU9cKYy3NL+Xdk9eIr9gulYlhw1sZZ3Sju8SAa
NMldmPgjjKFM6mLfBRRKFMmIey39hfEqLyF1cxiACqdeGcqOmEb1WhBLjus1Zy6JYSQ/apSskCmd
JHzipNdKfnT5BFN+hFFQ+ojmQn/zha4BHCNaOxIiH6k6OcOiHzBIl+0R1BGyE5Za/IFjtdf9YwAd
Pma1dQlrYVctwvpYbu8PrJmC6n3lixePWHHYmKkSdz7HQnxm5PWIu+7AbetrhhwcO6kQ0mWOhLaW
skWfxuF4IsGRrEGm+cpcQocvgOI1FvnPqGm738p9ossTbMUf0Oo3oQn0zClaU5j/bOaiSYLAt/pQ
jNK0ySst+oKkmIFVR6hdh7KrAv3jyDsQ2ywtNMkm8qn39mvmq+kiyzVDPJIge65tkNW8BHDSSgzj
+CqLB1VPVIT7yAbkPxvspnCK/+GnsqWXVkG2gnn7NuA/LkUs6SrLCr/MFoB6a87jljDE8rV4n8z3
m4T47AF7yc9K3ylQYMYnRSRQVqTJ+7diYjVB2poFhbqXMw8z2fT2PQ4zYBKjYUaYZldnmKcRmPz8
GtqGZN1UDn9Yh53+RNu1Jmol9nhNZXbDOpowQbicf+PO2oGwStd6t97SHZLEB/V0JFb7d7fAwJlb
vmaqRJEzO32fNZSRtyDlQ8fJWacICysYwVuLUofbaH9Mx9qX472nWVVUryRQWJzltnzxSZFIK9oh
EDMMHA7JOxVABpeUKwxq87m0pir8J5TvNLb1ARAqMYKCH3LsWZWGbhJlyCpupylTXjmbaANMlCk7
G9tZL2idFnyvTXH+nWVrkjRDV+yLpBzX3pzF4V0CaibUbcWuZBaSJ3Z2GelAWb9iEWfBCFKp4d53
AEI8pawj43Qw1P13pCZbxYU49Xk32xwArFQNVntMnLGpJmj4nPfpircf5FaPBvCleK9388UHZYV9
ZgN5SwZW9Vv53srXeM/c8L8o1Y0vtruM4ckUDyNrI68GUSNuWvHgCz/IKp3lWGLwqcXkRoknZtpB
zS5fWbUH6d2jo19miKjAyVB4Uj74321KQPJ+9TzsZ9UDdYrJRACzmKVqUbxIw+UD/HzMt2b3Syek
TL/CJvcKOIBnAxsq8qv1laQO+B+FFw4IoIgxjbxqELkIiOrDQbu1+hu5M7uEBzwmI8ad3LbOER/r
U+831DHVc9fUMGSbsmwb4DzNI4Hvip1GBydXyxJdAI/i2kDx7rJPWuiUyVQskwGR8KSRv3DFB51x
vGvazfe31tT3XBE7ntaS2Ai7M2hh55I76HKXCz5B+rUlwwT/wfWw/Ib+EHVhP8CMRH+Z5332rs61
v1xeARwg356s4hdXAmksDZBRDdJ2imRyfCAe7D2j24VhYqzJyIAbRtyDMS6IPXAFG3ugphpBJflj
Yo8O+dY4oGjznqBGRRczkqFxS/0fptz5DMQ9mysw25VwyJVM03PLBTUxh/wm9tyhekM+HcGHw9tL
nZpsKXVMJyJ16vWiiai3xFPRdNlI8fZO7P1vTLWjlLlIwfmuZDGJyFi8qfjHF20+FFXYdd5stIcD
CT0wndkKeHx9KqwbzItPM00KPL+1gQzSOucOb3F6WsYWiPEAH7XvpTascIbj4i5NCJ//uFlpbY/g
XED/u/wsEEdmvo1LC2xd5GFRJ0FjyrVfXDB5wWu0JSgDnt/zyLBC2yKXEzKCs9eMY3jmk+77Awlu
rcabFWOqUbEEDNuYe+k1IHO2LH3wlEbOnh5p4vP/tRHf1p1L0Q454lGDCdaGrAi49HuXF6sIBi8E
6h5aVMsSsdi47sAi/4JCyeX11FmxKEGvWA+4HGHBjVEmef1t2fhHaNXCoXITREl6hxuHfntvHiMz
O/QlT/11FWwuFDhIKq2sSyU+5g71wJW/ijRrBY552x7CgY02Qo7f7VcbkpHoSkd5tjIlnXh265uP
kzDnU1GUCofq1GrYwu9bpEYHfAbEk7cceyGzd1Y5tVTpUbWxnkGY3VpBqbfPk57/D0JQdM92qp7E
uG2IaGPskQST+B/+CUpFIY0k+P/FKp31YPK4NhRm1ykGTtsaNojFOknUdprNUx8+dNlX6X7JhaNE
aB4eb7+NqyZJuYwFH2RL39BD18sU44p71kW8Vlw5eaEC8u0hs1SfAMvE1wjOWgYmj8rfyry0UBnu
isoi7pMjg2kQz+ogbO6Cs9TrL12mJvM8JZHaMKnQEeJCHZ+heXUOehPgg4HUWzNW8aBopVrxHX15
+06Ogv7mvA+bHixCAK36pe8PWyYaLE+DYEOmL8S1AUNhoKyGsYIL489epRSnSrie5v0cbuySXsTs
OWDhrjiNWafdXiaE4itDXjBwp3mGKwSOuL8KxxOy8G7y6GRfHVfuqWvfVY9imDPlapXb/9TwLmZz
SNZ8R/HtL/ZX85R/WuYu7PIRpaRNpuPrSAwZSEjrP9h6ad+5/fS44KwEUGgZSCZFzRn2gAl0WJEG
QUkEMUvLd6cP/wSYHXHleFj8gPFNL8EGZ0vF0wOgty4Q76JjpWqMhxBKQic2SYnmWYxkp/fP/7yE
RyBFfrouBW7kV6zWD3QXXc581nTYhirHD/QAVUJlRebQAN9pZapiOLRGQNeQlZTBfjz+udYo+5ck
BeX1ElHBLl3H1ehimjnJWS+UDcj9m5GYRm/EkrbUdlfe71/Wi0wAfWWbdfJh/GGcATbkRjogmusf
P23RCkUEFWGIdtikau+j1FsIG5YljFg+RsuqC8gAXLEQTMlWAy3WTIazzw+x6Z/V4gcdQ3CdAQaG
Ig2VcyovDh4ySdIaYY+d5aISCurjAgiZzOqWnCqBQDOKBUss0vbG4CntXT5eAA91PJ8wxr8LCSYN
FHCdU+erraezS1BxfGi3MpHqgusLV5BMRWxO+VZA1e9upM72aSlyKkJb9ZIRes/nt972G9IXXSev
0G7/1waZ0OCEk2UiCmbYADzyb5FGwCZcTjP5OxCsYpNxfLtX2jqPaY9gNpKBb1yWXqlxUtb0FMU+
HZNF3IvB9FaD5o4GQFjlSc7OrNbxhzRRIeUgC4GyrENl7k23h664UJMkjPhV5bPcvO7X7RyOb1/K
/4OiSkVXnhOvU2e7T/hEnhfy+trUgo+AkMXRrGbxyRV7lbJxbfqHQXgPVe3NgqXx2FdLkYqKte/H
0BYI5nRN8wN+8uHBFZV84jSTOskQc3Rc8h2MrfsBB+KcFnGc6Rykk7lvN86IlfjXinnCFxrOSHHe
s9y1nHxX45TWdIKx2FYLhdrrDxej+aUl3Zz8p+yfTAjUSwqhvTCDI86tdyfjgPco70vI9C0qV0SD
MeZqa82zLm8orBruC1cLP7JjDl8Q19f7jKVtUjBH3j5C6vxuK1OsQSldIwhy8yyzNmh3bHvz0xb4
5kn5yaTa5VEs3eFkjcVEdopoBc7Hsv09o12Xs5O8HotHR706L0OR8hn7WWh3Ue4S0M6nz3wIRaaw
997JeAm1kYj/N+bJTAdvaDb/usvHOgxk8CfU6hix1i/uCcQnY9r7kkQi36t/JteoTcfb4o8wMaJe
VYyn4kqjqwlKlNiksL6gUcAiTeFxQUQWXnU/sVYhb/nrU4K6HIGx4QvOJcVBn8dEqg9qoTvTO6qe
pEu3mruc1NMtM7WLG+vf1tAU4+m3MDjLKxQQbWIp3VrmeUBebvRKrjdx5hZmhJRfwIfREVV9GJ5d
DU1DJt6R7NJpCqqm9pKOEIL40jBjQH+WrlLjwdFZUcI98b1Rp5le/DueLBX1B+IpsiNMbae1rpRZ
Ew2qBchvCnYZNRSqqsSwUzJAw04kI6+rCR0MdpbN9H2CZNcY++C/6qmu5465YknX5Vl/8NiYiV83
q7EfGVZHxkAPDqYQDSf2KYFC4+rrD5nOtUgVcmJTRc/GQakeIhkAyIb930Pd10LzTBUb67n3xQSX
MEM09DEBIfjxk4QfojTHS+KR2FcqsxpSfZWJ+UkvVvCSaLiiwVWidePKbRUJJPlMngLxJtKyJB8L
X0wHHO377kP0otgClipt+pUKgMtzULgVNH4wYnNktDNBBAdHxnPE0oQF//udhqgyfZUfz6/+PM2I
9B5eL9hzaKPaJrEnspyAr1r9KRXb/9EEHDnZP6WG3ziJZDzVTPFkRsjxNcTr0m+pnnw5F/x/sKZf
ObrsFGIQhm+CiySlV/ESwefh8rPVTnUajIhWvXXP1wSIA5ViW3Bw1DjoIGC5y7rm9ZFT1U0Yvme3
2EPJ8PmljxqQ7iT4qMvc8V62/W2OJgIGjsisFPvKKgJAIAgbapKWYmc8/AqaRDhXy6dlrnil2uS2
mdNqV6FMmnbCqW2ArWP3Oe0ngZWQgb0K53Vq2nUmq9iyvgCx5HwFa1zkwBZQgikWKR9KaNryW1Mp
ElwSIYD+QiFgTXSpV215WBEMFL5fgOr7xcLzw5OwpqFEw/YnDqQmbRZ5I7srcHWyWBuCzwRBg11a
+LgOaWimBXKygkleDNSDO7Vq6Wx83i5mhcPZHTObCj5nGWBANxfzSVtOFhIIBDK2IqxQXinQreBt
Rd4fMo3ERK6v4tr27AuCgoArDsjw9ne48RXZ6n9/g17aARZAcHHSX9Hwjry/IKojTzm2gq04jnnm
fK6MhAZsJOfeqF9p0mmkfIbobs8BsS90E7iGcde10SnwsHaR2LwKmFy3zDB1fUAbSGGbj9J4kdhT
FBiz5KxetIV/WDT5yV/tzvZlCJXUk/1HD64brOuxcKujJooIxD6Coj1oPvOuJT6xefnnyi7pZDm8
ivHHfWBwLKP00qsbPfD9ueCo+ngjhYBA29qZpfr4Q/3IRGVbPJZcIqtZMec3QuCRAm7kPROK5eJk
XqIoM1fuo7d9OhzPIIz8dVu5yE4YIMUbyaPHD3/Fuf1JGitL49GwncJDsOFNj9DCJscvZPbbU5EN
qEeX4t5usBDdc3e0rFW1a4DZZjuSf0F5tgJxxCnRG7UwCt1l9lyOx6rGQzwPkA2tLBOa8lDt54Ra
R9vTW/di4ySz6oCCF77qej3oUfIWD7zwthsGN77zj30b/jbvn3pMeyN3W6rJyTV8bCyakS1fr+NJ
3/PL+TZeL12MputN1kBWerYpMwvH8wToChreMX8Rld7r2S2kJf62Y8f9/HA4kgON080yhXuq+3UR
piAWAGQ/HTwl7piDtq39IaSDWXhSwDo7B5M+mwQJJtGwNF6qTXd4L/g5OriX+3DaZnmMhyBTFTQS
+JsG9K7TNrHRg8AHpfiF4N/Q6/ZIZxEI6cRRHcIr9pPtE2NQ1i/SPol0R5K0nJf3EZ5YNSqvt616
/xRpc4NK8qqPIhu9T7Hn72u0KifTfY8LqP4ovuIdPMTVKMGj4yp/8ARLcqQkE4GdMUB862sXXXzn
UyDLmm1x30KuFz509P5m+gw7wOvtpSb0GuPnVQrX2m1RtGRZ+ZiEIT5mfNJnjwDVMSqwhuSVnkc6
25sgI4nzlxNtULp/gVkcolhRk7rqXBEjveWV5WVRLh3NSbBmous/y4ISTFxRk2ewtZPx34c3FHjm
p394QGuf9tTy8iDm8N2y+VyfzVIIUGdgF3/TFYCcvW+8dWbmhPP4gA9vKReqRO8nOOD+jYw2y9ng
GEiPsq9ynOCOo767WQ2f6Ckn6KcRULKbRo97j3gH0qMZX1bDhqLC1Rn+Qyz4jbo7NacFC5mWhNxL
9rZ0T6GfFIVQgi0jqBqK9RtQM1AtDIAkNLT1fO6FeXCiRgIOTVBM7JMZaJSiBJ9tT1Yn3Xmv+ayQ
TV5aajeqrPGLw62yKj4tixjlpyB7yl13Hy/7B+q08Sc/eo/b3y1rMP2jDNF4Q8S55fwyD0dtB//r
VecNaFBNzGEkC98cg6VAhdEZIE1x712ho0QZFxv+3+vr41y5Z5MY/QwZzfCmrVjj0HrIGe3ZbUN7
7aBJS4bP18GpGF7rFlr4rLd7ngqJ93vd2B5lsCTpsSHFyZU1YvQ2qMQO8/5e7ZMNgA6AMQtDlQF1
6Kor3xEp/OB3of9emsa0x75EdbpX3SwqUMa4EZ5AxbwjW4V0V4OJq8KtrVAUcfNTBwIVlDjJ66Ik
NEODVNlDWtNl44SeeEc1u31Lo4703PLhlJ/IIV6qG1Wp8/UXiHpgpv7utoGqzbOaIMVoYXPw1tal
p6yqiTC8YaE3BsbM72dPePjBie8uDYfZmjJUoZZXj63Cy8SqDm/EZ6/TGBDV/lPAjiINf6vaQu3V
sd04aMYPiMAsITMwTiDAKjNqH31w4ijzxeQFaD2NDwLWLKdPBS6t+vLaGSPbi5rRpBX6ZFmY40Lt
JmxxGFHSKHAwLgWGar8vGpdp/4guP27QCKy12P1dwJXRG2SsCVkg42l2/DEsiuchdQttF9nS/8sQ
pbwBTSJxVoJxPGC/t2q5YjN42O1CKmYaD8IVuS04UY7hLckcU56Q5wlpn6NegON5fZw2A3KOVKR4
T3Oqr4x7UwPa+Zkgi+kLi1T8Dbj4JZw8P7CMOcGZTIVSTV8Cp9/0fG2YKSjnelaL7Lgn6Sc6oxPO
eHP2wF7ND+3htIUkVynZuWH2e6/GP7Uxa9zhrzM3MtPnxb6Ni9LRDv6kP7moCnqexQIntgkgVFkG
F4GgDM9ydw9vTNk6Iet8EaAAs4/CsbHgWZRzyDbMS1je58TqHQtUeJmoZRW7JHLdz8GimFJLtt13
PK8/eiwkIFK3PcCoAGsZsgfruvJT94ia+X03n3J2NL6aq6RInJj8+pW2oJCe3Fvnkt3mp/o/DWZG
KIHAyLlEV7TAtknZuaUM839yin0ihR76jtXK3HVblhYSdS/Rfiy27rpSqWMDrp4k1IoRxvUWw/6v
3f+9MM+8TE1HpI81N9PxgGR6v3RZm940LJMp4+S5ICXv7P2DGPCdppEWsHZ/Ni/DEaxv+csuB1+I
zC4jfFSirX71zXL3dxP0yophGZop3zqgcsAXPPPMwakPJBOt752DlDHI7UQawnUgglGbgdmoSOms
23eVX1bUgH5F6zRB0pi+18qyeyggsexkIKaIaa7+F0NO9ZF27DVThbAITOCxtjY2uzwXSJSZN+yT
oV6IYE8vQyS0kc+QOt0vjjn0Fq8ITrfnbz7gPzevXm6tyGNTkttPrE8QtJcUY2nqk+qAA4JiPWcv
BlpNEsV9e2GxKwyxvkQqJWXi8S/JXxR7vkK7ehyUYzvcumKZA+wKtGjnGl+MrIgX2/XCJZ+OV4Pj
9RvUzHUfCvM4c4Gfjzt4sOOevGjIh/u0Vvwy7u8AG3QlBDpd8bc5LcnlJfu4VOfEQoq2wQwH6rnE
ny3OBc+d6jaXX6Br+BRSC+xOYuJAYqFztFvK+snztLaZi7blVya+EyizY2znd4G//2oJgv5QY/H+
Ukh6vJKdUcp6ZSrLosQwf9oKHQkt0ed16fO9CGdGdS34yJ77NzLCqOZhsVEkdQgK5oy76dAZuPcj
kvNo2UdbRYsFlZu6lyQ0TwTYP621Cer4dItjEccTRa8bQcie3tSadxMDiVCjXiqBJxmcLZ1+QTPO
Uzjsifr19g+a6y+f0xVx6WrsPB4waxBvXuFucAbH2bZ8ynxoyp6AMdLXI00rDIRF1QDWvZ1TYbIh
8x3aayOieJj1ptorEnqc4mTgChhZPPdKUiSwEVljHN1d+HBwTFgr66jTVwuk7iKz86+z9xJCNc9A
dOh0I7e6kIAN/u/0BzFSuqY7Wy75ZPUkpHHvACb0UvMB1zj1l/rC7QC6dJUrxFMZZne7ATwmaukr
pLoyuVjwbpfHhfNK0HvRtpIfco8X/M5LpxmBxzsgFBJyb8CfO3BmHTwv4eqRifkYdOEgwuf/XJNm
1BLsD8MZqjzb00Jr/7N/cvvxLjQ5RVYi1cCLpSlo8VcltoIqRgjpXAwVPOXkpeE8KXoVvnqiKU7K
D7DJv5tr/PLot/7obmQlLy964U+/DG0sz4UT/oOcJR/PbH4b0UOKWfb/B8u6Z8PRY5Cb3FxjyCfF
CUL43wlX1mZYAd759eUV4cFjequxeUsbORGOf5rEHZdrrWlUk2CmH0RlE9MnjSaPMIfY1FHb1TZz
lFE+1RlVaP4Q8cuWe+K39kh8inHraRB79MT4BuOqKQ8sP47IOsqrGdmMXowxpshp/be/gEpE2Z7y
PPI0t3KxlYmYnDZimY0bmQBegifLv8UhvfTakGkVtcyBzu25OuDUVv8rm/6KUP6zghjqNQzNIJs3
eY+3O4ZHLWsbeLHp+RN1Ul5ErqkZQfg3/cGJgwtt2UhVgGo2nd4yNN98mf8tjeMq/fs7A/Dfqjlb
i5+3LOJ6I6bJxILFwyvn27Wv/zFKoZwTve+ZieL/S28GWuJ1OuX6ZaHrJl4efnLal8ISG5afOJgV
RtNqJ1VOKK/yX54fo/+PEgEXSxL3FqrXJZo7I7VM3CwuexImGkpOAJRMLUcrqfEN3wLvtctDbExz
OR6fV74CsIam31cnkmOzg0yK07NYahh0pAlUsT+gvL7s3fx5FiJtd0wDh/a78qqNa1KoFYAmE8Fz
kFT+W7CjnfhmX189LcSfh68s0XI36PWfaeo2eFkignhhaXC+wj6TxNcboGZokSY7efQbtqS2dJ7c
qwEOngKFJN3TfkAA4NKY7eEvyQMNXa3hfe0FtCJAtnEusoTxzLmDeIx+fFzLy60V5yAlF01FxVQP
J+Iywtvb984n+zGDXSukskWe5e24JIBH1cdvp+DDi0hknxeiiYeBBS5eUP1o3WgCI3hPcpW3DGfQ
kyYkUOIUFVaiuOpvUEMnSJb8NCb8WO6xZhaC3X+GmewEDu7c0G/yh4ezZO53pFh3GF3MuSRX1sp1
ZkGXmO+84dGy5PTZ034uSFwwmMaZPXm/HrnJzusouemX1EIScPN3ckx5X4hHiKgfKntz+xUhL36e
p6xeZeWjdJgFcIMqZr5q12FYz4+q+mrPuNZVpH7I5CqM7DUBuDCvIusTrTtLI0XIYoiiyChkw2ru
hvouEld+WrHHXwjN9wQ6vR+o3yE8+Vg+14C1JJfelgl2wPFPwYEONcab1ZDApKnotggIejiOX/QL
YUc1m/UBD5m7xxKEG/96bfl19ptHyL81FK2/gFkmgOl9LYNSeDCCzeh2QYwXcn7D8KeGH+AMl781
BVxm7p3oYKC21eL5DpdE6EdoyLKRMvrFmIwslIzXDrMuVDrSdyiSvrlLyl3nph05f2qlYXzlzvqF
0Roh0q53RbnklAvyQAx6GBn+Hv7hMCixZUabaSRJw6Zq8EQs39MgrKUBTbGg8npH1ga0fQcF1Uu8
S09iCqNHgKPZ+DUuudop7zeEyNbjI0Y4zRRs5B8kdbqlGFt8ry/ehkDFGEC1lOvbpTcfjzjmqO1r
m36Tq3OGpXUuTDIS6n1LdLjyHcByqysbWvbvyCucgBK+5ZFYReb3DxSCI6S9RYC0oBo5Lr/wd5tG
om5gTlLbGE2dUCDCU1pgRif3aB+K1ZcG/f1oBlbGJ1J+Gtt5HQWQiYfa0JRM/AWsKHcnwwB+tkMJ
vJQiexpGHv/2okJaRMPXve8bC7frLLaWjW22huFWlMC2Lpg6duSSB3hnNHKAu50tSnBgNWWfnNFf
ckCGZaSg7OvFeDQwOhSwQvCkzMXDdEiR6NIhwhwbuqO59T87uaNI8OHTx1Xnrpq8sfEx0ulXMKuQ
Ie01a4aHdQdhQTSW+O0l9h2JVSmpK9COimeoxENV/orCeFTRQi728Q3kEf4Xf5RfS3fjOda/skdq
d+I54JBZoBEjpOx2xTLzOYKvdxa6XBBT48DxWgwqFH+8qnjVHEB3T0qHveptgYDMJhL5GZpm44Vi
I7rURmvumzA8cYg7jG6EZwlOcgfxNYWGjJ6cKirzUWnIv56F8JmnDNEv3l3s/gW8aBa753psud0Y
wMhuGnsG0o8ZEG/xKsRC5zW9EZzIIvFPr3fSmJJm9HkteUhFG/H0v5jiqls8bbxqeJCbZ0g1P19f
5CRrulqhP+mMIG6w1q9yz84/VoeCfyCmHOZMxRwNmFrjdaGlfhZKGA/2g28B7WERf6Cc6PIS8ck+
pfgFTAiKwFF41MHejs9KvWcCrX4OQb3xoQeNZUEpqz53C30nk3bRNFOsj51cdiwH4JMawKxFm49s
R8qrKnUm6VYWudUvf0CExfMvE2hgcC/9v2pVtTd1/WuCMdtiHkUv9m7WqUkDk9t4tuQw+WRgcafx
G7rGCpHCnAKLzaVw6wq96Hb4qYzYhOm+BSZjLx/Aqs8XKuIk6TThnLFH4lsaNAY6lsvF4CAiXNU2
xYiS0H1W17GlI/nJiR+A98IlIMJb3rZGhsg7hWHy+pC54m7x8TusMsEdM08YQNXPWT3Tn7gStxS7
XE38ML8P5Q1bJ+j0UPGZ7aurRQbbnb6RIzPi67f5smLLOtJ42Fp+4fuL03Wv+ResK7zlzMSC2gas
QqXxgphWX9RT29dGZ636CTSgMQrGMJg1ULGhFAHqb6lk4niN7XmZVsDbfRchpBDPxN3bm4vljRER
QTKSUkEn0qA+xM+6lDh/+hywflrV0g7qyveqO0eCZ8h5pKHrTaJrdb4jdQOqCNfSmKSR6izmsnLn
eguQXEJDEQ9iJ9jJ5/bc5XMsBjvFo10O/KTkgQT6xvwNJb1i7Z7wqUoptXc3kDc2ItbERLrofpo+
bgYL2/zJONq/odObQ5t3elca3btzpO0T+h2+Qq+KGdiyGZ8jA2RD/V86tTTQuBL5YyvV3bjdrnFA
NknGmacnE2jDzPH4URpCSgmJlqHw5aIGRSdB2v+2xFDeBSARlVYNDwNekaQM6LlZgHIXBiME5hb5
v4lnbJZxl1Rp3MzHMmy48k85QDWUsApJ31wrAGCbfBEOH1tQJvxHobEE/8LPGL7bcE5cLzA+NyiP
uLLTbCJOsudAUr0RKXv03BOy6lsZGKtl/Eug2XbA0APnTpPPNsLVA7m4yRgc7Zy7FsPvtr8IEzDh
rf14zws5nZbLSHp6J8P3DyCKHJUiScasY8oAGcdXJ01GGRfJTzZoJoNLfCG0YydWwOHWivnxtbc0
2K+jGGL4aG62JGq6RBHfO1At8p/ZZc3cIHlrZVS7RYDEqjoxu9W8JjNktBoI6Hp4IK3b32jrin71
4tvimNnD0xqElo2lxgfMbfsHkW/JeG2hStSxjRH1NXc/AjvLDWJ1Jjd18mlgq0xlBUSI8Qjh6GPA
QJnNqMTXndkUkepnbG8DxPPD8SaNm6cfIFSUTzuVHQrHbkrtaztmuMeKlPjLHsa7woJJE8Qhb5mJ
pN6blAunomZjMaY0lAnrdG9JTc4+mnDG7kNr6CeRx3Awa92aZoHu+qo2q+CF3ot3oy70eaj2AHe1
qg6TKHBEv2/M7ZWU356rgqUURqi7NAnlV5dOgTsI/3EYmbqWf09JByUT/7BSK49TM4nAvAOpqHSo
Fbf3SH5Xg80AZU/3fGlRGz9t9UzSqa2yAc6Z6FAtu2gYiu190x8N/27CwWNqD1FZLhF6+Wv880Lz
LQQ92wgsLL2f255npXcdiMNkPxQMBxtXQqfxRf3gYc+hIaRp9vAEe6NO36OcdiQCtTEniBP7HsGH
X+Fhc9RJgCvNTDwvwhTrEwN04uImU1VyivaF8MvmoENiQS3qknHD1FmeabLKvPtr4EXV/99/bpHH
bz2Nhkz0X/fvN6T+jl1vFKEsK0oZz9JJAJV9CMCw+oCyyKh8QFBsnKwut79PxLuiqpWzREPnmvZz
TJT+et7aup0tXjtZ8tnza5gxTKd25U6HB4vN3Bd6PhImEGYFfykKPW7zlKIfyTnubHk5kkEQ5Abm
OveFW6Nc+0BbFg0RJCRlEpPYjVke9Fm7A8InjhhsuExSaxutIWsgNv8cneeEp7ZmNPzPXqJhINQW
b0QwpnfPz92vEVfjONgPlKZdI+ogOohHYboQmvKQtOUk2r/iueZLYNbk1m9splPv+WEQF2ZjcCiZ
swWlTz6DGnc/anUWq8ygZhFi8q41HnKGdI6BJSDX2Qv2BSZzZhq1r+XEDDqCkFJhuqXtPLwLcu9V
7nafqJKqrtjDXf0F22QHZty0piMRgfEhk/JnhJ8hRmc0gMEkYNytfqL9RiKDOVggzzYN4+89tH7V
WDXiL02dsbxxg/9osvQGhdbiq+eo0paGs36aV7WbVFAw+NBfk9/LhY5EBnLiIdvadaha3JDiB0Ql
Kp9uc119dcmRPPYXJsBIgNmDiNjb0XJK3dT/53G+H25GPA5bzrQPlRIvAFJyWfR67vgwKh1iWUCB
SCv+d82hQwZIWAt72rNip4PVMj6qzq3oy8Uon3bIjle7BRLtjYAhH4Cq3G4rYjbebHWlU91kZI/J
chb4plgYXmwGjMqJOI3Ps08AHQO6vNvcxieUffKY688PIXmxqEnaKePO5gyTbTipKPyqLpw44+Cx
SF7OcWif3UXm/VC0pqj6CR/o6e8pvcAJao3qZvaSPtn7x/zNMSM0QsnmUz4daROpdpNNlkg+8z5y
etsC+FZwERxlYWZtEa52ixcY4/rhG1k8IirpXF2cGRrZar4bRFongzbUS88oRIiBfkDdO7Kt9pp4
o2XywNy1u9XfQO3gaB+Ar6wFwj8qbH9Zg3X3Y2E/HJz/tfwMSYAW4KWoosp6qs8IHa2y2RUyTxpR
34dNxULWX5hZmOHhF8GQm/wIzUQcM/MUEm0y3gvsG/CxFQnqE7i1NSw7S6w6x7EVLlo/VIet8VUu
bBtvmGyYtmjSevCB591sMIAfIqQJuAL81w12aS4SzTlrshkC1gLz+49932w6jaWxkYBBqPMLwyFS
a+0wezauoaQb/LC1xbD7wSjA85JlCV7Jx2D+G5pP7UhSOKESmRocSUxsxd43akCIddpaHK8AXLCS
5g2c647CUXxvfAmEMJ1O6xbNlTCMK2abZCG0WsTKyHX33o02vDLXZUmr7+CikMBUWMa3H20pvGtf
IvoYvSv09Ys253IOqTAv71hOPgUO0EbCtDXPB5GuB6Fizdm0TsZrgcajm6f/cM2WLvddne5ShfQD
emgYFK97IUj4hCMHcZ+eu8jjn1TpUsE71KHdUBx3N6FP13tPCGPjIzMYqc6BET8ZsikrDo8tm4hD
D8hrDBzX2o26p3jF8obQVIpiCfKaeyfCzBjYPa900P0QaabHLL8rMalrhTl2Y6NeVAl6tSUVqnb9
fSr7kUhiaJn40m+oVuQCpgHySaEv5vk0fqb+jknvLXhrc8blX6uG/srmzsXFV8rJw3Wl6hv3BkJ/
h1DLKH0eqo+bJhu+JuF6Wj/CHyS+RkB8+V44yCS0HezAEYXE0vnGH5SbECj+4AASzN/OPRZmliMt
UBH6YtgxFrZ+y1LhGg96X+n4Ukg71nZff8y7Q5TAJ3o0bLqa4blPHL4DdJnvYUSLeuhbx7TCSL4B
wIaiQQ4VFGoNGRim68vKTVCNWTgTB4RIftdAekNZAmoDvFY/22A9wLbHXJVpwjzHC4Br5+EnDRSc
rDYz7zU2QZGzZWC5CVWW/az5JP/LH/UPPtOHBCDHHPO1HJc33xgKJrPh0sYT0vzvjdxprVFQE4Ql
C9r5ygUGKiXDP/iNyHqxEUMYQ+pV97Pis6DccJksn6s9IH9eQYy7Kvtqdk2O7N5D8EYv28sYxhCU
AQOJu3CVEYuEAUWtTS4KV+PbaouFJEId6Uc8jKzNjuC8lGhYoDp7RkAeEWDl7QyIQOzlQDhO86wH
RNOzjs8gVmwyGYXH5Av+65kDcKbJ4yeDxq3mxd5g6WTHNSu+1oYzWpNYWwaY+9T6EaATJ8UsENki
KZ6DvTq7F3+ubkVemDReg5q38teNj5d1BfNcTGSwVLZdGAs7me+wutybBwSTYcr0CYgCRLeMe4Ne
ZuPFdkEZnHUKuJgXdhmiU2iBWuzHs5iepblzxwMRv1LTMMetSDM+mgNWuia5hq6PpIS6eCRzBZ0A
PAKOKujFOxnI2ICFcQ5bz+TjoiKI07INvyLQ+08gUMeMOX7bco6XqdTjjmTuElPFW9XhGN+pEQpX
So/xaF62rE2cY9w/+7On3R4QAQyqzIomXNhKwrfRKNgU3XXwTaYHx1a78OwdCtNzpNfC8fm2I0B7
Fpqun7vtgj/Y/nKqwW70q8ykr97menEmwXTHvuDuSQTy2VvIbIsnlSWHNwRVZLAoNI17ng9E2Zab
3MOlFxT8BKE0HO4bXwthEHMZVk88Vxkg9x+7taIEQqTfQFz1NQ5Bv6pRqouJb0WTFtP7KXwHpJ6P
za780+b/Rm5qfdSMP+jHVJoxBi0UCKSi6OPYWHQ21X89jsZF9S0J/AcyhaGdC9dTxXmXV6KWcDUi
+I/wxNmYmkj1NCOaGAq5UH/205scl/e8B2dqafppq6IYdqhPVynvuCPPju02kOkNBSjTAT5p9XZW
x2dnGmHuAW+f+UMZJwr+er9COa7H9NVEKEH8RCmT8nN4UhUCqkcqYNFbHP4qaivBJWYNj+ZabV8T
JZOHRR0xeD9C63VoNxNa9wz3MWAe6P5MyAeOfRh/JEcJ5tCz2vZdfD9bYR+p/AnRfOKOvM+YDvwS
+bWX/lHQOYbieePWzehT9GomfSWWoySpbhBP4avR8ss4IsbQyc1eyFwTbxEBpY/RI9uW1LT49Puj
Whu9d+TJVWNGFHtAsaTgaEearRGMURGGPI2I54hPWHwSvhk8u6kgzU1djONvhv2m8/7S0f2uQ8oA
WquwVpF2hZ4FvtN/UoBUyp5YsW/cFb1mpz+eZUGYznkuNknhlOw0l/UhuXqxaGcE3zuOVVtJfU7c
O5u4pzf086eCoYYDcC60Loiw9OYX6IMaSD4p+WT1+fZVgsctwPCAx8EjOCxRBOBSZJpGMi78y7my
A/wMjnHyv5uGP4KmeNmUDodOk/7BuhifeRZ0CiN6uNAK5yfS6S92K2OXeTqKOSFqjYnL5SvV3Q31
WFOmJfiVQgnhxE4wY5nlmoLyWvkw1Dz3QOdBlQBW5k9UeIA7Eec0T500c5WUdITwrwPrreXzEhAa
55R9doav0pJFIRbIb7wuRspgDwivlXyv+k7VmU69kpmuGErH3Z437a4cVzSu3fhqQkV6wivALpSy
+yX0dJ7lW5k0R1qfJMYyaJbfY2zy2/jRAJ1ScPHX+qX+K4TR4bWahFUcYZ+JDDNCueSRezxUu2+t
1R1veD29pSipZq8du3KFXvMZtjDoxwA12VOasb/0PmdJF0RVdOgKizEaVkiP6PGBK8OSbux7eKA6
rMDNT0QogGeQhFB72acpFK/l1dccMw70SshAxt/CWBNP9HyKK3dUerpA/0eK1Xaudj1pitmG/FIB
74/8OZBl7LWSclXFkRVcdI7VOmTMZnucnEHY3A3TU005gewU4SMHpNzm89+16PFGI0yEgKYnHCrO
wg0jXIXd5Kuus7Cf5asVxGoNAKr7+RmkFXPUariyVJdP1xka0FUpxZY+pF+QK+UOSXgTIeUEzxBQ
1AbAiwHp/QO3/DoaOGaI0TGjTUu68yYxsXQHMBbgqmnLfRYz+RFqF5pNXAXAabZjX1HhzWOPXxrt
iQoPgO7rXtU6GTPexjG1HuUM+9Yso2bDDQYcniaFEoa3+zQgOSDLmorHfz+bP3VOm2Oj68srDxhr
udigDKpJtzxOe0uxo/6PrCH1BOlN4gfZ6Xdd0iYsPabDQ++u+7xpp1JgsRfRKe3sl20dwwVAS6lC
q38cVRkkCXHUZUo8cHwe9LdNqFVmP5J4XVEPzfZNbGS0DvlWZkx3Vf9eyMs17LDushk3cESR0Bo5
CwgBqnomymptifFiRqLEdIVbzM5s+oZc/KZCq5YHhCOFtWGABxCCTYVFTowDc+tfZlUh/8/me+pI
9oqZ1EDCmRv/FkfHr5LbOG8VaA8fNKrU0ndLaX+J+TLy4HO38whhbBtDn7g+P8x7DHEiYiH2XanK
ea4sG7WHb22ZeCVqaXGbqF2iJokfF0DaaOyFvTB4UuqR5oAYrHq8/Mh6xHDIfSPYi/sDVXmgdfP4
IDA/9y70mEuCeF0q3UmhpO3oK83vgShUMusmqIGEnpJQLlolTLjIVTUTDleSpHlRlLCj4u8EWSyo
Sv668s4AGDrSEddyRe/x86bOvy9Y82nj201SS8m40hBTQBBBb29mY2Oz4CJh0I1ciwPwQQxMgmIO
8B2a5NRjsH4Jawf/o3JgZ72ECBdBPCdlsMPdNB+642sP9NHOdFl6qnzfnlkq0Kd69jGfPviLw00Y
i/Z+VNogoXNhjFu+eDlxTmbTzsvWjpc7H+4v0JxiLUyYjcFC2EIfd5PkvoSUYCciY6zBf5x8XKdl
bQA2GXbD48dJRlh91Qa53deC81HVw0vlS6+zNcgC0vDHs70nAyBA6fKOv7szfaKx6Pk6mFCnDQbf
gBnIEK59v8Jhe0MCLJCa0iMcIyLwPcz0xJ26skJyJ8yImXlQG09Fa1DmTCH+N0o/4WsDO0Tzw+ZJ
cY8Phd6m780+J8pD+Jwk/v5TgEpROXKuxttf1ZJCUVmLa5qShZDONOS2KGca3ay/k+5T+LsVvF8I
vMwSMmkAFrJ1HRr9yRQq7uLS/K2bSNhrd9X0CJ0XdMA1SoGgut9/W+83J1tP0B7en2Qpo0CAr2pC
RL4wxT3c7KTe01T3+2wfTtBmxNllGYvcnu8Yrb+7bhX3qmj6aL3OxBlCn/FOfitve1t4evKiOQMR
RL0PXN+3k7ARynrc9RKhxKwSv69/PkgjQ6+VT1Bkm0fOEN2KXcHdP3RcnFh0qFf7T3iz3Y9L9b3E
TSfEkPaPkWnodcz5phEXjTfKFV+9VkRQCf9Mavxrkm363jkIXjGFdQmRh7PMpH9hFMLZq3n6fqrR
ayS+Jsp2eeM9DA3qZuqqr1t01nQZ1pcGETiO8ixIo6QSYQQqrVLmTD/0eqUPS4M1SXfzpP14th44
CBd7oTObNp0EZocWPTHnvoaoVbaozvZH3fk2JEYoT8GiJjGOxt73f/vHOL7ngfRVABFcZ2HXcViv
ghrlpTzamOkqfnt9RiMenw0Inq4g4VZseYb+R0Z3mRkrfNn2F+P74gismWFa0UPgn5QsFZHRHd8r
n0uO+viAGKTvNh/Ej295h+/+nPORrJOAGDHW3+23lb6ADAg1qQT2iLKsHvCt1XkVvQ6hFOazxGAF
mshIg0O2aYk+INs4kcXJ9Ymq5s3VoY/Zqq4Lhd2G0zxMySkUFAJgxGQiMFylH8R2StPg0dN1SyI2
sfibnV3zAMZLxa1VGFbnPhGbs/NGrvCwyBZdODKky0amBntLiq0CT1o5j1K10EsDP19/ABEwmzid
UkTNjuANpcvEBAS2YE6jNoz0M57ja0nA/CezKwt5Yz2mDN1IwXOAJUtUeBs3AuZougLiEDopCOuJ
G23lbAdHcal3S0fPMQRn/pjuWmIVYv6og92xGT1h+0ypBqffSrbkTlHlAEnutH45K+IwAns3u0Tf
CG2sTRz7s3vUqMe3yYE/O4iDBR+p6kaDtFnhaj0OF5lcpowhtCmCH6uBzt3YqSJyJRKlHkgAlvQZ
E0LSBf42VZa140iiEtUt4X/l1aabhgGeUXd0wKdZtZOpaylt7/ezLjwc7k4cfDg+JNmSRYyaDl3e
vLTMoa6Ubz/6M9gRr7lSZ4TWX4x/yNJ2RV3/W/cbrNlFi1aJbmQYkH5HPnV/FvXddfBESezl9C6v
VSmqS5txDHoMQYW2OYI2kAWEA0edQvKbfsTX3XqnISX9HRU26zgmB3s6Q7B5hKpB4N6Y4Bs67Dan
Z1OomNRSHU3YhsuvQeIUOG49GZEsAiTM/cnRvTU0gQYxHN6S6c1wVn6hGMncVINE+kmE0qGdzMuA
teN0Z86zxqwvOfebi6fWtjEC1YfOODrda36sdGFiG8Yxdeuzcq9/+MTyr+NRSdOEHbHmLJPd215a
hxqOEUC5/u5C1Eymk7CxKsFt34/DkD5/i/HU4ecf7rG3sP5qHv0ez4hvRPLSj31hSskpFBtOy6yV
bOPJ1+NTZH1Ia26C8q6suPhjZZAgF7axA9h3V8DKrKbaq0kfC9NlTXyKL7fPJynohX0QHpr3JMcn
r+5NhHjaTObu8pOgfqHpz319Y+mqsIKjvk2smpvubFqeyyfOK7Q0rUULCZ9vAMsUObanxk/mwldP
SSAxxx0bK0ECv7bVx7X9JNXYS0qjCyZn64GJ4s2q7Q3rgihQ4F6Jeenu6XnejDDJsFNgF2v6xp5q
vn0es2F1srckM5Ev8549k1utk2L0fT48YZoAFKKIe0N5heY7SqfqZ5veErp3XwR35JJHNoTuB1Vo
v5IpdXaUIFyIdJRDLi/z0Zp581KjGvudvDkxwqFyiNqbF9gb0azb/EgWszjGE1UOXiLrT65wfOMv
pE8bUL14ofHwT3tH6PDetNE9DUgw0J92J2xPODyQxDLZ+7hOIgeO3n3/LGa4Uqw6Xbt4Uq1kDqA0
AIA1625qgVAfUPA2J/dBTV3FVn1b05aiswQMzOFq40Dqr2HhKt1keDqWfieCgIiBSd+LQhKmhrDF
EVU8aXTboPHFkFU/DT50o0EVdTMYO8Km4d73RPydPruh/mZtVh6U6Y6CvI/SDY4drGemHWSYnle+
oUarQRBVzontYWE9oT0t7vxiYZA4mvtmNMhpEjsT0rnAJh6GGThSzlrwKlkYSoGMBmkCU97eO506
aM0Vfcbyqbctj7Dwvd39mDUg12XFo9iEoB2UEH5TYrEzgNxc+2XVUfkyAlqAkByrluyRyl7JaurZ
jDcaKLujQOVDmmfx96+QBbmktASTBgT1hTZj38AkG6kd7o7wOEI9hMTNrmxw3auf15288IjCFCF1
F7/j7btSq+ULdUQ7wYE10hj9zeOSqT0LpcmklWAD0IVdBoTvaZgM0gnBSEaPWUF714RC0dybJW6Z
lNVHaKJgFEFEavyFSawmg4C/+FX/OQ8x/dL66hSBo+5LEWrk/JvdsSUtzj2TtbS/IEZOvHPhN+Ko
gOT+HE0+/0Ag813MF9UqB0P4J1HRZfU5HQ8lwf8EMfpOd/W8pcHozIL8CF3cQiNGkh0SuUcPrFT9
LRGCiKmalpURE2a06hfsL6Ly5Hix4u8M8DZCuyFSbWvzfB6xHEWqWeUBPy2hyXMKbAlNmPIETtrp
XftJkdWW9xQsgaEMiZepw0bfJsYhQGR5nJdfBnj/OH3bRGP1rcZ80XU5kmycpjudrOVBr0T54sO9
l13S55TO/gKfYCygvKGvZpECj7/ZoIM8dH03Zje627z+5oo0DEhPuIJRBf0LMloDKFJTPjSeHrPo
z2g5O8M57tB7LaTW219ZRBeoH2HVDQjzH22xJkZT2dEGm59vJm03mWHSeB7HXLds+UahyWEenPbI
q5ub184UirHhkeucOO6uFRDTjdHN8u7W40U/zzF+FJ8qmOUbZnyGt8uQiUkUrzjmuGc5RKC0iGlm
QSG1uSE5u+13kNwKAomH6EbSjqM30hEytI9FFhE4hXvJYKE4wOYsWBMX10Fl+SFz8lweoQzcjy/o
KH3MSOi3VLYMnvX1l+noh3EKq7PrSkxvY6NoCA40qd9ojBwT4YdLLD4fsZtqeFORULpU/DVBHKNH
4IOI/Obb2IInq3iNGE9lzdduSSqZeGTaFBfJtzV6LHTRATO23FDuNKdoR6wz7mDXLYJ5BXy7Ht8W
mrSC3aBzjU90SQ7pbQuuZH56EsOh0BkOyO1CoSqAAXudjTjTClmgYru0tJZqq8uki93vTUqDEl3u
bclZl32XMOefQTQPYbedu+8FcbuXL5xBP+UCIY9GEJ1WEZxhdIp8iA88l+992fH/o/f0Wd7kIklJ
qXfwBlR1mwT8UcDLvTDF+tB9qlZo8gw53aSFiqKzuJxH9hF9UUNmvbGGSuc1KGYVzZ1PqwhpLAS5
xDrrP7oJFBMc0KeM0XC5GWr3xIHJoNaSILFLskPebNYyy+YeEv+qppAv7vyT0FkQYXB/jviCr5c1
3bSiq10fh6xFXoyvWvFpNq03oIgVibVyCky8wRLzoCY5M05hM1aMGM5ljaY5DJDmPBqCziIaAjUg
mpZgmRfQjSguVCyOEOOfaUiKf/lZHN5vNM+Uneo6ohS/U7DUnstmfhR+y+EqY5WB38FyO23+jdba
5gQ7cSVrcPy1CSqJ2KeJ5EwBuxxocP5CF2mB1q2IEOX49UZsJ4ZHhqx1DswnFjoDlfwPWIiik9tw
Nq/99WpgmlW/i0LtpojdJST/3WYY7gwJV2e27ceFT+dKMEX4XafucSByHmCM4oa7dO2K+D7HoXzu
XXzKHAixbr86XxF4KxBfNMaIFIVNuSgmkAv/75cq
`protect end_protected
