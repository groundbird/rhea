`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B8is8LlVX0+LCsbxL3voE43lzMa0KQgBeS7lJDrURNNUz/IqCNkmA2ztWADeZr2HbmJoMX6Mtz+m
Obh9/uUSug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ffb5YVmQHPZIo42T2PY1G+g6D+nx5Yn94Lvwg5C/wsij8iZ/Eel+r+994r2NKdQIyV8yNwcNoP4U
a0kg7t71xIr3tBX3TNs8LHEPfsbjVsO1Gzc2iV+XHxHpoCBPJ6TYRwYThzdB8otNfFeey3uOy77z
1w9T0wj4ZOyZZps/BDM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EY8p1Ce1StIT+WuH/tY+Tui3ah+Q4MgqdcnipTnkZo7p425BeyN4vLlD40DjhzKBQgdXVanwmOXA
M8atzoBC2/o2hvsTlndi4vz9MpyA/utavwPk+AAz1ez2lBFGZjvxI1ZEjGEutznrEIFhtHYKLXb6
iQcMiebqQXvre3aEv02q5D38xCzKgVkThns5aedPVxBqcAP9z8Kn4FnIPsZ06B0IeHDTeemt5Avh
Q6CniBIlbjWHuXy8TdSLOhTbD30cL/LPGaGyOGkewwl4mKdEDmeFkzQVJ14ELSg/nIP9jr3wgs7B
B4CzV0+pHX9fyFdR++nOCliDZu/bM0S1uoDEOQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RLMf7jDS/qBpFvh0mNzNllnXJOZwD7zb4FQrolHJgrEI5K411vp5emxCd8s5gDRkOg6MnVV3wKTf
SxoANCKXdnm7v9AJtO97AkGKNppOBlLETr3tcvR+lcHlqm+asaead0Jjygf0OCCncmWQR7rvsL19
5k0Rae4m/0j788FaF/Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k5MsFgP9wSYoyqINb1kSR4dSOfmLK3ounILYcX1rNIQzAVw//yWNPYMvPkFRIx7pymu2jcFG6nRK
rKU0G5q920nsfEGDFjxIpzKo9c2niCyF8TUT5vBFWCMBixMMxsdoVs/1ivr7IRlvIwKL7ETgvhVb
sP55eoBiwDMPrq0vKZFFTBNgFAUdYLTCo/rlcyp4bi29DoLPVhtJG5X7s3KxfXiuf3PSni7q1F+k
wfksX5lOk5/rIqJN3+Vb+dqAHSoZcjGqWMb6/acfgy/9rlJO4kMCHgk8YBNM35rGLZ+M3wRZ8kgb
AX1hWr7b0rFklatqfF4mHSLubmhiHWf4hNltOg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16752)
`protect data_block
BAZLpbelQpQBPuZEDB1B65dBWEO8+Fxlru2i5EscHAm7s2IUhS58AD4PLORAswpLBuJhw1J4Gm2S
R6nDFNllCZ6s/QBraJOwbc/LU5wS+0BQhl9Mspc32lZ1oXk0ps0NOQl2XomnzJfs0ZYRuR/ln2yw
oFa9zj30kt19bGHAKmlkRoR5Z+KnkN5AKGA5WB0m035tAFY81Pgr8NwXe/24r4k+l/5VQ9+I6uMO
8+aAb/lZO7yhb5IKOQiYwD8neYIpuhBnb4DBacNgDxubNrwuyyoVJdWBFrS212KH9xQrkSLt7Aqb
5ups94ryyXlkTyqbaeFjtjlsuwXAVw6zAjIbu8jz/Aj7cyTiFad+d05uD7ltoVIhxAN3RUDWc2gy
pqzT19TVpqoLQkg5psmkK/3zHCra8vrpzT5qYWKqcb4bgIOD2CW/Z0vmtuKqH7ni3p83N+daeaCn
LMSwEr6D7QxZBDCQqEqw7wrg4hh4ENHZSGeFmrnoEbipGORkJKqKwFiSsdLmAFlarl8XPelsnKHP
YYF9A9DPmzh2sX7v1q72iwjFyqYdh4AieuQQ1RRkcs4Nc9iGs4MZ4gdazG0uYwIwVsgfOQL4kWHB
cQ/o6Wn49D71U5zGAePmp5N6ri6kQrWhgJcLVX1G9fPJLEmBml1StO+27LGnYeBIQrFOdoOo7vZz
oOJ4DRuNOxgeHPdZcbDWk+N0aPIMRStW1UDNWZVVbsIQg3n4CBD5k9qLfDJcbN5yCK7A69xTaLcK
n/+ZQMGSIxGYAXvE6IiYPPPr0TWeXOCKjsoHalDsRdgxo80TSKf+guqsl8ayOS1GpQxCrekXYNd2
1tL4yeCRtWP3CcOyyy0hFXQt+GFSafAAWXDIaJ/JFTr8SuEg6QFeCnHgqLCIrY/Gt+szBRRJelvx
KZoYqlgYfFIROZWJYUIFJEXQPYq9NHQc8u3MGkBHQWOEKGxVYhWkgC2SCIcML59XTxJzaWe/rY0b
bS8MG2ts1rF/5ZC6LpNqGnUn+83me5xNz4VPrK8Yx9VVkUU7rUBxAhMIO41EyAqmwZPVL0EX+ceP
Q70h5JQwwy+2c1ygfq/f26sckJ9gMzPj0I3QMi7Cre7BYtXka+A4PcRDsYSZx4uFyeI0r1sxmKpN
LJhK3/SILpEk9W93zHyryxvz+k71Xwdow9CpiwEwsIH6CVuw4xpiO/eiDX6Z30951kRU1fleU38A
p84r3ldrVbT1IfG+YqhiYBbk2a8O2pyxXY9rCwbT9Dk2eXU6nCfjHToV/kQiWJwHre0/IDzwiiqy
5XF3oBma56hKWrznKOHb/aSiDgsDh0+1CnG9b9gD4H/Vp8wX9cgltY6Z9N1eJmF1rd+wc4+uOtgT
uHhDIvinUJiXVpgAYctL74bc1dwnXo381ipxeAfGxNjlpL577m1mHWnf5GhSrQDmApvqrCfjYFy5
OFPWNAEOgYmpxGYxWFklFEr6B0/cHL6dkerIDXXprPQgy0e2apVNim8Br4/veRzy+JGmFJAQHvKy
P/ANZBAiyqgQX20B1YaMuTLtlqpNECxNAI4VIv4ArxtM/QuDIAnDfaQ2RvAbLKZcZ5ZhfhOsTnPn
lkFlVU/R9Be4IBlvqromJWMgeiMOstY0M1pEdLR1jy9gtb0P1sb3hZw79rL7zfJ8KD6mFp8/apk7
g2yayBWklUNz5/uQuMRA47Cwt5RFFfFg1j+cdojqv991IVRKkuuOfonzSiPN9P+ne2AcGlc6s3dC
UNY5yRFsk1Xwl8vTkD4Jz2fBJTZG6kJDWQX9YkuKLpl4f9wWuuQt4ORCJmCTxH4ff3cOaOd4Tetn
w5YwLW0IF2NuMuEh5Ybf+2GUAQWbmIT8lHGKPoGJSTbsB+yFx9tO12q/tfJx8nYLMkkCfKg+uFgp
+tb9NkqgMCYeR9YFyPHWiXz+kn67jpD1yQtCpUSti6thFgt1dWW+j8KyYdc5LAW1jwC23x1H7l07
z4qCsVrlQLsXcUjOClcb0OTwjv3ThC9wApBJ4ZCzREvycP3+tTpIwmFLOfxkYKDDq4H1xJaRyrIQ
T6HdTb/HexUonuHDPFfbllzbEtprEkn8IPsL6Jhj5PFq4J59J+VFgcAwsuyO/vNv+cy/6KNnND+F
bo7yabhPuPfCNfgYjfYJ6O9PRIiDtLYl/Z7o9ULqcdsTIpbim5pX/6p0XsC7hi+hMzkfc0/Zddvt
YDWuP3eoVl3CydRy24lyoXr39gu3yQTLNnlw7fDZoBueV4E3CQTaIDheGjz91SxXLViU7GM0ERLj
vjazTXoAzP1bSEtELxkOVk9MYnzt40mEmgTDOki2dMMR7NY55DpA1G2soDE2rX9l+svpukQi+rgK
3DzRrrfWiRMGeQUW9txM/IrBpZDv3ek9x/Yq9Hbno5e9D4iacMeq1Kk9l6u3ohjOmX+DL00U2nsi
nsCA+VeumdpjCKPYse9YydHnf+xF8/iex6IZKuDJIvfbw8yNi/0R9GW5piC5EPJbP5lIrOiJ+L8l
GK6fpCTAmxTl+8yyMD2OJdO2zLLowPdGDOKxSexGSw+BCNXfXRDvi5QfvM6KLEukho6LSXCqNX13
tbL0jP4Bp7d+rDqR3G3AZtZ8Xsxe8PGPuDj82K2jmoX+LE0he/Mk20q6ObsLYvUmQLKmBy5mgovZ
QyMZbphFvSNHkWtrkHhRZb0ZScSSbGYO8tXx5Qdx0ZQM2gzBIZ9NEzVNO5bfx7Ld7lxrL3MKnV2C
TM1UJROlPXCRLqPwOBjySZLhq7FsfXkjW3HYXykftTUfpyG7ojeex8qZsAEA8s+XbVStf82HrHPH
HHgzMGkxJa9rlbEJbf0k9KL3Jn1VuvjrWIWndEPskQp2M9w/CGHNo/9iPK8Sy0nHAzq9MPQCJfTf
PGMQFQEHzQVocorZtqYbsP+wysfQLZefOe6Zdon+VegoNzpts+rCLgRYvjY/h35RS/ybPiwHZQXe
5vafd0O6ugGel+7V/VlQFeXdWAtN9G4uiEcg8E9oWjbwz1uxD4/86J+GPTMSFTYujxmlUSzqrAdW
KzTQ2I0nyv/UEQ1cBEPGHbzea3a6dFfviepUgN2NqtchOGVwmhqgyryBZEg1VxnZPhxfLPioNyz7
m8iw53vmG/2FTnfn3GAwo2pIytSNZJpFK/oAmDmsHK6vRWOCKAzCHkS6W4aFnRmcaqZOaYmja6jB
N3vTimLTTq6gqElfhj1S2It4LN+nk8pky242ehirLVX+q7b3WZ/IEVqwRhmpV9zk1gxwL4cK6Efn
5jddsOmbfbVYdvy4x2xz/8jIoIA5+88VSAn/nWOcOfUR3vX0yAEwUkIRTAphbYRP7pLAM8m8EI1x
YX68tPAGpqfJfEbZfcvyy+Ux9XY6GMtOjE09LXnt0Ox5xSz49z72Q+4r8CwUAvFoZwlQgQVXoEl3
4q5hFOp5dEiPYwBUXbueEaJl1GRf+HJVeFjOom9UR7CeGCHaAzFSbHEsgDiv9CM86Hh8clDC7rsq
9fm9Nko3AuLtbhOfQEWBfx0R84VjiQITaW6sbPtd512juDazjaexONw1jpEl7tunW5VhmoJzSepb
HjMgC7A/KVEvdkRb+4vuIjLyj3ubsimiVatn/bBZmz+1Vg70ckj9GRASU6cKeEw5AX1MRdhX6e/s
nJHq0g7bsj8aBd+c8Sn0TviC2v6JfRhvoPsbG9a/SSD/aqhqFYZTwxrN6TbrjAP+5Fqpy4a0HvD+
0e3JPp75Pw9Ke1FO9coO637luRyxx4Fd5hGi/wP4CMZLjU3VFQhsuZcobRyiq4KizvMVC2P9vD0S
6Bj8TCculfmzwRGbngXTL0/ufANn8tC4RYL0sfg8J5Lxu3SCFwL6Cipp/VaJiQuds4wC9H/iJDfW
QChYkzF52VZdjiiSapclPi38PGw7P1CvC98Syn19pf5ZWeyPLKtJ/KpCF4zqvQPanjiBWRm+/Tsb
YYLg5LpBJdPSvgRZGOsDASnjVVSqz7/B6oOaZwMkFCXUl4W3k7K8MXrh1OIHKdOQAyIcadAXLDba
cNqiUIP5C7nzBZMQQ7kTcPQApiPBczJRYBAGqZbGADQk0ym8WgQCXnd1TSPp2+/qk2ew8WVH06Fx
7VNvklHi+kEFjK7lJnw3LfaGd0GDn0BN76XInDrtvUoMlEJIZ71aTHO6NDPj5y3hOChwcgWwqYSD
EkZk6l47w+oXExhQBCFhhH6JLnbpTMKADWuEEWuLA8/n6ySMfD4AlndbRQYwf2x8/a8lNZj1T6gd
YBUOz1mIuDTBKXAL7p9Rl0wg7jXsiHBZ167w//ihYL4rHbKdh70fcfVd1CJpF7OBy1cSaQgHfxFf
uT5eAUflxdnOzQny78bC3OtM5ZAvd88py1+V6p1R7Nclo+rzeEKCC6PaW5fftuF3VZx1mqN52VrV
iaHSPAHoH2jcF7ySO82eO40BJ4EMD8WcyN9205mtDK4qMJoQNGF7kjqvJ+sWG2dYpyjg198W1/Bx
yjsJwsXg/+frXdzpbikiIxzGzOibE2eIFpMEfCoaFz2WlrRqGbBAbZxx1RQf2/iq8o7S39io2hvZ
L7SeRLvGl+EUG+ow6drn+xk1HrFKB56nueGYeydqiG2HOHsh/mSxmLjU1q61XIHZF1r+fO9A186S
xsozRJgcFGtjITEo+tQdjpFYTE7/YGFJOsMCOtrPSQ0glA1+Xk+JLXiH6MgIzehSnasjK13a94tj
SftrXYFtxSHJsn2DP3E+QRcqWtkXiB6iiZaRsyYVYJAYulNfcnUOCAF+e5W+YODdY9Khljvr/yVw
OUrIM+BhVuvmaV+Q5IgIo1ZragwND4ixaPeBdbifVwIUzOs1h0XepdXgFUtRaWnPbb0Mw51P8wls
e9vn81kxyDHfk16JFLtMLLh0Mi5zUK2entZkKWtphtWXxSaY1GjbPiEjr6ChB6Z9K092BApEJ6ZQ
fZ9kxWyB0i1N6BwhJZzkCL3tcjmT6pAIgpCsbWJYMPozaS2LOcqc6vmmJQTHzeTUIoPmd/SS22Cw
SGWVar1TXA0/B5g8rBW1c7jUobEgL9AAcAlzGWuIH/Q+yibr4yUqY7QeBOM87YouF1u/9ovhvv2l
cgSmetTpwbt/E/wZozhPSIhO1enbYSfMucviJutqSTIWcjzAMe1wgYuttpovhTb/WRCAs4rQlRT+
l/hz8kp5t3n1z3KPiLyVQ/aBVY/8pwFziwMUMLIdERZEKlgPN55OUpG2M6GdCPkFOa+u2SZQSsD+
Xh3l6Xiw0rQj/rN/tQjLkQUQhSn0n5AjjAMu9jKTLs69mQq9yZi8On36B5QYs+UsnXYPvMiD3cUg
gG0IT8l/lUnhRYfv45ux+L+oh7MJOkDZ6HrfF4dqltedYmueD/RLKmYZqo0NDwdSe5hYUesiyylO
X2BHZHvNw01YX8lSiVIZ/XP/wpCOOI4ZzNdN9U+3FlJnebPm4uglz/WmocIB153XxOqlYbkJVuGn
dOUnvjc5lsqOxqmG2L+WwXwrBMTLobk6XSyaTFiGclkRsyJoTpfQXExp4DjbKdFvZqWd98OCIrs8
FYWKdwUnHbWxlmMAj9DDmeAJBzcj5eLK83/MxZAjEHCrpKdCfM+ha0oBkBpbgiCRl41ZkIeoxkPL
e9Bt84h8NCjTa594Uxive3JE40mAUGn7VtY0KhB9rPIvh6ly7W0+XaeKzdaYiKe9IPRRbD/7Mrsy
lMIAGpKsiCZcxHChdr2ajeDd9/Y3//DD+fbkw0/I9ekH2m0fMI21r2MTHyTe86HsTYb/x3tykaY2
IVw4xDQZYstQlXGL21GjOO1LaTvSgUlQ+MAfKpMhf3XrjQNmnCDVNjSggt8cBsUg9ynp/P85s7Kc
SURQbdoInR4vIk0XorKoUBrEFee1NikD20ggsmpDPI+ZyQGZKoAE2pROWNQ+EO+ZH/nFflgvqo/c
GWQel6Q1z5Jx3tFrkA2jxpX1L5QgQ/rb7zNczX7ixMN53DIaMKy3sVa+eZOVvYAtV19YyFgvd2Ih
TVQMH/CaTahHKguBOXCL3TiQshJMQqsIl3uZXe9gOi+2ZBjl0qdDlcbpqfO0V8hMYQtkN3IM3uuk
YvC9ioc29ERq1oKtEdxSByt9Cr9Md3icMeDhTu5hZteLli2a+3cxTDpjxCuVZQG6IFyhwD/kvAHy
RXdpqTpK+OdPzZ3WUulwm/t/MLvamO95f2bJlkwreAobkymz19WVt2w+iINUgaebXJEw/aFprtDC
mNaHG0k+9c7cO+ls+zZuk30EKhWR9TUSkcQN3YlT8UJL9lj1Ee46yH5MLEqcYrFGlYzOOrKey9rR
tn+SGfWoXMiDCwJc7pzwp9gA0HualrihWCONFgjp+aFOv2lLXliZeP66IL/EaNmTnB8aiqyvTekS
35xvnZCmCFcryjbrOqBdJ9cas12jJ+lpi3BsPd0sSYPAwd6+cmmqBSOA7RUy0CBl3cBHSKhrP/pB
AzhZnu8G/1KL8ylDqh1x6szoe842RlRZ5VuG2OksbEe/9C4Wz5bkg5DvW9uRmrVuCExqHdqnJtTq
ZShqkLDr7127W8rU9tObVjJfKMHo0x8OSgqrTm1a5BYGtYjIkmpO8HsBSbGAsZZnSwqnc2wH8HIs
oUHo+F41VrkX8N3vNodMTrpvYlgaUWjVKlak2HQQMXoJo2jJNxJWnP5/+x84T1wcn0gGd6ek/DXC
lmmeBNfOh8pLZRGlKtaoplWenVfQkt01f5v2E+qRLz/B6yqLPhJRHnT3pqwxEwY6Cf0PgjN31ODs
b+ztWPIxbgCF6+IL9v7xOReOPi2OQmm7mCBQGExQPS2xizY+wIEAUD65HR1SDI4BXRvmY+MgGqT6
wtYXG/OSov6FoRP9o97duzas1jPRn4UX3Ox9sCyzTVnBQWGbYx4q7BeQPjKP9yEfjgGU7ePxuhzV
OUOqPHz1F1B5aEUchHMAGkLIR9UzQNYDB3gEY8vOpwGr2WgvguW2zwI+z6CooomoJwBcnv7p2/pu
vyQtn3kbe5SD5a2IW9FWIM83sv2k5/Ctn+toITU59Ews0Ng6HrmkcGlmk7DDLogW5g2P33mCznpL
mHoRBl/RM8iGK89uMasWA06EB+cw0ndbm7PTbCPu+RxqcxDB2spvvpblAWOP/lX/JrgGCwSBC4tu
/Hhyh5yJdT2A1X/Kl5IfO7ZQrbu5JglzebfRzY1TBf2UyPV0at5MaYIBWQOa4TOZA60olLJtK6y1
iWWk0HhdFQkgp4EyXV+JU2MhQiXUYosq7WLXPuToX/ujw4CdJrlSeyLg2gj14PBiZdHc/LAOx1b8
jr0jy2uQnKyhQDuouDOxN1qI5JZTWnYXt/GeBRC9belrp9D+iWQ2havjsX9oHVj5+61GC4TX+a/6
B+2E9/rFRm3AfEAWA6HFtFG7NLKiXAXoRZUEjkJw3dIHtlXL+vo31GArniSi/qcpyQP8f+LDFMfm
5xmVwvA8ot+Vmd1xnJRooG7vFxYti0ZI3RRwqij07EEqOSFuY3+CsGcKi2WUQTt9aE583Z45BZbt
tqvnoOiQCxgsuwrdtNNuaOE6+nKr/B0x0OnCbwuJWUKoEz3DgoxJ8fxC40MkYcO0JDqVU5Rk8obG
OJHtxEoh8HopMMZn6uzvB4jjpRVwPOmAUwCv0akqJNfD8Elv1CRQPHdpaaz0EEa4+N5LrXpsEpXf
oKOlspSY/7BmW+DFa0r99pYy6onHvZHLzomxxbAc9GMNip8yXOc/cb1UVDBsIb7qmt0HwxPvWIwQ
Mcev9Qe+FNRTsHIyiVHkqLoL22S4M2KYjIRsHJoSuBPSmEhg1lkSy1MbjtSgNNdHvVsIqWlrQSrl
0MpCdSJg9YQgtDv68F4KGnRLXMOjyQd6ADyGd4rBCO8jYw4jMnznFiQVzRRPl/vkANi2ON8iQ1hx
8eE1h493dZ0SDrDaVUM4m4M7vmbHshD+8x+BQSnq8uXLb2hr307btYg0sneGaDLwpF2fTegu+4JO
JvaQLdjQlM3KXSmHSHfuHqvQzGHGLBAbUmyaIMtPVW4c1/WzTlN0NjH2WyvxWcICcOXrLEaxdbjQ
eMz+ZTEEgBQ6b+E7f5Y21Yn+KqwQnjyuDzRCpAldxX8P7H3DlEHwKTmZv2ruHZx4fwwGx+BRSgOS
AC6IAatotOoSwsg5TJ099wZ/tSYbvc6qHdG7sZobFxnw6J6MoE8+69F3Nq8IFLyJ3j0ChMg2Yy0P
ZVrt+AgVq57CMicdQ3sRdeh3O1mIdrBNXsX1HVKdRpHaCJVPidkYmxIoDayXlSVXqqLJwmwcWU30
dChC3Vmc5W4FP3Mdo1JTAW9NHY3kRiUvwqdRGHh3Fhevxp1YAO4AFbUcnUeXX7KRZ1pz89wyoGnI
z/wisZ1ZbcwsdukW0hcaEtNhmtzkHdnQLrPXkgJGfpB7hrcSP7MTeDJljHO5sWWmLKDL/mbEGhy5
g7Z2TnPuiFQdrSHkaVAuILetjc8x51lJ8gvC724Eo1BMjn/2zfLO8qO6x9fU0DDalDeB1224E3Xp
LOWBgDBqE3CidK95o5Qc9KxRqX89B6HY97VGN/2IFeCVLVghbjXwtoVnJwqw7vHH6CLPR422NfeB
DZHXeXH+t6RY8xIhkFhi8Zdd8H85f4pMKzoGG/E6ceeQ3Az8nI83JUvEdku4Jpdl7//PtCgZqTip
gd0z4IyZJxbcdWA2oUucBNbpwCfN7uLJb/z5aViN6l07mFtIxAxfLCeCYgMfiXfrrYIMvQYOV7op
EW2lIRrX1mZhj3rv6A2lIH/bkE56/jM2rub3hGToRxI7tR2kEjcbJHQZdEEqxOYxhRQHiCWH4Lg4
ZmV2avrjGj0zsE6jIcqJ4w3BBtmh0l1hMDivXDK/KtHU8Eu8bX+mabTq4N94ab75PBcVRLJvx5Kg
Rms6elma6QOUXOpdTLYr33YWOv1/cIZSPcrtVNHkZ9QuUiuR+hG+IG+vt6bYgL4GRbiAjE6FYqBT
lv77qmr6Bj/ByOf2LSQ4MSaPveG1QjPYSWQQFG62pvnPIfr0uHWuD0Pbl/sRdvGbIcQG/QvLHQBy
A+QfvEy/NoGyE5CzwyrPpl0BYF398ErRz3PMpOqFeMtTU3Y8CqjoH4v3qkCBWiGO97I4cXSpz0oi
2oLVqEaZFpog7AW/9Kxj4Xqg/uITMP0Zn9b4UgCSryX8Sq2ODNor8WqJOcN5fOnvSEXREjhi15JU
Pz70zDroBRNIAPVIVpOOuGnVrqJGQCeU29Kgab4XaJo4/rgwogdZ1TTBUdjmogiXtbDdlhjOcUFV
6p1SVFIJVrVdgwVMztTw3aEqNFYrfxC6IEg5dJH8Pw4+qA4UkCIJBYSZRHpC8J7Zwrck+wvDkAdi
Nk38Vk42Dr1FCZdxJRkYoLXjh3eHIEUEvLUlIsCn0bu9A30DFXcspecZ1W2YA3hdFAbTPjuMtc6d
ucdoYFULl5LXFv4clb45xRfuIStQZSVx6d10kT34T8NRhSwBWxKHQ5Kt60VpcE9ZDWyc2W2t90Vw
ejqKPnIv+Ns1ScQtqOxjDoBX13Ae/0d0OQDNPrs3e33he4jnYAIctxmQjszHT+SWWcVJ3KTBbMaD
hekNs8OytRPV8xLznPC17E8Y0TpAlrJSVafpeveU0q4UQBK4WnuIFGvOXsTXf0M7+UcIxkLr768d
CjqKdm1b9weBQPdTNzG5OJ0XJaFl80rxY8RqoD3XtRJmIZljcYWRwoJKG6lx4W7F0ci30fzdfN85
IFjAvj74OAucT1Mwzc84EVe+HFkASptcUJ4QMnAQwqfVWL5Ipw/cGoJZHHEHOYFzQZqtcVEvqqt9
xcmKDAwz+IEAM+mhbs/SxmrQQIJo4FOAIkYyXiLvKpyCKWeofnE7nFyD28Ja49fhmXOI67r4B0Y5
6Msit9AeOwAXbeurm9dykX/J/HFOhlSyXiykzbVo/J5E4pHgeFJ2FtmYbPRVsZYfhnc0u6j30lSj
dASOYiTGsr2nZ+JLSkZJHEvOCne9fV+7laKNqzHuBpyD5d4U9f7ukxYRzBokwVt8XjT8doxdTbvy
P2aaB68k4sfaZ4HlBr/ShlEwZ8wluSaaOiK99em6PWcCyaPW2VCEURQgusURMbKNo86Ir8NJLleb
kJt5W31GOthAemmFNRbOD2GhCS5oqoCxChn3A+MKL0gM9vxpApERYvx5ndNqi4jAl3pjs3RofJlZ
8ogQOfzt+o3pDkzhcSOZG7cbUFD/WOu8qR2WZDTrqByNtyngHrWVu/vWOT/5RRcFRp33AvtZ0W/6
Tl4K+LD8RyZlwoP6TjxIvwoX1Cd9oKm06m78PniCXq7s1TkxK9ECoShxkby2RTVMiVZ4zlksu3UE
w+5Co+c/2ZpPAX71BueBaHcpdg/0YDYSxVL5zAPBSG0+Tn3soFnS2HGSl/woJsI5XyWYmD3CTqO5
V7Z3dnSfIIr9hZwuRnGC78O6Q09g8+bOqfT0Wil4/LM1clDE+XGVY9E022ghp/geOWvXxeSuZkHc
ynU22nybx2+xfGiQsdK5D9B2Y3KDDsGXEGeoz5+QVLe5MtspW80bM2LHtHOHmrDdbBAwfXrPBh/P
LNIGgdwWChBeiTnVxc4Hc3fFa+GsA76FGHe2crYgVaP4isKSaDIqVmvMBuOSoExa5UXi0ZB7/2+e
kSZFukxJFLN7ew6SQ9V9Cvp6bUHt/U5ze9s17PfH4jWLddz+nVc0IVrmh1mkJXnMRDX2vzaGcNAj
lQCwgweEN4m2Law0sRm0QqVT8Rc0jdPU+HmjrSXCUQwkwWJzRzmhIEJqSqbBcb2x9KYdhxy+2a4J
4GAo9VbsMmzqmnAR/Rp2CGhG40EUuqa81YQo/kG54ediPMdTj21p8EGVBzyPW6BU12aC94aPimTc
I22naQKw3Ly/7BRRAyV6Xaqk73a9abZAJFLcVqYSRn3F9ZIFwzU5df9xfj2BSlhmM1HSyqyHF0Q/
R+jOE2V8RHreXGMDyS+uh2dNO095df6uqT9A2qzlJxm4awFl3bXTHo2u4q+rUUlCvfumDfvE0H95
28wVysoJCa+1Q9eICtffL4LL4XHOh6GrMdFA9R2EKUizSde8lcd6Vk1sembBOlHg2NDvyXtGHWxh
4AEgbO16hE76iyyFDQfpub+Za/ATy6B0YIR5bPN3cey0BmRsugs+G+BZhJQR6VNI/R45X3XQfcTA
o9AwSth+PynPvOQdOG2DCCDhC6PoOe/BVmJ1cF6aAVcC0CpEmz5ArnlICCWc/zv1J1aT8O5mLAV4
4Jmy5Q7w2XC5FPl2paLxXYsG01+Ayf/80BPiH8eLbO501A+R8myjAKFVtARkYxF5NpfHAJ2PX3YW
/InOn8U7qCidtYAXiSb2zqG5r+/fOzK+ZErAITniSZ7vfemJpvhEFq/qaFm9F5W0eGPhP0eXdqxf
UONO84IvTLSqZh1Z/BPD6NzJXI3tV7tzXC/tJheDYxVtsLuw4BGT3LQL8+J6SebrW8GtfP86ods3
/DvRZQEGJmfR3nrTL+yNl/cBq/EcGhTdqJOvzhmfpX2oseYmsUibQEPAvSmC/mFFWl1ugbU95MeP
yFHznEXyZ9MjI91fn1MqcBjMcMJBs2caLDbw6Szq9cDRCgrKifwJVXWsX/5z8M94QB6QiilWlXY+
5VCd2aP7CNod6qJ5BhNwNjFrOgz5HZVLue+nFTZLrlmYvY9ZvSdL7PEcY0l+84A4XLM4egOD4qIE
LPzTt/i5ONlHJXRaYlsw2/gxEMOil1ltN5BbY0Zpw/D8JekqHyLU4OxwMK7ceV0x0epSqfx1wHxC
8J8SgPylNq1Zmmwcn/AYZi4EPwpUvj5XnIO3IVyUc3OPfHQF9+qsoqtYP4h4gietLaYOWcgsnMHC
aKc9YyZTAesIJrj5XwsktebXCnovDAs976JjrWq1TegZUvOv9hdoLavn1yX7G9bNUoKx3wj8aC3S
uh0pzO1rDlXwkGvM4/+Zlx8qhiAT5vGk/yfG/9tLGnv4NoExI5b49kMwYHSIdnOp8xK0ZtCZXYFX
6NI26oLwKPYDK5L8z5TTHHTgqgeCPNBXC2oTvsYDUEWH1akNAUy/YOb5qtokMbKAhilI4ogdYUPk
WcWy8z1w6gSWo2kBf4VyjUGCYGGW88GpsUVso8MElXakTITZ7ovHl8g6oh7edZUFr3GMKRc4WX4a
39X6mkoFlViZN63gOmmWZs1G4sy7gDGf2d4FaCRSGNum0kTdLz9gFqeiTGf15Orc5cX3JmTv3Nrn
5+S8X3AjG82xa7q7mUuNbuPFFC4OaV53wSLfgCS8z+drbX1wkX9zCjSvDhYYRPD+v98Ld8ACKsGC
8iTpSuN2oOnytn8MZCbo++7Z4GPj5hzIbfcB16BfEZov25YZ2uXl94VwbUx4RJGsQg1Qz8StX91+
Qh9hKllULU/vB1MeoBbtK5l48TzpuObTVeRvsv8KGESYNZmNVNdyIX/XjpG6oskZPtS6U1zI6MSe
J4nMorAM2Ao/fI1B3rfTn7mP6GlqIg22UIfpM2h5gBNRaaJV4k3a+/8aZpTo4cBdiXtYwIc+klMJ
I83mMHHUEDtAlrNqp9clrxo6Aik4QYef8/prS0BwRhZdUuR2glY0eZYl2dA9PqzCtSU7DTVk4fuk
+N8hAqlq2LtsQutv5eS2pJgE6JDQLJRwLs84IOE5OBGlgfcoIjFvGBRlpT26GnZsm5wMZIfYHlZA
q8j0LqI4lZPb8wrA18lKm6krTlV7DyjD8t3Eok4sctxxeBAVTTTWb2zcfcIqS+5kP/ip48CteIjg
ghoHhY66NypYH8R27ULJ1YZSzU+TT3RZPqI9LKVP9Fvr0Ykn5I5bWakvSU3/X3M8tCGPqQYn0BTd
Kxxs7exyu28wtGLazCvu8Um3w4wUHr6mjptXyc7MyMxqT251V5nvyVadA1cIjZPYdZqqYSFG14ae
IztE5Iww8ul2yrf8o1cAUm/L7hc0KWea0N2K6i+MKj0JcQoVGL6K2yP9lTFZ2xTDtpx8+CVh3FuB
nyVxrvTtbF84MPCmayOmem3L2J1AlKuMdSAxgsrG2FNA1R0Gaa9tYKN4Ay+s3bQ9h3vrFHT+Hss9
1KeXRxaeyFqa1yxx2CqctGlxzW6gL8BS0CThHZcYR8oJuKiS73SKuEFrUQti1At+iQeWXAldQdWX
YURTBE9aZMe4fRSbED/DfleTEmXti8+yuELJAjdVh+sdiXP2/TL1tLbDiUponJs33JVpX3MqKy5D
GN3MNb2HH4pSioTwabmTyH5OPIYBVB/V9dw1MQJbgJZiZGnAMUe3q7Uk8dQ0JU/e3x4hAFfJbbfp
hnhMo4DNXMwwL8ZK/XyismD7DZwvIRjjY1Y00Tg1PwdU+2uD229x8DVVqwgIj2C70LN03TIlz3IM
yqTAdvvsuBG2RZ0AY/bfll8t4Ft/7Jts8zUZ8eQAO5o7fImR82dR5Blq/RIb7PMpoQr+rkokOwDN
ax5Dsn8msL/dPi7xPp1t7G27Y4zwdm1l8Uq0G4G+pqTiYqeKMzApeDyBcIZ1c1EXgHuZJq/tNMnT
QEqXVCakgHBVhzLpgkSHNCBc2hXUvoy/jx+ZEUflfOfkM07P57IQCMFJPEPu1fEyYcRB20sND4Wq
L/FFFW6jOSrBzg5uAakcvNe+I2mm6CGhOLFu/2R5ngNusllpHtccDJ72GzObwdFG95alV7SRGOaL
dBOOyOaJdZY2VlxSHiASQWP+o1goH3O31g6nkfz94XiZbTen636oCuO7JG6exxvk6TWCEiDiWlEz
kmuJYOz4gyM4T34tmVA3kQ3Hr6Ywr+DBnk21PPl99wjuStC+He7tIgn8zz3kiGty6N9G4ps+UFOB
5MxO9Jp2fnoLMZRPT5NAXj6NLYM2fbAmF2v+BkqXEkvKb5gYHmvDMn86hC8jsiykIjAMBW7DW5Xn
9zZMjRpOK6JbHWNi2c67/memxvHWCc6xEWYaeqUBvHCsB2Qw9THpIaIUIrTzdkB/Mw8//xE0JFN2
gykjSfwgUaDmhNIujw5vpwwKN/HRwIRqn4bXMqlG2M/a6Npeds8w6S+rH8NvCyDZIVMu+473ZfLR
FqiNkzBH198buekvCCrTro5Oh6T14MBtn0uErtAv7PSZVuA00s4OrTRU4VnKZ8UaGy5a70yweK3I
PG10atl7igU86wg82nnNYHjeYwxKibF8JvHYUNM0AD55Rxh/0rmt1uRd85kKk/AJLClRCaw7gtuU
GN3STQDOsoJL23WHdtU1Its/PB2SC71mOig6yaFq9JlWvR5WvK+Y5cMg+CrhMassdixwIwMjWHzU
RP3l+9DRe0ofGMQGOryUfj3gWcnVotKoco5pIQxUu88bTkc3kwiOmQjNKNyQvWeHR6FHwDO8/Qa/
DqwH/tToif3JLHlGJEiocRL2xV4b+RSauB7pnNjNfh7I/cGs7Egu3Snv2IeXWNBIVJ53Q++HzOhd
aRiwYyQgCun5yfZ7JAfHTJpI0O5QG4E0hfd/eZ4nDRg/tJEL8uqym75zLb+aXJgf5fPQyNiB0e8a
8bBDo7iaiR7fk8qfCS+6OzamcRqtrmoCUJoFkSo6+y7g2DPHKfwZIhM8lpaUBAc1AeJDRM4aIHAB
CYorHvaqe5tXHMvYgL3MT8Mvx9vZ53HtJtRyVN/aFaSkn5IV9TErFCCzJ2TR9xYkIaBOHnZf/mVZ
APsxi7iCHvgD5Ins757rP5S36Nhq/KTjhD8tzq7C1o93YMzimLdMXRZhZSIpiFS5KHc8Q7KdXyLm
bo4fklImw6PmFSc1k0kUcocTFyZxOuzeszMILH8h7OMh1/D4rZ7NlYs9xstv7D07B3lz/MEKG+dm
hyaIsPXwUvEw5HTc+i5kUyporad8KaeaW3ALrkx7L8jEDEkaKFe9rawn3hx8XPrhSeaRl7NexoF3
pOVlPn5LnZKJ7FkpUwT51me70fCwXwz4BmFiB0YnX+6LZVpds1m2gvZnZv/uLhp94BSx2EmKt51R
F9BRMXk1SMZbmp85f7YKW5AFY99ntmt/UXV+tkfpmM1+rB1mltOBiBFjEMJJGYsEA8X7X4RTRbsv
ocuAl/ARKWemM+NgNkK38kV18JoN3JW5WzUwIiop1ImjVYcUiVK9H8agYkhv8Y+m0RqS5c2DU9q7
3Zrl+d1vwDpG8ddH6TqcStOmMwjDUXTRt6f8IeS88cgYPY+A1ftOx2fSTu37/zoshBE2Y6dqtaBH
hsHRd5ldsYfAzPvvB0MO8IzdREUj2xtVHBwU6G+GBjiNF3oj3gXNS+SYzrn6/Ogu3pL+CuPCNzot
ppAW66kI9HWOQrRmC2uHu94+bQuqH9voud9PcyaXHvgn+7y2RFf+sev+Tx8BzWPQKvOCbScTdQ15
rH/hs1/8SQYvfWgGsAaukbqXYNzqPprkd/VYuDaOnZVn2eE56/cD/JaCMd8kOHVHb2hq2kQDjVfr
hqpGX7plwj6ZpE4JbBKCbb//knUyS5ZiJZWoSnNiJe57203leYzaHyc2VtSRX1waPAyEdCUnN8Xs
hz1/NsIIAaGjnDB3JR1t5OSAHcPxH5GMcf4YiuVoEDSVkYY5qYo7+ttoKQfObsZN4n1+sfh3t9ux
YODHVn0nt6+hutM1fCtB2GRt++Yf3VY/7an4NZI+l2gS1swqFxAGRRJgu0Th2MJOq3lRmmbcWJLR
vue+pRcrMFRwS2V9z4hJRbOkfUBvQ8JwWxMteAKGfEk95f9CAhV075/yw8cerJJ/28rL+7z+9fN5
zcoVHg0R/Lm+OO9IwAfBWfGgJ7fJ1LCMA+via/shFYCHjcPddUsk2mDO50hCpNIi7rdKPYRHBkYD
Ip/+zZqpcfN5j5hw+/v7K/S2ehSKiDfKyBEYg7u4H9xVQRDON26lS+6uEmrswSL5kB6r1mY35fD8
L19HxDEU++k5+Wwv/ju/lg7ZFHlO/y9cN4l2oaN7PEwvgbcufArAxdM+qPLIzM1O0QWE9d9kjaTU
Qeq/O+fOvA55vHgXJt/Ol9o6CrdwHaOStC5j7nYDxN0oOCkJSKTJ0jub5OqEdgx5tYerk5slsBVA
hMYvXtM7x0DSrqLoWp5HQ8fgZx4kY8P81Iu3rIfPlYLUC+dw7/byRr6exv/CbEpsN6B9cO3MzqVd
3BlFbn6tFVlCk4LG56cz5U4+vVRFsrSyvFUA0NuYBLEyOP3ZujW3JemCaAG7m9UMDibSoeiuAFaC
Y0mWskZkZy/7MQp2laStCLaut1SnCjJUHSLGle98ohlV+3ytV0bt/6wOIVfbz3iyUFhGYsnRgBuP
u8mAFufQ3d+2o/rNdSL/MkK8WsOR+rKvl9OH+d1nf9DzKCpgFIlkvMg59a1Kk4EtskEg5cU0arR3
REvoxaB0axG5Idg/HOJfvo0d0yUkck0piehMuggdKF2fo7kPw8O6X/PSXkGZx1pi5lurjbP56H/H
nImMurApe6knqPW6qPYKa8RumagpWK+b52/YmAQ7ocnQAEMT7Pr+pbLTOHlzp+iVWt91Y08M+70s
W7CLcqXCVrPOE3QPHEZ4gV8XJGYd3kQ0KGUg8EPKVq6Y+eRJdQI5549gOKuldjN3hT/jAl7hx2Mb
nEUYvrIwIB5rXm6PoYaeEFxOmvOJ14s5KnJsRurtxSyaddANA/UoF/0A4rkoy5nPm54vGxNoFSOh
VEbA/wf8BJ9eRyunojl0HqNNKuxN7adb3L+4QRePTomuj2ky3YAgNGJvmAX4kUU+4AMXaLkbYMKT
GvU5VnplFHhgvaQOQhNYgMy/oCPwAuWpx3jPXjZeFQgonOY6nT/rss14fQuzAJmlpmSEJOD5z2e4
WgJLIbcFdYKXlVTDvUQ1YY3pLfpb9/GiJ9sIphtDTlk6i1iOk3ScWuodZqAT97MMXq4kUHk3c+xO
FVeS77p5lBOhDYkIsSTHIBl5BjzG0mm4td3f2b3oaG9br42VarZrp4THYCvuxn0BHofXpulRK2gi
OTeHRMe4qkKXcHiMMWetF4W6iU37w0YEGf8ndDJDEraojXnktyMVpDngEoZEEKbeTT5RbSNIhw17
3Jdgcgf3bnun7o+GPPkyaBTxoNzgaXflDbSZOF5SOAb1PJ79EwiSrLGNZopClhNH3aG3v7uC1P77
u62HZ4zIqzMVgastnzaqrVA0IIKkOg+NrID3LPqwsBi6ICM74TVloE4CyFWh+lxQJjpn7hnplzAs
UCFQBCI4EV9rzIhKUPDvpw3cnlmcAyYnouOkzGJcBbfBz7GbQGSj5xoxGo/TUeVDR15gwl6G/MvN
jpdbrqjWHlfD48hULfFCJqEI+tKew3FDUx0E2njCoNn2scrKtbgCNZoVWqjEXt2qfpKHKdlYXKxB
tuSdjhJhTqgo+7sLZi0TMAKLD8+RzhvOoIghy3qw/h5foHWE1g1x5IEjRvW+CYJXcuGoreL2VcHc
OJQwdV7INdQktBT+ZjDQZS6PGcprvZxuko6t7pjK6isiuYlo6XGRfoAI5cujzFxezclVWMhspBEd
FdBHY/bO6BqEv4ZaZ7SpSZnFB0Q/QyJ2+8tPPGaM0mWx+UCG2WmAMXcCU3FeNMGaguj/WtzZjCA8
1ZD0nHH5Z2Zd5dyjL7z3OoLhfNl4gcB6wIg1KSIyky0v5ijg/gz/+9OifXifxSW0MM/KyP6oFP8m
TO9ayYl16x4FyE+HZpetmyCF8HMWsstSN1KcI5cYEN1RLk+RAXYK2iavqi+7WtTQgW1AnmeftkBv
kzTYJZ8aMHt6sbwdocWy7SCL0dQMXgoIdpjc04g31rdNT13BfwEn4LrrEUWWb7vBv4UjlRpdGGJO
T0R9kXS9VI9C5sF9PaNfJTRn0+fpg1iijxMHpiPq0aQvA+Br6HA3X81qAwFJoMDODBdWcxhwbY5K
60ztLpe/DYn4xSPF+PI+JL1nTFQzG85ReGZQY/AqcsKyfFjGFRz4mYXN47CcW9NZwevkp9NJBjwR
Vsz/U8UjQQOkPs0qlos9eB9TfP0rB3QDZrJcSDP2PPiHr1Wh+x+zidaE/VXFpRu+Wm7Q61K2v/X5
l68bP49JAz1y0rMlBJQHPGFIov89MYvBJegymIfKGrdabn8X2JwCFOrK+xeIFaXaLFCrfHyS7kZn
zRSf71T0um++wou63YS6oUofF54BeIzFYWqeStqozv1/d1zLU8Ke/v+o0Pw+VnK6ui25EPTa0DiM
ezt8syTX5iBAsvLO0aORKPGUHQwMGnzYj1Vm6dxgHk5NB1BcPBmzTK75D3HcYLMGEyEVwAYE+OOq
rKeterNyM/q2UuLWMnDdMHxjlBEtLubC9irzCY38L89AW8f+FGrtzyLLk9PCCuoAjAgKwPjVIUuy
h5YZWIXnJRcMi3MX1I5Pnr1Nl0XCQJCe7sqW1Q94fJpmyoMmDMppHvOrx79DsL9oDhVZZ8f/E88N
CB1EPPQuAS6E2feJOkTnT6R2JDMbYTum9Z7+lIEhtDeBTENyX+Vf648n5/9iJiSiHcE2AMP4wAH/
r01YxYR7dIGPgttPGCVj07P9PHYOe6s2y0gmxKBKktPnOTeeeVmc9+Hf71/7qwDtVYrA+lZXE7iQ
rIWdF5YGw9xhoDn748ArIQMDP2a9GJmOuDjgCbSNITGP6UvZNf25mkrJEjvI7bChlVpPl/itD0kw
NlfvBxP4k1J75bSEZ7BklufvfknhcqL2v9LoBYVZQu9frfHmUKv1XWIdsa1UbSnC7Lupu0x5SNLR
IHDZW6jvVUjrJrlR9mNgdlXLsnUhjpd0fTr5/Y+E/JGhzzyGj/5r/odWYtyd7ty9peP9sTcBY85s
5nC2nuCBw0vxkCmD20cVoq6IRurombhrKlOZcl8Ib9ShViK3swiT72vrlnWQoDj1ZZFNB3SOYWDT
lVDgv6FdATFqaxtRohQI0IFKmpNogiTUcj/dw9uqLSHdm7Vz1TDvJt9j3MjL1K460Y8wmrc4YD4v
PouU73W9oNujcrfaYUpX2TtfhjpeEBm8iK+99C54I72cfYRpLKB0XvsO3azqxB1p3Gu3LJqib7Gm
QGfZ5g9z552V9HHXHcV02lNgQlxKNqWmVp2CaSfDDDBcAboZaN7fLV41UaZDT7pyopGrikoeIbI1
rvsDZk8krE7tDKuNgs3El+7tDgD/8U/IgLzhAe9qYCKran3xrdh8zvcqONe7IyEYxmRuD0JLcTAW
LIkVu9oWj1BFO7+FUIFLHdUku6YuNkqmUFeYwnEUReQ9GNN9OFvwPzHfsUHdYbFM75UEI0G1OsqD
AXwT2WVzPrqX0Ih763autewTYCCpym1J5m/xVJWqOdqUBEU0QfIW9XZjX/S2c0DfeokKaq+LVPOg
OUW6E1ydCqUfxKzpRLcV43GjjbmBnx+ZgL3tdrW0r4OCiY6SKdbk/iKzPWoqx97KhzhKS4LNCyIJ
g+00QpKg3U5aq8ezfPCV5CJO5cNGNrBRfH7WtCubZZIn2sxvIqNHbdpeJefd9l8RIXA+Q1AeSzRu
/Vd5Qsj9n2vCWkQ0IIQ1sN+EiYjCK03avGXiYSw9lrCFdRqPSpZyM9jE3CtuRUTEXx060YYbuYWq
JtXGpp1iVwuAhbf+NRhWmQmP7blgTsLQtO73YGDGAVBn1BFCiRbUzWI2K+fcvnBdBpgohpOuvJXU
6+XnZz6kiasDNw127+9SqH13ZfbinMJ/gzLBLIdkL916NX/dJqFabBEvUKxhM8NG7+UgeP5iH0cy
UJEFQH9AfFJXLSrK6Oor9y5DY7QwLG0/vpjh8NJIqqmvLBbdgbJmUsJ/SXX5pm5KjCR8ydi5JUUW
wyrnmVEfF4tSNidMeZ23HXQZBDHmgu1Ec3PDQPDXne739WwsPSg6UengRhpKsKtB5g6/hhbVpHx3
NR+zrHkTzbo5oL0drEcAO2ZtCQ0YwSPIx5UvZYTRvoj2JA26sd3i/EUvdt4F7aCBTSy1fYmGJJRK
h+zqGZP9r6cdIAabYmyf7jnBjn3RwsuOLfCcBnH5RcG3tFpIL+aKKtzmObxm6tox3G3KnnbkpB3F
/o8e0cDiWQKb6U3VvrRXhqVDCyOnxeaty3i5MGDxuraJDzcCDXQAoJOMZRFsl79yG/yj4JUGRxqw
5/qFRAJOonML8zIM7Qn6gdfSN/yK14nciktFW2j2azP1q5MuduAQaMQt8IVUqgmmIJyuql6E2HOS
0mXigk2rgMuEZ75+1ebwsqmwRAPcNCjMa9WvkJIr4RGrJ+zUMgrihIVJuRYXzN8PB0wAMZ69Hl8d
su/yag6I3mwzSYzF+D4R71TlgZoQmn/09giERLn8Z1cGuakmhtoAREh43rZvyEXcBZL/J0y0tmv1
wM99xLvZ+06fPU8REPwc+o2Y7ElTuV9Iin6E4UWG1pZP3mPu5Gg4DgqCmikW7wJ3imE45O4XEd9k
p+WSTDu8tzi1OZMfaBlyY3fpJkX08nZ0Hwmb8udvZzHKTQwWU7UXtcVJ2oxtZAoAWY65vWRf6SZn
l/mb0ymeSicr7uFWCJG2XNFYv6dVCS9ixrKp45FUE9A1DAUXeXAB45H/WvoSB92zgXFqd/AdOfys
+42dmbz896nz3MDNsIkhCDvF+/h0LDo5RwvrFnHu656RqAP2xiNruGhjxuz5uEJVaJK27UkBd+VG
akMfAtUpQEo3VtDutVTAd1yYsB17d+BNGYIomj2hR4N2PBd3bckHIWThKcZoTRETg592x7ncN4Sw
DDhxjJ7Ubb2RS+vUsZ3yROt0PLUjHgwem8VBQcBfpf6ROAiqeek6Krl8ZgiGvJzb56Y9W2hu6ulj
/zB/XlIx7iBLn/ZVIW33fZ8fvr41EuIZYe4RvvxJ6s4+2CdFNY2yA0j5KqBPJ88cokJeQr4dzbfP
CUOcO74LS1HvY9D024c38vcQUlV74IIYACdNSaqavFXsoXYN72gzHjVetbUHKTNlUtYeydlrwAfJ
yqDMi4OQcVr9Danygy5eZJ26+anpA6aZgjSud8OfewDn0cuxrTeJHtTclUlgwdQPETvK06k6PZMl
fQQZJKvL15sEbeUpSkdfWHYMUNHwvme4GHqim4EH5UlVLkU29WHG4EMqjYKG4r1EodKhBDjO7FL4
UjnT9hhlXfoApGAnvoKYi6BnxSFEMKqjuAucWZgV/kpndFjptgXFGccSpDuOMTpm+2pZNat44Xuc
NaCSAfE1XcsqAaH0dHZ2NPW528GQVTjrDHFWpS1izPL4NgCXNP9YOGGLXS4Xpv1IEPTR29desz1h
JqJtQ/xBeWfaZFIM/6niGZS6U2L5aNMyvUHfd14FUKFQO6p5Av9S63XOCLBUABCdHfleADqZZ+GL
PlQThdf0W1jyuXtUv8F3fexx6B+hMehncFgBISCz8Uu9zqPl8rDcPIk1mQ/1LUO/8YR0oymCPC/8
Y+6gpQIpAFu0MBzc5pIENaSUk9QIfu5vaF8aaHziSb0H6aU2HAexkIfG84WpTJKE9xs92rFkudVW
USQvPFn2uqpUg6rUejlGDZCEE1VZhJYJZJuMoO6MiJxEh4fBtMPHI4YYtKITfxs8dzz9ODOUWOrX
LhYPshN7vzqSc8OTySk5bneSPOyQBWXDkh1aZnCA44tm958uqF68zAB+K2twhvseyawA2IR79MUJ
tLEGNtJvkPWTaNqAaX4jAHZp6nxrOQ0wN/bGNqyYMgTv6DF6TvNEwbsNGtObhqVwMcG2gq1Ijk2K
rlXzERVslfEUea3lUNC8XRqaGMD5mIUPe4FIAm7RKRT3M2V1O6GYAVlBrl+GcCB0mHWBXa8NPip5
UZopLp5UNttQwUJ8KoP2/ekkMqfG1QL0M9uhphgheikecoa5d3bGFfoKbe0eiea+Yyut2EvUECl+
tF1HpG7TiPBa9DS9pXy4/v7twlMNdmwv9aEeza4Px1TMdo6VWxvVs/KKjqXE5zImLXkRDcY4Gva/
Sq3zNRkpxKfHqctvHL8bpL25SOwkPCRyZCrEmei++FCTkRe4UEKdzjLkmETCw/6hcSiRJ3IqIt2U
kIh8P9aJQHbVK5Ao19OvtO3itJ/DgF3NWlht1/hqNHDfuqXaptJKBFMe4bmzFDfgbpl3Jhed7tCi
FkkpvQI43UNVaOXaKrfCohi6OESTmpbxhxXG7s67g7miY9wIriglp4ihVNj5A0VomP9o9Kb4Bh5X
+QU6vyA21PKfdx93ELvZkQPsXv/19iTsGPfCb7YqjER5W0Tf7ocGUcdBHtoWi98yF3KP8bl24Jg9
J9unA/+uPoufYXg92iQatEuM8saZ+PMDyovhlN6zuVxnAt5rNWOLrPXfJN+SsJJKVI1mT5bFxEBn
6ro/MsvO2GEK5hvbzjRSR0mqKc9bmJg+mw8EXjXOqNET1xy8khQ8Wqa5RcJNAKGmGagO
`protect end_protected
