`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mL6ya7LNT0XPJgdwP+Qhpyi9/xfwyNN7pNwgnBNaVc4iqvL4S02E50vZCkVVk9Du1j0loiSALVCl
FMTq8P9gYg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jvvSK1uVFrRsmh2QOXrUBxukiBpcpWi/eNtvRqJFK24YFGCJQ3+n3OOvorVM7WaB3fjBFMhVRg/+
exuFDoPw1e7fMH/7zsMbUmSSskhz/NwOhrIc64W9bnjCjBPOh0hCSwNFM3x/Yw8bxxedLyFVQFW7
EMh9MDUj0t7f02b6e7E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A5YrMJlDfxUAFuiCBj1nIdlI2XBzbZ5W9eBFy/7HPZRvCYP3jZ06PU8A/+ab+AE7+plaeM+l77ch
aZA7O6cQqpGZUWv1LHca5Whha7qvN1FBsPsDhnxVChBX5wRB8TioJis6bec5Yd0eMrYJ/eSZyBDa
jY5/RoAQI9sgPJu+GKiUtFRcqmFmw62m46AX59+lyVn//mXeQfw2EXRsyBUPsINEOq/JGnctzTNR
AZS+A8htRJNQEueygBmctBkWBuXSN9o8RoLiISUrTBEaUBhb7ZuVGoJmlKqcxoG90jZI8/T/zZS1
d9EdyaqxE1iCR9LEW9wr+iZ6wneijYN1L4sgBQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mja+I/qiuZA4ySi+3GfJaT25/Guq0XsXnTl+VNZxFsFNXBcvGpWLVhF9BkOGs4rsEcjOu4IXKl/A
6i1MpZS7hak3VcsWOpN1tX6Q0qWr/k7jPK9NRZWeZ4WvZ2y3UddFKA11NQJBZxutgLt/S5ZVcclx
qLNyL/L59OX8MLNIPHM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jx9VSHMDOhn1BEN7mZjuhg4v4ONyxUuk+BnjOOqgMXpVm+REwwF4x7fn2up/zkQrxYupekPKyJWj
/wLN4nkg8dNY3dNDTbQF/2UtR0gShRYAcq+bDyL92NIogE87f3c9HYc7YQVzEKr4TlIZgfg7EDoT
wpTBXIZb6Rb6nFpFCrTWbJbtVnNSiuitwry4kcXTia7zdfy82VclgqIXmMPvw2SqejRINQhZLNWN
3KF3V543DGXzxqrz+FjOAxzPAUhvj+kf2srT7tjJodAG2b+vJ+NIKt26cH+GcK/EWJbwLWFPA9s9
9owlY4KFaZpck6n5nRpOM/YS2GpTGWWywQ7adw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5280)
`protect data_block
zhrNWXoj/FhnPpvERHx8FyYSQwYFEavId5aSGxplSK4mTwLDGeSAYUqx+O1cHf6UOIODeD+KVD9O
luqTTtHYmyG3rGmexcUYaZqLw+vc2pWczpUodstTIuWHcYIzlT8ZbdYjD8B2Q1OafmrmisyBga0Q
7PO3D5pSrH+UfotfphVdcz+wDYDsfZt6uzLN1nyRhU091KbT+KsWcej3YvumTr2VyAxwo75myMzJ
ms4LwXEPig55Ywuy2PXE+D5CjvVnJcvJB2YFU5ZVgLNqTaUykMs3XcpCkGw3MKgpEZ3ro7UYtYz0
zBofy63jAKZLPL1dxmCOHDB7vzMj2bBp8WHH9tk7aoqDwHd8rxDEA3Uqy/DKelMF2R5VVfD/3zbH
dLnVMeiNl6eQgrqeWVLyUvqYva6Cb3ZT4JBvUItpSBeLuNINwXdf4LIknSpeD2dNVfHHL+v91Kny
3gaWLLPiZLUou8XZo3Ob6d6yAnxgehASOSjIxodAfE6lmDD7JE2VL+aKEdHXkik7uOmTXVakIJCo
OIN0wPhDSOFA0yoqPDbvYAM4qwnNrp6DdpomwBzDZYHO7eHsRLVRPbkheVKRclg59O3/vnL5aHZY
1170T5Jy5/+N4PJmuNXZTyggG2rodEV0asHFV8KdvJyYIHY4oQxr+JiZ/OaQyshp1KBcBd2ZiB/N
qIPIH65+tBuupk0eLkl/T5RFmGGHH0pYwyPSCzrsdvBGVI213wARGa5hWoUTcQQ0lAM7M1z513RY
B4y1lOmOwILc2otzFaxlvi12YtTkr77X+kXS0G2KSmjT/UyRi7RRyuhDuXR66Qk4kESpqElHjL0U
oZFiu84vdp91LkVXcKSu2Pgwmx5d4y+CUqZ0O7TqJE/E4kna52CSvQdiKGCuIF7HusB/ckvDuRQ/
hzgypa+vplLfKLYVY4ymx29l2Cv+dwmsgpKI17ugGaA/SpPCo45wVQ1F5IuOyiFih3mUgy7CDke0
bo9Rk1+9EFoyUlcKGPw0bFV8WYkjQmxPTgBAYHQp64bnQRR7e8dRb7W9gyXmxM5mAqS7MnYLZiAy
P+HVeiQVjk9O9dYHysx3iLKw2GMggoOfEPD9UJCJcAR66gK/GOP8lxrRBXrj4qI5iJpTcOg7TYhC
b254s2ESHGMQjlcjEcv9e9Y5djjVd5Y+s7Xtp8tl+ln68b0QZz278qt6n24sAcqnnXyPTdF5LDvh
Owtv0XkOU4AhergIi4HWdIHNIU2DpXx3uU1tbLcFqwiskpr/vHG2heNBaDtQDcyfCzVFpqupT0Kh
5j6aJNSP1Ay4OehwNWBd2SK45RFmCGNQkNgMHF3nQUIcitz13Ct+WB++AWHfyKC8n3CS+omR3tiI
hBwCHojbfK6T15VGYW/oLipvvQsu1zC6mtMo6f/7KSOETz/oAv3oqkAkNaXitPr8wfNXcKFUd8pf
fOxu80hWSONOkHLi2badRePoGqeb4YsB58PTnpNH4l+VUuk+76itkmxUrx12SY9UiIg2aHVp6Prn
ffmu/XEclTypMXHjobNvaVG69ZbH9lBLd7KdbabHaawbVPaD2gVmOyroFEzgMQQtr9d/y8c2eu7T
t8IGFs25pAABBswodnFdG9eW2Ik745vEpH9ZenKmUe0JMCDoWcABEUQP/ls40OQcg7wnPVgb9u2b
iqqFXYh6wvfD9u3UVKr7bo0P0uQYuF2AV++H6Ubsj0l+4sdPSu4MmBXtD9kyhiLehNqSFTIpg0Vs
frL+3gMHKfZg/TzynxOrlJ7J6RIcqevNZggoaD68H40PNlJVxZoRBkO0RTW37D9RVlzCb3/u6Dni
7Ic4aDgI2297Ne4mqtTPSEYTSaAIHTo61X/2xhKDsRGfOX2NJc3s1Dmg17SXgGZaaxsfSpwYxDOL
EF0/5UbEF4Yifv2f9ngN3gv+XDZOGUe0eZW/QJXGlTX0NZakMBPR09ZrOTVPE/ULQwzsOzDddHCp
tuUzMN344oO0hZUnr3J93LfFJujfQEWScxstOCdU9eWRt3EgL2W/zzhMcopwR+NiK+ZlKQeMzPej
HWPdL9LyzOm6KrkqQolnvXEXqFhAv/9K2qWSIf0s26AS61BpDOMYJ337m+9LNlxlwDQ8hUaCh/MZ
Arhts3ggYbsm+0hYz9yAojWko7YzRf6/M9GRvsvoJU6mSbVatsEA+YtKry1z0GeGQEWyBLV70cRK
FlSWV2T80wbP93Q+zNuxlzS2exzjhMTPE2wAhWNBpSqU/RxDD7gVjPArvthMR9cihNcJZ3EhIJse
FqIea/6DZQlnatCAWXz157nKOwPppYPqJbxneR6m5zM4XtonmxnGRFWjnVKzlHbtzwrvKT1jH8KO
HPEj+id6o/Y5DoKE5t1kzQHsdy7M3WtJObF1/kwbLepNcnr2i4cxFOlENhHPB+ZCc24K6AmhG8ct
7Mb6cIo6SkDLD9v2EUi75H6wfMLzbvCWbVAG/aLTTxYV+7DVK57gKk4H84+6b6xfnFcEfzCafADD
Y7rvOTdxZeo7y1Wsuxaa9027egujtI2fS9PrFBFIdysO9UgCfz+bAy+TRPAOCYl90WKLYY0x4keg
3ty4I7SBpumel83S5rZk81SrU9MHCoKeMK5EFBT3uIBZWp90qdaquhXFWWjoS7nksZjsTjESTWpq
jicbx/ED5U60buGMDmE4F369OWSRGgjMKMvT0a+oIT+NWyYUOXcGJf4Sln/ctwU2MyX40MsXh3vl
Pa2TKVGwbgHj1VJirPgHhJZIXDYoGp69Yjq4PhW2l3FKDUO1FzqTqydXJ+2f4PqsGSdcnjecU1wr
vYBdCs4FCVRqe2MwtlNVk+XoqqMzXYeJDt/+IahhhLvkjnOM0/tbKy4aGgHOpCUEH6YRQIrKz0QD
lip2FD+p0orfLlyKLKDHV5gj9rJVjxSgDZ9EjNqSXHyItVv062Q20K5blKuPUsNHEZVsI9Sskobf
Ya4VizuG2kimpRjRNdAd9ODHJXBBkXBEUvBcggA1RaBLweXCdRLj00wvUQbvzne62Ja8Cajuzllw
M4N83hOBwPvx2BJbWBORxsnOEP0lEQ9ja/Z7WoMSJAJ0uMncy1bYsIhKBwt+zFB3POxQfPILCcm8
aLSLbet2v0yP82pSceCZpSXiKgvG7KTthLen0Pj3y7Rwt7pBdytWkZKNt0HOnEDzkv34CoWD+vrJ
KYc4OLLk26uSG6Y3KJ7tCPE3XLPIM7txLk7TkX6wgKy7+P9dE5wwySiugU/idzt26aCcPna95KAD
iLkUs45B+ZG15bA9osCFoCg5zr1jxdeES2hguD+yW1Q6Cw1qvTb93zJl03saX0qe+NQJM+IPXXpo
nztsbyi9enTcwfbAMy/vg1+KcAxMwsLjJW3BRS372gS2xuP6yu0Afcx8ywl3zGW0//YQOJXIa7Uk
1BnCfuOY3U77j+n05FusPmwMBxadDIeKTfZGDzVpJcAb8rnivdXHh4Mda0IMipaU+ZtcDVGEuF48
v/PhwI/RaY7mP7EpCc6FCwj6QVIUq+7gCo1Lc2yDSvWj2rX1cSMpBy1ncKSnh6VDmU9y8mOd7osl
95oDNbGj2bSQlPBGQGrXI8Ndyq4MJ3lX8aH+7PksG5XesFg/suPAbg3g1DUUTJcrkkQ+k+pnR6ig
sye1u4bE1ibzOGRloEtl1IuVfMTdje4ThT4GwwC2eZu0hmPhAfO5ToF4FarQCL1gkjv6vlwhM0Dg
ra5gOL+bQKUwNRJFvtdJ7nncCk7p1gyDuirqnWtLYCW7dfzWplsuEkhlslR9LVjg8S5SzIaxLbW8
zJy/Dq6/rRCVAikEvYUoGfRkQYiZ3O47CAhJTWDZrBR3vNQkMTq3z6KjNOSTsI6UW5IhBBGOmSli
Byi3fdOIZijThyoEyd15v0fM7ahjsQTNsT9m0iYOHES0YyGkpe8qjhyaGFZwLoZH0LQyl93J8AJW
k44u287el7w+LQmdQeeObIBWB+OWTSnb1T5OuqL4aBBumNHj7VS2SZwUECepf1+GC2WwLjNJ4ILa
qG6IgvczRONO87E0UUNC+8G0CVY1OPQ8EqA5hHdTk7lWpHCWlXSBitz7gCypvvHQjFDzLLx7i9WK
oKshfkf1s7moab3uyK17DLjjAm8PN49LZgWl6RJ6ReO5cukdHKzmJsDEh4oiio3+YvIKNwFo+zcw
MVx6FCo8MgLofG5geQLPSFIksv3m1RX7zvGbkycQxGhvDFe1fFNMiotNfcEjffB3YikofeAJ+MN6
YL6fw283vQEJ6n7DZiHNoKEUqgR//PZBq2r6D4QNigLO56cRuoNfxAVmB37OzSZlOUBPijHhuj9H
XQOO4Sgg852Cm5lKVZdGWbIqo+39s2WyGlrWhe99TjeSTqfZCNZ5TQQ+SLRfLLVh1NYEAIIoNmf/
Xp6z/q2tiDGvvYNKij25XbM+UCT/GJTljAj1J/4H2L7x4zvNJ/rz7ZsPQY1yNSihl0MFtciAGtTF
ufkDopVwEFOFxCHr0uSHk5uRe9ojhJdKfh5lZZjfUVr2cno81UgkcEEI36SHbNWF4ZzqEJQ9P0P0
DbaZM8vAoBu4aV9JtiGrz2OZSVg9FEBpolDGH6ULrOyb1qqSSHLnauRG2njx+DqkPyCh0zc4Ebby
rwXNEmVfqIhfUxg9NwnA9qafVnxoeN9klAQxC1u6R88HSrKxFNKtTzX23T1VnNI6eKEpRHJlsIK2
jhGvaVEDUHnlg0ihEZwZReTHTP+WPPVduNnROz8WdxAaIgnTfYwMPQUm9lgu2sA3Bv6OhG1bMpn1
rvW0kmrqu9TjU/UGIMczlBE4XpikKxUSa9NxsDHwMIz1GBXGg7lsE+XhFY3Qc3kbOv7+jNfJuskw
EPWjQKQzDWEWOtHILKkpk02cX8tzKix5Hr754fC5mqCeLihnLDRO7A59To1iJhFoPQGGwDEVF+h8
lOikkPeiS6JtWD4sSQW3iv/8rRZc6Wwtdz9B3ch6KJOsup3XzanJGX0bevFVmnxbhULzpMNEoBs0
uAvEvqM13Wq2ikGWAOaTRy+tWVF3uOkOiUI/h1x8s9KUDJHmqBmOPnzYRUHRNxVzG5udiAM/ELuW
yAzPNbB8lEanvjZnWgf/d8aSYyRDe1nCw7wOJ+y7bdNnLUXHEEDABpfM0YoF9BC6ytoJZIrK4iZc
KPQAQtyAVogxEbwdHfb6SPno/dqJgIjBobT6zv7PrqHWZfAfh8IuinEORTWLRkVt0rq28Iv99dg2
KKqh6Dmaa5mMDQXDtzT/FBNOf6sYkQ/teeSXpfRUblD2otRCkgVAYJ11e3ysxyeR74HDv4qbBiGL
7lph+TvJ+QhujUWRFnvA9EeumFMB/XI2APRcPzgs1/1+YlS/6/DY6Ntx5UvRmtAn3bn/efL7IWCX
Hj5y7yRpdR5sK/kxrPphdoIP7My8SvIagff077POxyMH0T4vWKg6hAGuU2sYGwF3p8n8VzFyugTU
YN0K1vaIIUdR2KAzRJn2vjiFW0MEo3yrUKOfYobEV3Ff49Izr/x1uMUTGJOvgXf8ivAlrJB8FjDX
baZ0oETlfcoKl8qMxNs1V+JVKg7ptNeqM2ePa1MZcqd76JDvrLeJY9/6mhU2OwYSZLr0/5BBZcuv
AdAp1QCiFoFRDYpsJCnxWrb8jJ5Jp+BlWtmpUN7e1A1iHL/MzxrxZ6Ps2uWw8OztqveLUMfFQwxl
8rhEpoEjCHIWdRYqytLHJNXb6lNlQV5d+zz7KnTn0AZDniNjPCqZFmxIMyiKKHNuJUV6jYlQcbii
p//JVz1jylBc4+XiIQ7FT/GZh8tC7/hPCrH0WGg9YMNdwly0I1U66W5vrlMh2W81cOPzbKJACD+4
/RnGnDgsAMgNE4OmJUOg6Ek5UbA1hpZsuTtFvUDh+wIhvmn3C59kBNWyofE7uEXqNwqwLpJGdInd
7VDEec+vJDzxg7s0mcda2FTq/qD/D+tPKyDPAg8EUzAGk/r0icN+jrtof6d0NAzlJXp8Su8e/gbG
zcJkb7CLXmPqp/nqvoZ05g5VKy/M+PLAn5SRbm1xNnNXIY0jfqsUutkyCEd1b/rsOkwL1WMEY9lE
Me2kiHUm+Ht4/LKR9dbSZWqJSHbzEEI2fqoirDg8k7KgKq5okb7DhSqUcQdP+FIezVusoHsRL/vG
Aof6arPVeCrV4o7Slv36ydmDos+RCUAL16YJU9k0uFmc/Wmm+Dl4xbXNmiT+mshe9IoNO6xnxU3W
bpbU1k706RHO6Dk894l3nHpUTM08nWRTfB5+gfiNr6RqFOAVjd1xaKmARFSB9sz881Ksv+a8IJfP
B3cf+cqOAFgS7H5iej/7eCA8nkMpUZHK4Os1ULC9A9TOcQJLYXSOH4KhibNK3a7yqwO7qRxRQxLU
wtrxSbFR9zwlMZputTqM7O5u3bj+NziQGMtszqanaqultsmstCh4VVofFIjOqcVQlLaPzKz+T8wG
wlUeD7hcwvqShDFl7nqrTaVHI0rePU973i3l3F9Rl9kVAguiTd3H6GUJ/5tDvC6bmlHe53eNcgJx
t0x/RhM0srHt5yJOLxZYYiM3Tyfgdk432cyKUIJQWuNb5f/FjG8lqY2ZkAcA5zKNTanUwnyVH2Hd
CYnGvtEeQE0Qz1LBdTJUeYkORdiE3JJkfX+WOiuPNrQIJ21bmw2m1OZzvJCsGeDiSsVFm52ZXUkX
kcSghG+zQo0w1XhpM+6cRyL0wZPx02GYKVTPZXnIwApmbh1nPxh8cFDLP4LPgiM2d2cAhAnFxSLe
QB0jlKH5u0+i2Iqw6i/2BGvUUddvIwDI5kIGhN2+0E6CmGXIISLf3Oe+yfh4KoM7LC6BLLgf9p2t
rhqd2sFwBk4rJhL7PQ9G0hozKSeUh96/Yy3Lh+UOKt/ax4OUBAPFSWk6qg4VyQ+APZep7r3HGoHn
M2e4tKolR8ujr7jqSSH3Vbf38GFq/7LdJKOwnoxArfDaaxSYZxxjwkCbP96/5lzdokoB99DvDhHP
Jnx/iBHr1CU3+0SIjrYYx4rbIqSHFlElFtqq4ykV5qb0cK1e
`protect end_protected
