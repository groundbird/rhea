`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pTe7EdXE2zbFpfUjtTJwH3vrv0atBv1bftxlxIitt8BAzOuk2bxCaT+gZPyKL7j7A73DaP1L1OsX
8x0LWTaoGQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lxcG5iMkLXbcTWX8zFIk9TYEgBxL45bVCEHbUTV33ROoEr2OcwZLJizqJ6ebZTFjxLLFLqc0Lixw
SZDBuWwHBiTjQNxmoNRYKgVm+ceFv+Se50mly6S0vZ8lztQ+sWutcQUwGpxF4kDJQGxvp0/HGmsM
7ev/jPMuBecLBPZNJsA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DT2VmFqFOyGr+LijHk1kPrZWhQs4V1G41tR+giCaP7mS4dE/NqQ2opiQ4eGaCVckh0TOjdDxiCgr
vn0W1v9cf1D0vDeKgH+tpPXJtdTMF3cTkHWlFAWVYaleX5DyfXD4yyQbulAl6zsxDv/lMoraoIud
VNhd8xLrmA1v4Q3SJh610OPwmp+nbELVmZiTWb5te5Byis6AEg2DvMEE5/V+paZIw2qcBomKaPtl
KcjsmCzLpd8BLXpSrObIx8PqjN/I3Anh3zQfbsXFMc4oi17pUqe6fBEOql7uCH5Aec1QkzkajJWb
dsAlwghqY6xQFUFiZnP8MWX5v2xep32X9mJv3A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G6KlV6HvtD6+2v9BynlPK1rZ6OoRzMewUdzhMpM+DKJJ0NrZNABRCvT3tGqCnNqxElkSBDFSjAwe
9igC9extNsc1uKF5mMYvR8JRytp9P38p4wUa4F2GpfmgdN/GP2o917NIE6rwtUvFPT1MNOQCN8Mq
xvJokWsrA+FqK44UICs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a9OLsubH/wWNP+GydPktnO4vYeO2+BOnpq36+PF2n4Qupz3YXt3cCrPvdQx7ldQb7kWk9FGKHg/j
aWn8gjlMhEbkvPkzkzuEO5XQeF/tSSWjHLyHQMbwKihm8bZycrbf97S06Dp5wuGtlDqLqvzp/dGh
ynzPcjqGyVeZKhkv7yOQu9OI41EaIu3kzujU0pMjGtsZTTyqnQXRdMB7rHIIruAt6MeVCU4vO0/k
/n/Z0ZIsRlvi8Abu+4nOBIJSwUFbAFTsO1VJldhPwnw3+7Yaw+gxCJlURY5/yCLY+PLtzPjIk0/7
cZmffq85lKRZU/WZP12aeqLJD3iVNTAl6JOPWg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4384)
`protect data_block
dxQdY21Xb4VeBgom2blkosgOb0GvEqk6xxG/ZcUIleqX3U/u88AaHvAmxaltSjvZqQEpssElCSnc
rUi4I2m3swBW//IEke8jrln19BPCs00ZFX1Lo7/tennjivC3FrrC4b6/bFk98t61dR7d0lv6WuxC
/WsvuLS0Pprj4YB9lZS/ikk2jETidbfeGQOpVRPo4UPdYK8ZvyG4TOGPiVCDaqJYbjLkfzy1VMoT
aUVdUEkYNzyDe47ljE0MdZcYAJGtVCsmeXR5A0/T+MdiAp0AE50THbfdpZLrb2Ge6yWmfEI1dHtB
Eyh7u20jM1TM6z964XAGJKj1xMDv7iToZPnjV8HvBMhhFNH9SqV9QBNY/1xKj4/oIkWWKJadOL7S
4tnz5WTkXElwhVy18ug+bNThNjfRE0uOFzS6khgZoJWpbpw/Zpr/O9rRB+lToMJ1zbdbVP/AOeQo
utkEMU4tN5MKfQWFgq0PnxIB0GsV2SvLy5fKJ8cA3ux1lhQe/gv4ltE0+AE1Mh2GXrB7WKR0Ug4t
Y8OBiWOQYOw2jt4L7cdZMBV6TD0xEPUwjdlnM3oBZD4SW01r57TPIW3fLzSxuzw7NACeGhbwDVS6
yeu+ImAfvaN2Cs+SqnYjyUFWtM2eDBSlLcDJZGB1FHUZ19tT2xDnv+kNwWqibaVDTwnHYTDZM5FM
s+9oVFdn3GghKqPvAw7emgcQ77FyKbAmy7Xq4LRZBOtKixG4sJj0rcBSK/50WWKvy29tGAM5rfs/
0F+mLg696xAei7VJBEsTXh2B1IwAfEo9ja+gGiZbiBud1oIyJYqC83a8x6wjrB/A76dzLMnfNRGm
a9L2Od0Y7N5uzubtNPs/M17pNsTwy1873d3k5EF/B9jhXhMmoV1kDS/cD0v2X6xrdLwlr0y0eSXC
/XF8bxCRBCZwKEO/hEIQw1phndTHeszN46SZWjhtGMPGfPv+riJnIDeHWJIboi7Pc8hnz3l71aCM
mRwWaYLXNN6Q3zbCLCk7u6ugCU2PFVEqzxJKfiayL9tOGuog63H51fhiEqV5E0fhM1G7+AcXwZxl
a5SSd10BapySParBGxfmotLg5bNg5DpAWTLrmkSR1ldeE5C4xRKni6zFK2QBWKlb6jjVTN1QwaiX
y0G5Zr/k7HdvOY1CDUidsuY7ou+Hr9O7XU+vp/FzzIDStNl1AiijjDKOhR6Pu5B0wFhMCSD8lMON
lbtMySA/aNNBVAWurUvYZOcTTmZ6I/gIPiOqq/cof/aiEzmj0NlBN+2Lw8BjsmRWW1xO8L4wMF7H
Vz8X5tTOshqFJIZkps8u5rT4DO5Fk+MT84ULZUQJMVG/pMb4OMLNYb2Scr5rJNEJjneDljGjdJkS
D4jugdc+69d/UJEjzrd5PqnG0qUkCBG499B25SOK3pGi0KKUYfEMEOMu1GIkIJUyrN/Hm9SY8Lrr
TIu+YISkp6srm0SMdxjjTwy2I3AkuqfPpd3KIZo7Oe1TNH4rygIIXBa+hgAloIKJqcEFiTpOIBFh
YIBk1NXxGfYE4CyEoWNfHB5IAacccij35D6jGlPUnwwtwpMf7TqxEghG4oNWglaWi6k720dOcCHJ
07IoL1M9WbH+mvITl5w+tL8yMzsh0jIcIkZFxuExJJ7XSfn2W/v8h++DhwLzFD7jwADiRfekajNN
D7a5Hxx8WMg7TgA8a/JR8Doy/8sPkrXa34SK66KRDCr7FZmvNjbf6I19yzmwlCzB3N8hPE819Fsb
LAeSpOvkkHPLloYmZ4V93k6+wOkgCJ0tWims8YEFmxhOyeDeJVhxO2cyugyJE9bMP+kEvR5TpTaz
BQpIQCqubLEtcG1vhQm8fXJXUQ4itNjcKE/imv8T2Zm+zX3DiXQFbKz6lXG4ZR7OQ1r3UJiE+PUj
Cgl2fWk+fFlp11e/XaUM0lk7j1/qKchCIApNfwCjvRIE4/AiEAm80MNXVJ6iDWsflDcm9lrrg22C
FEsz+kyVbXuxIFBW0l+3BtM3PMc8pHhOF9ksaz3RDrsbqFABF3f7/hK05YGmu+p4u7eS3b5ry3FU
SAggvC/okNkHdzT31eDSKIUhFkmFv1FkTi70PeXwhvaWV9x6eQwuu0MqlGrAr5kNpzFZf1zYcJS3
jR8Z3DDuoR3GZRXpTvp4wLVPycFSmhoarIaZoGufkj7EgrZ/Uxp1e5CO+elBGNoNGGJtFxNGQTq0
KmiYRaM9h0olrqOeD6aQ2mXgWh3U/oXIW6IitoaMVzZvGS03awRpf61N0qewUMVewFWdqJIxeD2W
nZMQCTscIT5FC6n9yIW0KNy3zZ6rMIkUTh0b82/sFS6GvwpFxoiNtWOOMgpEN0njs/SNOQRssm9X
55pkMk4HNzK1wrp0WYrUwRkCftqECm4yjjsq3cnTE71wNPRSyCK6zOU4/vVQoC+7WRnCStppmRpZ
GAvxQjm0Dz0Yd8bYHV8Wr7B2q8ZIwDeappuWfx4H1L8RqVM2cvtqXPId7N3asQ1CU5kLD3l3v13h
T6xEqvXUZiN6FWFnBa2ilYeFpBruc8MYHDW+ezO6LUl18jolmUvXQFEVbC3fXROleq3o7GRuZmTu
/nR2nG6Jus4oXt3zqWuttVMHYBfZWvYFiJXdAW7XLh3psbTL88c8gi7H1JQYUnGuRTh0HsC+039z
o1+47S48G7f8HUB+tyG0dsuxXOgTQTFgfwXP1ykFFvuQXM7Mrdh0NubV+Iy8L2qCzXE+yVljLnYD
lxsOKTAll9FPzV2GtyMY92MoikJTjXXy41LUCn3SKPRL+cCyOkNXImv98OufoyiysvvvsECnUb68
x5OtkbwUk9c40OId3AK5HTvf7o9A2HwrMgCrLH0kwbN5Yg9JZnKNeunhXfitKaZNrVxKXRDy+v3L
PUXnHvAES77BKwPXD4CTp1Ebe+8qzc2TnBfxWOhwvpF6iN69O2sL4tPm76Y8i/5ME9M/ZEef2aO9
HYTEC0vfkODb2zPBzMnw3iyU06NcuO/NeIhmk3ldOuf3arcGd4wwiIdRvWo+e7KqpDHDY91QJAIx
mk1jKgPgxjnkIIgjN6EeoZ6teNc9g2Mns9JGkRCQegKk2QbLk+vKcJoCd2bFFHeKrX0qcx35asDa
on+delsGK2gLGoYvXZn7gCzLY7982HqXjWTl42ugLeoADpMmQjwgW4WczH7q+oB8is0SesleLfB6
B/rKqC9z36HNkV7Avv8JAx7MK8ctYNIuDeJZXJ0PnHsqGGr6dxS29Yk95XH5l1dKCrastDXZMv3D
7R1peAvTNkLRNKRbO9FbqnIc9ec1SPV/SNjCDP5sc/uMxUA6a6mX+y/tQXrdhLQT675J/k+3FjPq
IU517dnAzH8sxx4Eyat6V9zRTiPHbxg9v49crF2G0XOQO+k+WCzvki/5OrqKqdasON7xwcFnJeju
v3WLNab5gGSQMK9Q0ttiJqdZBF8Xunwe/sBHTXnddj/NZf/FVYsvKzEUoGfPKxaZLNX66gkeT5Rc
2h+I/uz9m9QiYG7TdxKfbK2QKrQQeaowTZJV80oZY+r0CW2Sf2C/dBwLf4dkjnaJhBhi2cmIEPxw
xvUB5dzmlRZobqVPb4vFjoOy30TJEzv67J0e+h+6mU/sUhPBAWCudmjxSXmxGbwVjspzIo7bHxNl
PEbaA/sL1XAGmXO3B5PNTILkY9GgHoafgNics2iEBfm7o+/pedAHmcB3z8NWRhM7vovPVV9gqXVF
K6GVeAf/FV1xaF/CZSpFHy6Gv8XhRIpoBGpvYkwbYzAAORmXIHMDS25c4AADPDZByicxXl4O30IK
BCkDKWCUCp39Xf8sb+06KBUHVOm+zJZYKfbywEqF6SmhPmOXBArMkyvZ3DmlQ9MjZjCE8L9qJkbB
jJavLcrV3tEoabdFD8aG92dclL1HFLpxgdHLJjt7zd5HBD6sj6Kd4xwqSOQaztxl/aIYGanQKpea
Z0cdDKjzR2nI+zvyKoN3ERMom45JJrWqHbkHZTVaIUSrVxTFwSH2qtpysXKbHL58aIOBXgidxR3Q
57OI9EJlJkk9ugjVdsphyAhmZlEJ2cRrHogZbnP9Fd5OFVc2spO05ogEe6ohvQWMOVfIKiwpmSxY
s90VB+zcsJke6ntrBVtnmR4MySadcoZ+prR0Xq8i+Z5w5BMAB++/3Rt+1T8loHMu5Vuh0u9U0Zow
k1scZ6MASFN237aGfQWXH6SCPrzsAjIfm1Kpkj19VPgCND5RZd4mbvmb5bOuKvfTDq+QW7DjVtr/
n3ynoV1PE3aSG06hZw6SjlqIZtQ67N/Cg1JADk8W8qf4tEh0sj7oEik0E5LaAYFzl8FraBG/ZsTH
6cKEArs/f59fApmG+Yefw+h2RgONmM0avUkqYMW2cEJ/qMeGfdushRbeYho5k33i3FIg5kBo6mBo
/SJLYq3PpclDabKcWAVP6p8TPBjKel2Z3mOmR9tQfUZuAK7oRmkwy4xW0XrC2SXY1sktbzzNBpt1
9MQGIeKLQOHpskF8kdKZxsCYpM1mBxSvH+ULnBvyfIRhfGPV4oryZtI43ZX0bYTrxIQ+hDFXreIG
dR2TY5meSvDYvMbcaVEiq4ZxmLS83PkZEFn2rtQV2r90GsPtYqK/nADKsqc8c5MapKdNskuhZWDT
qQJWsrysaAe7SSyImv5/iIjRCUOOCvBFitWIKoOaJLX9DsJQ/wlIgCu5UoTjycHIOOwbsnD+jVDw
h/NA0y83P2Ja3cpzzy7SRdrg+UTjDVdYa9Lv8MbSs+67RxMDrYcjwgawVP0y9Knt1NqCUlXw9saa
mtgz+JDg2j0rQhAskIX1xghiJxvPL2AtfD2peRXHScTG9QqrRx4oFIMCnrI5DyBU0nfNyB5T0SWV
J/zt/z6y0cFkxDWLU2BSdfQSSsBP2rmHmm1MpqcpL9fjZ0fKMDtK9dgmTREikRGFmauT8OQHSHEH
YnLuVMlJRC/wqbqUfq0wuPKLK03VIWd86dEQdE5IzpH1x187HrBITBLEAvrWh/wAB85U8itlrPH0
0qbwHT+KdtvW4e8xJ1E5xE4CMt8V47DxnjMd9Kp8fHRhBZLcDYRM+kne0xINPAghowIxU3oQgMgU
lrfWdqLBHB6/f6+uRfzMJ+SNUxI5WaoBKQeh1M9yto/N0d0XvrEU0/8woLqfIHeO6TrhS7qPda67
w4kBArdlxM2if2fh4HdL9K2XZ8/hRbg0geXehwbkHxXfpM0V/PwAwuTyMOdzgyd88b/kdb7zkuQD
KMZs85emFo/O3mq8pTukpICq3TLjBLjl6kCG52dTZI9lJNH3pnLLj+Ggl7MZ6pdKtgUHjRFfP2bN
SnolBYujt67LoM9BrXDJwR4b8OsjS+R6EWcHFXORLyGdpuesDMO84nZhB5FAKvrknfmm/4rb/ipw
VZws2qQEi9n6THmJCfwFiQ4BML0JNNvFUyJXSMymkKSaJk2r6CJrSkgdXYWWktA9MfFXYEPvdZyr
7ZwHBpnA+teBZ1Ra9ZRzlM7VMoj1u7wny4ExqRpltHOFTs4j6XlqIg4LNoOhjBTSRXzr2urc7yxF
XrNy6I4/Izz6ZHWEtBk9COSRT8kbSY7a5/mMtJYbZSdYUQK2I0z1MMDdSEOopXrZ3EnJhiQPQ01n
z4L/CH139103MbQh7asMYXch1tq+qR9KHjuNBveOPPLWIc6om3a6XQAWq5wT4RPgKdJRaUUpsJTG
xcxX5NxjsiQs7I+PB0Kz4/kd8fEz77Cj2URMNiWzWsQr2wR0fgB+AaENL++jKet+eOFc6nVZSSGo
ma2dI4YyTdx3vUpIVYao2RYREO10sUtVNdQHVphTdurpBaSIccc+12eMfYvtBXa0kH7wyw==
`protect end_protected
