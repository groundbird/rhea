`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Tjf29iORrKVIHRvtvrk6aRDqmKeJWaLqE1aCHIa7FYxGytOGulU9GnP+DRN4Ow5dJ6Jp1iyZrjQe
ymvaTXXJjw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgpyy3TPo/idL0RHeTQR/rQJdwyhIO43/HQrJDFJpWqO8q7ttJuy2ZlTHW9q9LrmnqRRiWbW2Irg
QsFxHg/47mjvd89BDzQBpdvWkTwG3IGn6k/sbFF2v6BUfI6WdylkjhKIJXbedVukWBl68vW/I4Rj
bk+yAuO7cmWdc3a3Fuk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zl+eTIIpOqO4rV11m9bG45TodRndMR97jnZCKF2wNgWgUqthyc0QOqR8l5fesrSfQFmldkdI4Aof
Jf4DME2EaDxN9G2zq+VgK0o711fQ7DkW2J15l+qhDYa0cITKyqrvJWd/Li+FqLz0tefkpN72tBOm
sjbQypImXMtkGCRSM01mz0vvzRseJo4OXyjBk9KP69bDSB8Iiz/KmpgbH1TiekFd5o9bci6/SxGA
WOOdpTTlPk9Qz00l3OigR8SoIfCUUQTkIyhdjqHmMEW9Ug80lKUNz+xIidgrKiNFezYMx0KUHMKP
Unri2OeUgvaFgsZL9EnMNbIyPKaloqHHuC64Wg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sVFqhKafThpN3kYCJZc3USKnwjYfeMNcG9MlLTuMpwNgdcpouFKfXxycRcYhL6K19lHY5TOol4z5
sYHEZ0JPgNjzZY+6q3g+kc9yVP+rLv97IDFczDE4lyAjLpuj7AdTpQDl4DS14M2VmZ0vp/bp4vdH
g4KvtccX/Au7XWYNjjc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rqUTz6rDUDK4KRpsno9a+KOnh37IXTSclFTnVTGDj5ZZGO/4vKjZsLvOVQVi0jrv2scezLOZMHAF
kA2z8eT58BkjPHwGLyPXbfKGaiHxE/Kd/dGXltHrhDGc3mlJPK7oE+EWVwV+i9aSYzHuMPs1hNuY
GJbWOTMjVIHYjrlCfoJeBYQ67yqE8LV0IJYav9EIOo9n7hqx/OEJEW6sAUxsOIznQJ4NcmLky8hu
KX9SOkCSjltdPQhqeFEr1YoVz0z9RfCgr3a+6gZMEGL8lOwvvMyOJ8ALuZPPfC3m8xX+zv0OX89U
45DdRmgwSZgkjxY0Qjah8z+eFyW8r5ZVZ1+rnA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4608)
`protect data_block
e1EimmuGN5zoP9EctaLn571RCwJyBz9HgJCBbxOQvUstFbb3JBdijUveGmEYaeznGjvnGI8WT6qA
pY52EGkx29AHCVtp46bDDJTzEceyaMQ5Q3iQ2NHeUbfd8e6LMzbq6GlqS+caMyf/iqg240TNiAvT
444NxbDHlfSSVBFJje95uszSi5JBGkFsuby5Bu5ynYrpXYhlvo32/F27wdgexQ4edUnel0YvHauJ
imn257XtRGHUSb7tIP1K5XICAo9gnR0qni+zzcEOGHrPb5cFdD1zwOVuu8suyb6U5gp+TawgDhkg
xeu9q/zuxoLKdaf9z8JwEZnOeAgkGyEylxZfYtxXddF9KtYVmJuPqfYX1Fgh7BtnSOu42xcn4qO6
0rJio/5gxEiFEe08iXchE9io/8tnpwVksS6lndlsIPNDm1Eq+ywDuyapl7C5t/2FTAODrnoXrPux
g4s+aaVtw8E/UUX2MnRki26kVWdeRUrj9Tr2ek+WJ2AdPewA+CMg7G3x1FrcBftGIsVkbZ1Zpy0P
vzk7FVHhaDRJJsEB1m6ls2tnp2/dfdDy4gbA+sANM793Q8D3rVBHe/TyJKB/DauSBL4BMMe6kmkC
dzsgs1CZGwx1WPbM0FBHl5mGg2L313K8bMoxCzcFXhtEuJbmxS5HwzZsGsP+c49+N+CV6HS4Zm08
lY8qafSuyhEEfjxtnGyjDrjNl2FJCeex+T4qzix19bBomQrUX454m3YPOGdTo6iIyNuTgP67UNYc
XCqGtZj+bDcSCU6bXhz33x0QvO/VTaQHbHm2ODC6cGHenMLg4agYsp5AuD3RVkDKaapHijw9NRef
QYfBQSml0FlwoBkps2akqKMIUrd0JYM7QfRgalTy4KrJnstxGFEpY9iqLlkt6Iuq/UZsvSUg9jB/
eye4R7YEcbWmIQjmtotKp80kQoArcR1sn7cTrpQfjEE+x/5l3b/zFBEyE6DMJ89Wjfo3OoZagl+O
H3HK422Kz4i62mRYYgFpGkMd98z8uS9iFRRvX0mRpZVt5ZDl0JgJrOJaqrpPfbcXH53KSuXWsUKk
iX+uFAXjZnCorOTcr7NUE2nFk2I8E1Zq0xqyFK0g5v1UpcX8mUZ9qqvcQBqVXFgwLERAgFwZOyXT
uVOdFA7CHtfJ0fhjh2+Vw4eCKySnE8FoGn6Jdb6WHyXh0rH86+vprSkoKs7gX8eslMcLZ0z/j0Fv
RmuW5y1Lzeu7lu5S6sK6d99DFWVXI3GsqpPz/giH0s7INESFWIcTXbT5X740cIHV4pvMjNO1lAfj
yZ3YWQwzmVaZTCQlLCaUedcvWObtr+NCvMMGDDsZb9zNTicL0FF4OqvUtE4tbQ8v7RJfKzXR8rDV
f9Mha4B6ax4eEam94TMjpbaGXUTZZ0vjeLc9jXehE/tp2ZUgozwQOgnyNvMUKmsYAllqv2TyCsgR
nvxS/Kxks8Bruz4H0Vudiui1MceeNpjU5bnY7mno1TRg8oqJSZ/l2kH1gM+ktTCjsC9eblUg1wKt
taYsRjf850nbatdUeNa5UnEKxs4A5deB4/3k6I5hhsLpzdAonuRHvP2WJchMHmsPWM259hakwlzA
8zlzwznTSclDAISKumj1LOURR0xtltFHXdd0rHExFyjkOTvUQTEtSQeKPt0efns54JQ58RXOYW43
OTU1RQIpOKCR6Q/dZJgvb/cTTThAuXTNkjiDK3wXDnuP9wI9cDyFEGeJZGtNI5GtfetfNDCO/WaD
2HJo8neHFHwlybMCqo3oQKVhAQKU25oEj0kBvhkN/oa1dkVTPinXjWv5PDOX/Pk0lwXNuCkpxHzM
lmu/qhJbimNneObvpth8v3gudyPMfpgtckIPENuiNcZTbEhSFpZCh1oQbM8PpsrZFpMKqA+T6Kmo
2jQ/ACg+61EweWRKcKKYlpMxnjo73D/k4LnFQWjgTOArtfi3A1mE0YjN3+w2ukB9WH77YUciI8pj
8yBcx3fmSqgUISJcrCGChIzQLbytiORa6fuiVb0/JFYnNUd31ppV9QNfoAEF0HBCZL7Xru/q8Oe9
404RMDowYt3H9py8YQlzUIa+mRgSxNmpvqumO2WkMeMFckuLa2XheY4VAogaobZpGF5SGo+qOL5u
UjCIB+QtdtXxX+wlK5R8qB0x/E/PBSy9BXvod896YtxeI224T0aQialse4NoonvVjxgcHP+hK6dG
O2iLPfizJofcw/p6SQDg6Hrnd0ZsW8t/Ez8RbEfqynpp9JahX4kM+PhoG6OXtWHV/R9DAX8J2vLo
tNxahLeCWs3pVelBIFPVOWIIePSjUrwzNXsaPgeKVOTTJ6RR4f/t/0sdoqvPPgDcpGCAQbLD73RX
Cn1ivpZ2eXfJ0Eh9JmYfGrjtr4K2B6YCs75foFexIpOG7u4/xsOIK/DeXRU9qUJOcq5M9clM/Ohp
TuV2LAc5EXRjg+Za3GCbGsUPfhikdO3LsqkFG+3hQm4aDPA+rftFhR9473KtsbMM+KiQrD9rGAw6
ZOpt4VzLw72euNVQlxq9NYsm+JN3McucEPviDyS2JK+BxMyISNx5hUoVkLBVosDa/H58tLxp94AO
If0aNI1EHVaU8k8UxYg2xPe5HrtfC3WIGhunTSvneg3bQmR+YOOPt8XbiecTETGMvW1XNFvT7ZJM
HkJ2EMN84KlACoA3pX5atfjGDiFnEXkqIjoOgriQHy4yHh8Y4AnAI2SDOEO/z8oMOsAIjVWONjAU
jE8jGPwmXXJdFQJN/w0TaydAd0zmwjQBMHYVj1WJRfmjcPMRkWxcis4l3/gcYBILPD3hDzZRGugq
RpMLcVRjG51u8LwQRN+g+hadR2CNqpsl3Eiv8gtLitIVpy5n1hR4yQRl42wDIXjwQVzRbL4SY4Z8
iilclqQ6RH4yv+bMGHWL+ALlJKs+Mc7WszZ4FdrmePFOYx5pIny2+gJlfTZOhw+Sa3HcUxXlXjUK
X43Rg2egbT9FGJE2Sm3aNyS+GXQlnPnyQ8SQ/6ji+DpsSuqt9KZOn+ayy2qEKY53HK7hurGdQsFR
BaXURaHAINbXu0/S3MtMIbDOwrqmHeGyEBxgJXf9+iUik40ZbjrsXszphpicxXY43bBK3uZ8NPpx
sjTlxvSns/TeUtUFL3RcwyY4srCTtmRZEYYTz1x8XOmUSHFOj8k93JbypXd5e+G3sEVXXDlDQMGC
TWGeiMkndbPnAg4lhJ0YPrKjRNq5JrfCM5b2MIigs6pR0UnX/ffggGdUMEwm7yjTQ2BbRNPZ8Mg1
zO4jPW1mHfKMcCPhxh8I9G7CUk8Ra+awavlXzJwSAJYJgWPclE1bfEaw2BnQLewNxvNGkFV5WFSl
mhpZuZA3A/WPvRfy84e0pBocjWkJzw+MAyQU63CKfeTbXcNa3pNqTZ/sdjlLhrtiwqElWsDPQwwz
Xypyirg6YzNOdXkYh+e7sQ9Cw4Ar2XnTymL7oeDvp1UtdYXohkxLOepzdk1eX1QO2UCrLC0BbWZg
tOxjfg/5Eq/mPLhnsPW3pzX+d48ybUCz6AtiVMdSMh3ErWw56NxNsQZT0poNJCqLEo3di+BoQRP1
IqhiGpdz/nS0svVuAFD231gJVUap0s0Jb6f8sQTVTedzzWvpi2F4z/1RdNnjpEJp1gnypPr0Ao4G
Ju5e6R33xfQtoFOOcBZvb+IS5FGeD+24Vek+c400JXcnq0DRWO+qGqk9qWjCIPvPzLmiggSPaKk9
pHkLFgn1klcds4xQ9ENfhvTvhOpHfPycSnprUZt7bUfc3LBibFPyxsNb1TWq8KbxPxuhIBpghwfq
N0DFwPJgFscM5KplIbveakZIfErYFH/idPV6pR9fH8Nk4j961VxlFePi/P0Uih9rrOo86/azdEaU
Jf/CUZvTagOhVZUy08we3wVtrTK9dIXZA7y+eadcvwlxcIeQ7Pb+GipgjDVhoWvHYvYQ4c7yYrhc
uXK2LJ7c5UzGhhnG3+KQaK2pfyQBBoFWbse0fHce4bk1hXWtlaiOpohkvDEfjXWhtg+SBLSYtWL3
9jltAVYBWkJjAej3FmpPmguzOvWfZsH4qJbP4tLyYC1vHpBrMkyqH0w8NDNArFmzqW/hNhzDwyxB
EbZEtLs+qfvJaPDWx5i6a+yVNskwrf1szX2DDyIMCmKiowriYQXRfLJai8zWcxyncXY+TNKbeUO5
s1uKgDVZgFFIXRAStS27qCdJujL8pDiEiAStCUElvosp14D6KGrHmWesLcfGpUE9uLjvcm8EacOj
IdLHpxmEW+7EqJZpBA0H3rsyJrDQ9wplSh4F4QgFlSJfog+T+19WVgcEFh61jw1klq8JtGYNWcj/
fBucDE8WvomL8+y7jzG6X1/tZx+8nXXUMXxiWcoa9H1vbvVLmd01jBjm7qulQ4KW0ueWZ4UCSCsy
iJbzVtbm0L2UvrZYga5X64Vwyu12grE0S/KZrP2WeINs4xg8+AcYvZ8/J+2HSQwk1CDLt+Wwxcv/
Rew61K/ecCFpRJ8zSxkob/2z31DSoSM+Aqf9MBMCHYtzAd6M7q8tab6FZISKCytNVbE1v4ehGk84
gvlLtmozlT+xN/F2aVpdqbl9mGJ+xaDefODmM4X8GfFRuGGQ6IXy7/bNwDqWOdZZNXl1Bm4+E87S
NcqB+NZl9gydkeECqjXTbgVxIpfX1YkWS6FKcMsnOj/tOSD2PIMsBesG7/Esv1pKegUbxAOLEqLI
GCPJZSc9LvmOj0cb6aV4689YpQyUrjlE5vf3RlHp9MKLWOcsfIpeto9fNpdP0McyNyVukX+j+/iq
CxCkth++IHUJRB/igqyCpGX+nk/EIOZQoxui3Qu2Vge6VA1sLte0FhtO58cTrXz1tli0RSjEfFsK
wkSLRHTLX4x8ujTSSdPh4wzqMtBcxfGUSEri6vgtINF/N1gfvjUu2eehZhoVOPcBYmRb6pwvY7Hd
gtrCrT5KkZ9di8rj66HIivPrpJWvvlJJ9Qpq/m5D4w0Rv4162lrR0qxKZ7H0HYf3Smw85GPVEvTj
VNcxNjVU8BZKnNGWdwjDyVLbfVhByR9RCrCLBP+c5kxCfZw7sWpy75yfJIYtJU2nMPo/xnGLwVFW
JWXUjVM1SMD6qXlJqa26UJz/SzmLmKaZ3qkATxTMCum/kPQ2ySWFXzs5zUfUSWGFjoygtlLhe09m
1dCjcVsxs65jInArh2sayZeAPCP7zGPiid2gkzqtyNeuZX3WZLhfc2pRHzgnsrhQpa5yIMapzJnJ
1HKCDOctpPResunlPs8ug3QtuyQOnOMz3qFudohsV/ImSa8eESGipifYWczc3QJgf3Yj5sBT5aIs
b6JxfY2X/tgLyWHJMmaQyhGVGcaJ1Xdhlf5rvxiuWzlV+oCRtsFlEaOk2b8RD0cFAATC2pdP7Tlr
Pucn+mkPDm3yW/C2eUjN+SGJ1P+s+KjAJi5MfhhLBrrZHzVU7v2ltBj2rz9ald8yI9cwfRf+fTU8
3DDhxWKnyHD9clnnqMN43M9QwGRdBL7LK162JO+oNZ+QVlOeaNdwvwgl5SV/UcLi25B3WJZIOtC7
2dDob5mrNVlDr9WGXzTyAbrV6NUDyk9t7mJd+jF24n7M8CBWEkGtPP7yl/NIebKhK/3j4Pzq8doK
FNTzKnHNvXepQUj9G4w9lVLGimMjont6aKb1xi8NOzkkokN0Q7A/qjtL3Mv0pAoH2vyIbcbJp1IS
b4OB3hN9zibA67hLQSXsftu1tsE2le/1Z+ntpcKROrTbiFTSzZDWOCZby48llKH+ForXbl7UxOxw
5O825PWH84qzTYcU/vxKflnYhVUqc4/QPvQ3tfFGsNxPUTwL7e1rO3NiTpgm2V2nWwJ/klx7Bev8
E9E8Zzv/wvfry3ZyVrqvKkLKePXhgyKkrk3tL9kq/GBcc+QOPS4Ki31mdlO294dmS5BqJ5+B2Z3E
KsHSFb1lHAohEj3cbe5brVII/PAm6zSYm+MwWvAPFaFQ2JRKtduOHZleAtIgdJRDzNKqrVmkJE+v
h9koMhkMOpnGpRBLirp7ZjdGqWinKQa5lNWJ03EysS3pzG/elAK2aZjKrZG4J4jIiBF541YlwZCQ
wSUbem/uPGQw/g9Xfnc0IFumbFAFcmQWbKQbtq7lcV5lpGAZPJsXDpt6HwuavVTU
`protect end_protected
