`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NYkQi5kVVvgHTTD8Ugw4HEkVLa2fTs0B5rSLL5OLX1XzrgAht/vTG1nIL/aAlHgyBIJns/j9QIni
avdLPKkseQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HsDpfx7ao5hgyYj9/oxnZ+wHlfhu07UHY6semw9Ms17hNIb2DyYGZ+JjjCMt6Bpsf9rQR76SpTNZ
w9zpuBYj/JzQBR7vVrk19ZZqdZGBHS3F3ZBTJ3tnAA8etgEHO1wYHa0X2vJ8codLogJ56f7sgppd
GfOLA4fMmssuOK5MYiE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hNo5aozyYVUTb2dIYHnLT2R0W/7vD3YjCLn0MjSEjkEMr/XME8IWjSOiL0pF5UJ1iazugMVYSUUT
7G3qVkMD+1WLm/DbWCBUl+0YE36nHReN2u2LcJmzoWg524T++h6gMZ5luNKoSDaQoE1BGTHi45sT
rI1sSuTRigLG025d8bF7xZcGXFsxoxjzbfbCAYRi+uWtaP9P1R/iSWVrJWzpbzSw0CMfdFTNK8vE
GV+ek/CXph2Ou99cgVZ4XOa1Up04wxAA9LH8SoO2cbzoKk1p7Z+dJ5YM7NybemTDClk36kOYoWAv
nBaj2m5xmRZhSdjTwc8nqV/3GrXw6tIoxBQeGQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z+WuLbm+998WNnvoDJGq+BYvy8iy/n/2ZYTDsiM3OcZQdYTBxqVyKG6mBgVyBQJT6TFoDM6O7Dg1
aJO21ElnnDbArTzeUhFEoLNZ1nmLIuBZ93Di40Xiy+piefNi+iH6NC1xJiqmLaPDa22SLlK+FNCS
WWgLsaH9rUKMxs1H2HI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b/vY4LiEdyGWFH4aohsD8SMKOP33IDQya6qlZ6UQPHahB5w6UsKIjq2Uv5TrmHHRlCsiI96ZSqpI
3+t6zKWiGxEZ7CQ7w7OlPRnAVMa3GsLBLslvFij5zNYQhbxrW8n/6NL8omBB9vXKAMyew5GBiA6y
4Jals2kK5DgziHKOONKjGnqBP+5lG2xr27pyiGAzyvFyMT1oYOgLJZzuFwF0DW4XI6yyQipv2+zg
OQEbhIHtI+VwYsQH8dPWhOOv8MQ0dckz25F6VMKmhKaufKgjessk6dTZk85CMg8TULbfHtXrJD8T
PlnCfYY1qy+w+5r38DRITpd8y54//d52DgV+fA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14272)
`protect data_block
OtzBzyrXgZ7FqJOUg+CDokWPcN06JszowKhZAVfv2cRuCOgSy0LVcg8HwhdJ5+qS+L/q5x43LUWO
KW0kKxze0OAPodO7PxpkFKzl0sb5LMJtDzpuO/uftXKiC5DraxCWnM7/znLY0XraVwqCB8QXbgcG
aq6kBw8pZ+plAXmaQX2dlYNqThE+R3EzjGqvuu5fpBHmvfw1m6jmFI8puL7/GCNVjU9ZI1/CMK7A
Y55SZ1iCDSB6ebrXgRyMPEZLCIensAkNZ5/mlpiM7BkWjBWNZTyhNcKiBEKM5no5hlbh/ivoV7h8
7CNY/117VZe+AAMFX+Gp8+6u9Y2HhrMjMPzP5iQgu5eezoAle0A1HukHrlolUEOsEC9Tiz0TeThU
aD9iorqks7cunUOsWpv2GKucbowNsJTq3CzEDv/S/Aca42fXWr6fX8nB34imszooDcCWnCQVk3mq
gSLQlJ4+Q5uk+WQDiEnSIsGHn40Nz9NNDPW59MXEiQ98j5Ax76IiSLcxyXJVAc8z9v0wasyWa+k8
WIuYKG8h/FsJukZpRqLRgDK8p34XVCkMASOzbjPUAexLoBfceFn0zZDuG0ZmMWZQZmcpjvY7QtCg
g6qOT0znenIf7v0mxpmDEgz52tWXThImH+vhq/MxjKjBKB/ZDV0Hs1NQ/5w25XCV4rLuPMioABSD
STeMeyYDnjoTeNDXmjQJttnnOILjtYSNaldPrbSasWg0LBdPiNNlvja2/it7WTVV6L37BiuWoqve
QivYPr9fbtHAZS542SsbzsAN7AtynIOFF3qSvPAqFIWo0nofVHszCC3fLoIZlk9LlxCZWkS0YTEk
fckz1b7LP8RhfiexC268hXv+2Dmi+Up1x3mmOl0aNqBufIIHdvljcaPOwK+TTCpERfpjWxtn2xCQ
CJOTAUIZAQf9YXKtFCd/greTuvnVhkADJU+5H5rSKQ5VVM1q431JXHONOqDg7qk5u18ASZKGk7kH
kd4iuxPK6cFvzB1FnG1VCAc53DnXSfu5+cEsvmZx0Y7EwA9kz5TBQoskNqI3AYl4cmrpc3mcLTE0
refZKlz9nP36x9DxkO7WdYL9qRI5PNqpYgu/xQqujmWxuwd96g6HqalxP9kj4b9witGH9wu1clpH
lE2Hq4iH2jF2bP6b2cdVyfH87qNLh/iMA2BytUYMNU7iEAdPHGuRwqMmQFXesyh5wR3JPio9c83S
BDKUNCN1zUvFRkdcqXANpYIxsbOp8oWV+96WUe8G4WNj8XWyebZKMRfEI0WBQ9+V8lRnXlEUGfUZ
lmwQfAwqNCwiynEhj8q+00/1A2X9phPOBjJXhHfrBxn1K9cbVkpVcA7Qix+5wyXegoeZtMnIugAa
QoE2wZYADEAcRe2wITpNV3BSO6dR/k1tBEQV9A1sY4W75hbPVcOBqvc40+04fXYCdbJR3ePrrD8c
KqGCFgiKYC69IuAZXVdOGiuJkpM867gaCZsDpDfL2Xnmng91z6n7/4CEmZNUeXLJEHTCXPwBFsu7
y+VUNRqfHKSvCLQiRvPVwDLKER7luxhRGbfEO1UPlKpdScONbu0whkpb0Dwk4Yx5Pl2hs1mz7ngU
3GtogdEnADsb5VBVckeJ7UE9snALU1RXYvOcaC/aYZcgEpyA9Rw8cMNGqd7s4QNqhFd/xqJY9xy5
sw1HSTHhmP3wEVqzirKMbt0OSY4DL4S2+u8oAPHmtzHBXVl+PwTH57l964oimLcPyILsBhHIYOVq
7dH68YvuNWFk/FcmjjUjuLMOrizAOfoAhRZn/Fn4MwnOWjHn2oruDHPmpQojcihaEiLrYj+SB4Nd
TCTAFsP5BbBGeODOYj78Wdd/NbiWOGJAJgxk/q3S5/rEejMoG9OrmJ8hmj7j3eexqlKdhXBPIDpE
mF1h3mKRQUp4AX47GVcgy/XU7gO+KE3DQTT9oGPv33WjqMHL7rbBseivzAZVKxLvD3QRRFSkF3Eh
QXBnsCBLfwJzzz8xazxpggjJ1FKCzK47Su1kNAml8ienkjP4x83e3C4w5+8iv3vnidPtAB2i4FAy
WCtYuFt1DtwF5M4mb4Uavd6zIvmWJXBB6gTsP4Vp7KMkAbVr9d5uwITgWheQ6VZO3dzWDLKtxDJ+
XHbGWqYdLQx+sgalzBXVVDZiYGNwx3fT6Jn4yOhUv6TSpP+5EI2dkiNKYAMsmMGKjtm+XxUWiw42
KymB/BgQ8yI9K5JEsqrDvtQlIEPI7UNnUsGfuNTBc0BdwoPozBcfjJnaiGxPkQR5Zv5yw3qykoXg
jSpAtjW51nctit9z/DiLMimuV5ot8lDQtSrM30azamBldLabPUaFe9VvP3UuKPVz9SA6cv28eBFc
RT0DI8Ksy++VKoFaKgFtaxIqaUaEh679VDSuSLLxnZHd1P7vgIdbAQyLMrHBBYwG2rSMYVSf2q5H
QB4oYQ4RQ19kCJX1BLbjQTA5eyF/iDjDZ4HkNtlQxCoLjcWkeNJtehJcitUKCoiEDYcop1r3YdPq
bsd+O+5LZ3vVD7OZttrKFGTdB0PYHHgI72VxjOd39gsThPF2bfZ3WM+96qldX8gniN2v3raJC8Dw
QzKTrN26s9kOE4r7Bn422Ymt8x0Fn1T66dBsVzKv4WJB+Se+i5F2AHa8X4SMkCmDADDcolXm9/zJ
PPX5MSw8ZSGEGHqOIgf/trNYJZVfdMWdrAIg6Ep1D2Z2NIop2KAb7+xfCze/neL/eBl67yjtI+Qy
xoopwvSjjJgI6WyOSgq7PuZiGEhnOt5dIn5b/hd5bam7eLrZKi3/G9KD7LQj9J/eC8YVtfCaSV1q
4sqTHZDXW8suXFGk80H+xGtAM2wqsrFSwP2v+v5Kd3VKH9mIxajhQF2JTTuJtsbc/TLEHnRtPAaY
p+O+Yu/6LQk80D+qGLhI9ThKbpZJL5g6UZ5naCqcpgCVM8IbwQohcoWLcYZ277jKGQiz5kaksid7
VW34CU3selD6DSSHzk95Brtr0j9QObHWhTrZ+vmRPFfuSa0bl5j4PhWKaC1dltqr6NL9f+Uv/K9m
ORnIqmSkxW3csJrxRivDLaPkW89wMKofbPzRShwffPy30LSq4KUPiXC0Y6TFJYz1qBQu/jBiyJC9
7tdykGECUsGvXekXkBy8ttSI0yiIqKDZr/hUqsdLgIRXtQtd6GMPEljRg0sF8ts9JyLhsIyWfxnu
wnGIqxIbnrdcIG8/O/M0LmHNhKUCHon9NraK3cBbjg3Z/Mx9t7g9VkGS9+vRuKpxaCTEIN+24shE
Gtx5lajXfulBHrIRcNsWmJyJucKfTsFSVWAHSmlUMzD0wULaepPHBRUTq+ZBbb4thmKP0CX4zQq3
9fJnLNVJJADnY5Ng16MAJBCZULxsKwsiv4MRECuhcOU879R1bfJGhHoo4WyAsHVu64X9ylY9+s7k
g8F2FhkQkuJzlgL7hhvPV7X0ij+L8X8PKYW6C7fWGcuk7uf6Nuf9s8/sOwy0efjCGHXyk2TvgOFd
OBnS5Et4O8B87ZGLaYUIPr2IBSoJuvpJYkaeroerEVNO1v+F5Aatc9pedMUwbjTi348E4+guhJJN
0gzCUVwXTOitsMvslb9aFUtrk5SaGurUGKAPaCMw9t8Zhe6i9Wbqis7isJTjLQovWk+VKF7KPDPU
1IDavM4xdcthmHZENRqkmeJr9tqzzeQanVH7wLTKufEZOyt6h+Yho6T78dxm5ySyF994PBB877ze
bXSVbcMmGpalZUXpuRIkfWM1rRDCfPpDDG3gO9MdIfrUt/WIGJD+33/JSZdTQ5Q4ccBo2eII08TB
Yu8Umw6xp3zVXGQNf1aSTJZqRuYOzU5GuCcbl+vQxoTunB80rULskZWcEGkZGaeeNfDLf0C6GnGP
CvuPzh9fyjcJXInBq3/Jren9sAlN+3LwMZM9sSrrBBRu2+DiWeAKMIEmj3e3piWBZLmt38htRBol
GC7AyEOc/dUnsjQJhG4ScDFOcw5jpt4FU+tB7h3+S3CYW+/nimzfdmNHl9YqUZQSJZkSw2/jcBU2
MYrS7OCIqNBwrLNz/m1O8GSXU3hN+AA89SxKhDbkUs3/4IoXZcqzEn7jYTxZbS6YtdJJdNgycPmn
noXWZJtw/MQOSbkG91kLs6ulYQm6Hj86M5l51v0qR1sluXUQ/RLWRNlNH6PtN0FP/hqmtHgAUHXw
5fH+hCDYuptXNdSGIwxHSwnrQw+eDbVvTj649Ce38Af0Vv0+NnOSU1+gDyCRGU4yep8v0T4uOTiM
WiOGqYg+B1z8Twb0EeSmQ5ahP7zW4QDa1mTBmSTIkLxA1Zxqls7pzzxoGVTlViTaTKkl/U9Yz7U/
kJtxhkcXhvhqEWUpZqdJ35WpMIeWJx2nf8lqAwvz5uwDc/SMCKnafAvPlfpPm9Juj5KwJ4GtfF7D
5v99/ZPnT+N2vMZ21snwEKNRRb6sUzZPVNM56n4Vga4p0axLgxW6U6siiHa8OWvdv5NUZpJjLc4h
TqJy7M8Z2AS7cSfivQ+bssN1prlc6xSpgRwel3996Cr4OfkjujP8Aqv4DGd9izjgGbxKsOzpJVE6
2X/hXeG8jyZFmfnPYfzLOR0LVH0vSqq0240uH96IPLtUOVj2iVIIiP8IOyz1GG80wp6MeyrSFkm/
EEs+209Huczw8UziWt+B0B67N4CjFO9ayKMb3Kn1SmFkBV9GZKxW2j11Pt5I8qekf1sJ9eFbmx5V
+cILk734U93UlRkKcwe+ZyYLiaKvk5dliEXeDBfhhH9FqCCQqT9Ow+IGJpa3S3I4kapQxutZ8Rul
zTvw5ysu5Wyhf9PKZDbrnT148rPHEG1Zh1Sa347RNTgl9lHFsT+S2TyHd9Z+7ATJlC4yGh9GAC0p
ISy8122iYfnEdux74IRJKBiR1vOatsowBQP2dGWwlU8iPSSTGk4EP7IF5ldNBKZxzJ7u6+GcNfGX
ntl5DDvf26GmBb1RM9gmsUeOc/Bv6oFmFYQZY2FJbMsBifszOh5pzXWYHKSmeP2CvPHmoA/aRGTO
O0Ml9PkcHiXzKqIbpjRiPNpwPCam8Ok8D2VV9DV/PdYuMQPWwThRsT5cH020hG0MNS++Q2UpnekY
E2gCUcSssiOdLd33sAZHv0HNdYhc7RdENqJJ9UgBPkSTgTRYKbaOVClKv+Z/a3jxjEZpXIkpUKyn
9W4ioO29AScjI4DPwt2sLUpvbx3+dEOMEuZpc4ziWONUQSF9II+KAEbXUgaSPGieVrT1FSYuehQ0
H7ezINO0qkIQmNWy5N1a7tMD5QtOuEOe5P91+7iV2gWUTA6y/J6tODC9SvTXC/x5rsgLQDkrybKq
KVSWHGXe56+SiBmIxzO0cVqlj4d/aU6Luab61/7dtOo1x0tw4QaluVzxlNVYOR94GbTCikztklZZ
6dji4oAhrWXgquE0GoqUsqFAmznBsf3ZIvqj2IJY9tkyjvKUWwroKIAwBMR/DlMti8+VZsu64nsJ
p3jw+BDLEdEmp8WG/mRrL4wnnP0qV5RAnqMyfcANXwiOdgaSbpbMW6r/7N/bJrLE0+xBIsDUnRFH
GxsUiVF4Esm2EgQOSK6myFRSLvlUgDhtHMe811yBLdPa9RMOmfiD65QauXdUvyfDhUYjuUkO5GA3
2NMkkaL4bnHimDrqB2AHqWvcsI1AWMwZI/8KHYQQwRuZccMheerRGWVgj3LPahya78jF8N99/r43
m8/try8wvsjWkK34FRDs1sGPXOvkggulTbCJ2rb39rxq+06ULyeuuaGLT28vkjFwaRWPiR0d3HUh
xH8uAAnf6TK20xBWGQ1L1UAp8J7EkUk1wLIWSRRxV/bsBfUnVfPJTzBbiUWQkyopTTg03XeMepiq
B/at3qya3q+EEaXXJqGQIB1tZvwdgkRCpXsuVbWiioTM2nIFK+ggBrkuw8LnOlubwz3Lk9hXPNlO
RngZpQs6yqjabnYAn+IHt+OFXg4rlNui2usE/+TnVMMD1d4952F3zpPMMF6iXS05/8FFan7ZGY5c
3W6TDmpZwrmxozu3+EAZEwU/+05r9K4zyHnSrSXiaCtoaLwxzRkyK4hcHlqF1aeaYUzsnsfOMRoY
hmVx0leo1foDoTLiHlQPv74UXUZ1xni5iCblBmdTf3GMzYZnjtnK3QAxne8fY83OhUxBl3iHrLrh
VNNRmX374RcbaEqgTfZDDzw1vtD7r2GljuDgI1vqcM0yGjaXDuqnNJaIStvwQYVIzFA6mJJfGsFf
YfCjrRiU6Fb+8gQfUmJoqTUpjqKlJOSVjRuQsRZxH+vlVkgMtUI6wQV+L7fpLSCcdqC8xjvTqnaO
jJK+D6nJ+WWnBG4ZrOxvBQrBjY04ZX/vF1QtXPpcIgqvhk2BKRcFj2lQSU698RsQCSTzgQ560bXx
tkhdyZr646gyG1t4lNJtUDpQr0BFLBCMgYhUM90Oj5iIJuQTxwkEOzrnmFVpafYhOVpIHkVD5SaM
Ucssk3OOwM9QBObAF/gDJgObYnOClak44ffWGUkvoVPyxxf6l3VtvNV9fMDMLVVphKIxC4KkXk9v
Gw4zukGmptn8xs6e8XgO+853YW4VOOJyqcjnIR/w0UShKuYZRx8J1qxLYiim7VLiNdoO4bBGBZuL
WUmQ5nsE3iQEuHge4bZikVq1D+9/LKJN8+Ke+YZXzbGSsbLb+WO2C65D8b5y+5+Wv8cGp0msW/af
CsXZIWRSUXIuQv+E86+9ua3PMRljIY3pfAlZjDzKaPlU/u75pPygtxlJ+PBDsm660N6v3ZwFFJ1Y
gsOip/WL0x3gIZYC1xYz+ZZIxHDWMMvsXe33EeyQvYFVLuHkdXN364Ihk5lUaW1aUHRKGxYM7tZv
xvlnWDt28wAfNwakVxL4REljQkbv8WuTkjON3Z8cqhpf4yf64UJgUPcMwvAMnFzhFlUbm7aSoEc6
AH1DqvLJn31n+Bsnl6GOo2/21QInmFW/V+vVoPnR5vBMH9s04pv4VX/9sGAGSuP4vkN0k2ge3Fyz
xtnUf+c0ji/UvLt9Q8aIjfho17h+iBkEIN2ie8eJEnpDJFigAYDrLOR/EIGbU8pGO/uHtZ7AbmQq
VDdHNBFz8bUfaUQZ3u7eZlf1Z2hgEi0COZw4sC/sO4UAcLX+LppsvktbVOT/cXvkuXHzKm3aOdqh
7YYuE8AStBkfHIrC3nJ9nLdCs8bVoADScQkp74yAgRxFYPOnewEr0F0WmMhb6VM1kAA+vTx17+jO
ApgkSSDWSEVdgNn0trmP9gagrJ/KpyNlGF4GUogR7+8Gd4uLCEabJNGZd92mFjOUFi7cPwgfekLK
+kfxifFNL0YH/aAKNo9TN/XBRiOcpGZzWIATCWayHGBlqnFAvFLe05buE94IDYzpxUzkIwWXCjDU
o++FOj2R09GvaPtU7DawfnnL24so2NHmZHd8/5yNykXWLSeEqepaF2kLm18NsHTbcYoRh+6pZhkB
Jo7Q45dgpjIhRcdhRmnLtE7DQL/h58RwDta1DTMs7SZ/MI0/lKgx3xyjA/lNqSNPQVB/ba47COrY
I7Djfg9LtfNzhm2tgw29Rn2JLhrJVXEQt2uj48sj7Qkfnbgdg2W9vO5elbQI0J0t9C6lLrO10Vsf
E9HrFSfDKhi6pMoF8x+bYdAoVV0qWg9Cgp1vlIas91yRU83xRebXuI0apX7eAhTRVzfqb2NE9K4H
VYgDlQivuYWov+uZGUl3qTAlWWgPnlbTWOpFCPq/yO7cQD485qpuZXq87np9m3zyCL5EGxInu4bc
uveEE90scJK1NEPfSlOMDOSb5k8p7Jr4EUhOX/Ie9BhTUeTkjIvoJHyrEdLRTgTd0mbdXKacSuNc
ShPJuHEVZ/dlaN3D6vRdKILdx/7Sai312JMus8d/IwXekdYhwHboWVvVBND1iFT5ceN1alCNBkvD
MACSsZNpeCmbnAfoXXYsiXFYWF4yfeOddN+x2paerRBPZn5ikZhOPftn4d1cDDRZANgv/5z9bvOs
6Xxfg5u2Ggs8gAHjGvokMtvFluwJCVoDqwG5Z2HpgDRJmW/ySAdPmC693qffHg0BF5w60Ka1DGCW
pQi81b2J9eeJDWwjzAzACzpxgUh9G6JYLY2TRO4CFtM8HJAVoQ05NIyrCghHuYIdUG6sloi1cJG/
mTXn+4PWGwWtJI3St0gJb9mHDwcefLQnpqvxafHTIj0IlZTe2GpnVd7PdhOCE/YgxDHMJf65PdpO
VWbgXGNmpol+lN+nZBCQTXDmUJq/JA2e+DukipZlQJJfCX7shaqkUqvzZ/lA143cL6Y7UfnAEXqS
L817CtMMtCOseioGhEghOLSVck7vXtbbX8Ia4JzVDXvRsOD0trCHiHILrcb73v0YhL8HWqV/Fgmm
j2HVHI72NstfpqYcYGUAHB6qZizHp9z/vP6WbPhc2XrsaA8FbQjsj4YO5FIZ8KL7443+IntxdvVU
ceqV9XWsK59NpnPzeDsML60F7D22Gr4CW3YeISB7/aTQXy3KvKGDNr4RasCNRTmntWHicf4k5lmk
hTCoqBcd4q+vtj1Tzt8L+Fd5WSNvRMmOaYCYi6WxOj/m/PlZ7ujlhsCxn8+R+EIJsInkchyTHTtD
FikdyxL8VgA78quHSzZssbdjfy7DRDM5a0R6sKrMlZALgCansBbLTSYBliGEZTvVe4RgMsdinc0X
oxyGQgvN3ZVZX79/RFbe823l9OfebixfVXipeqn8dKSdvr8BkkZYFAlEVHjrSofk/rwxAe9fZ01h
nNheEg3so00eFfmzbc4CQ/Tv+AyIZ3+VK9a/KJ/dRLXekLGKKv7KPf/MZ+1pbl6rEkI5L3JpZF6n
4+MMLlI8RSwmExn4kWCG/I8Bg7AsDq5IBGLfcMsAa0RwK9bW1mryTA7X4kAZKNZbRffEDoYC8c/A
pDegMrlGJdQAtugZIXB1YpmkxgGj3wVjQbGglwVI2P74gYItueF1nLNRwK382Evd15mR5HDETcKb
mSUAfoL5zrlC6e49rS5E+FcoidAiKuTKjnJb5WkaWQAapRqs0aHFhk8+8VesUo/Ti4t8FpbTWbSz
lvw6i+/kb0nlTxBQKvkvVioGQSjjJ+pDkyHTP2tZmk4opM+Tso5aDg/uFIATHZXXau5WbYSBsmRZ
J4IMEjMry8ePvzD/A8TPIaTZ77RALzKlSzLcw5+iZTGjdMHCzfKx0bsUDEEsxn81TtXTKali8NwR
C4+tnitbgYeb3fQ74hhM32xu8qC8nAx9gQ+t0C1Ceuv8/GjIMs8PBbNkRFHOKDxS0feXirStLkWW
xiIeDJ+EIor/bnU7YKnnNX3yTnhPaB/pAmWvbMKIdul3BlpgFiV+RvfADlViQb/2AEPG6Z2+3ivP
7g4Yua+fXzk6NQ0P6FRlpNLqsVClbeAL7A60hVLURxRONdNvDcdFPi7u9rAf+Y/zBQ486lkWaOeh
FQc+Mh7o1t2ed1PTpTIeO/1ffdo0D7se5XPNY4nUnrCPE/aN2uNG1tAOLwkQ8UftjfQZjQH2GFge
WJ9FQXmUAnoxPagkLqLLs3WbqZXoEETcB/E7FoP36ZVjxdJNznCQYoqqRoh4ZrNV/En6sJwLF4ZJ
cupquqUeYgKH3C3CAOy+I/IBq5Obn55sSSSvY6shA2r7r6+lQqh1yrH0CFHecqZzLGBrkNIp9WsC
Py2vo2mhVY556AdpRJ+kIC2USemkvR5tMmu2vjwFZm1XOKKsCnoiRvzuja8B1Wxw0MlQaiH+PQVU
XTfdXbjGTkT/pc1TUV7zcA4rFKkp/h5XwW8+TqXodX1WhelQ9hxH8Mc1Hy9hezjjOut3X/UGBrWm
5jZQbbLMLiosd0SCPLdvq0ackhX4Xmr6/LdhHhexrq5Mj2ZzL1B3RJL1doolhccN73FpAT338leo
ZY8gDzh/FGc6MQMDT/CzBwtuFqorec4G28Wrtf+omhCUC+10SyG41nL++gMS+EhByZkezOLyIniJ
QFtw/uVxySce5VwPKYFU/WcmdR3YarMKvViyAYVxEUyXNkkHq1RynAON7SEAa01GbjfnCWQjj74B
eKcL6HlL+i1O3x/G6Udc8KdL/LLN8FdkU6wthTlqiK4lpsfl40WjrSZxrUtWr/T+5QrKvH75L8sG
706nHwzZ84U4FbSiBxEcKizqGJoDiH+aLFPVyfS5skUdjXX22pBjPCuUssIM0Xj4MJFtEEJjV5By
bqkFFRW4xmWSVF/M1IHpTJ2rLvTt7MO5gmrtSqQZxNLNNyUsp+qo9RGjKYB3DzPxEIM9fJdBP+66
Vkaw9OIdYj9tGl6Dq4p1xmy4F3ZR8vclKeDsy66zY+s0OEiESeWuthz7X/V6bmuHLK39Bd4AhizT
E9WzuKBTHvbxzcUt6rtAD957l8OIjz8tRq6+C0CxkZkq8KCA/Fr3nLAiulrGAtXjkIZSdawlLgSi
APh4Q4fReDAQhkoCPRrHnvC9cl1FaLWK9qgYbSrYwdv1vWbwE/3cDFIyVSW0d4H+aIRyQpaNFxAR
sKts3jegtAJuC41VdgKdHm5xLIuhZMJt/7FRvQwyz8VgFCMfrDC62Nnad0YY/QeIdGIuZYm9DUOf
Iv7nEVEIu57C1J+eZxAE4/evw8Bkxzqp+Hpam25lKF9qYwnfLJGu5ZhdnIFTfUxEskK0y4JEbF1q
qmfBTHAAhck+aM9zh2O/qXJGsmomrcnh27SkgZbJEWiK/42zmJ1zOD0m90Tf6ku6aFsCMaiIXjV8
3hRnYe83Yra3o1eBUBliOHHRnmJwNwMOpyvGYD1wn1L32CRPwixbW0kVCceqEgwyVcwgjnlf9X7W
ZHqc1Zcxy6FfpJqfEmub/3XjtxtyqqSH8ixpSRmgWVvWb8V7A8FgpTMaIWkjRGfzpMZiCvdsGQUc
+peuAesE7T8U4ja4TfudB8iSEhKpo51HN1asBd1n8u3k+DifKDYq8kk7NAyh+1QyEZsUpETe1BJR
dBYbuCiVt+GKGKYtvFxs54Fze5dRO8rA8OuBfpR3KEYuaWHjmYjqqYyMyha2Hj/XcrwQx6tapUDd
7o543Op6vMhwFeWkA1RP+SADspQOeOYWzRKbmmWQbg9NGqM7KG6/7+NlEDcHPcdzaQpyJaQHeOe4
F6MBSZvTxaJwcqelPRv2cey5enxSH7iwnwosTCdIe3ipBozrqni/npKtYujyYWFn6fHV/NNOWnmQ
pVckeoy8lgh1ujomS2mavv0h2OPNn7vf02i5h2nwOK2i7Xfv40gkonU+k2oIrDXjf5tT1Aq+SJQZ
mepqQy5q8KTknnrpLFLT5VTN3NvfRXkOb759ARxldw3gyqzoSN0UsWll3VLNKT2WLURgYNjeYwbJ
sRMxwc135NUfbtl3uunWyG/eUzD1OVOxjHq2J+OBJvt1oE5QsXT4w0VqPwV6qTarSSBdePAfUAI3
jcuoTfg0vGii5DiRI7c6xZa3Hl509HbgHOFzstgqzAwg3eUy9fNhvIeHIPacOdyGiCUWhej9u4wp
mTFMiRzTP2CvX1Js7Uof3M6vbHWRfofLZ1u2iG0guU8reKYZOBJZTzGDtyC3stDVyoTgUGJ++2n+
ioFk46V7ghkTYyzcTskl1WB1ipRN0bCUyquqwQczuw6ce/izGaKRxlW9iP80fMU724N7RN91xCUs
oGkB6kslsPN9EutrVX8Jne00dgRq0/IZ0LJsQE0/qlBTqn9iq98vomr+nukUulLa+cosh7n3JaA3
LCgwZm7LSVpPLSYuIe+eWQTfhvDfdppqeM6WI5zFYcht9dnOeOny1pROWGGO3tBFQv9JMOTlU1Cm
bQ5QKjP2EXcgStt/SI2udzuzIHCSos/aJFcHWmOEqKpFwQlgpM5BvULntVdVqaG7PyUbbvb9zvLG
fq5iWVkuh8iOF00N4FB+siZ1bwdOMDF9NoiMFKQ3wujsDNo7472jUVykrbaFzMOHnZKcXTrYkmpu
wvxwfj6Dy++1PyiMEvp2VN09OhEEdJYA6n69syswve108cchll9uM5Cmi/5/W10e+ulRddfTOmEp
sl/liYH5QxYJFY8fOBZnVRL7zUi0DO2j5V9xUIQgz0b8Q9aJGhJS9HsTW3ulwjvpwyS6FHCoKUNw
A68KBS4mYLqnoTDU86fOT+d/51xeuOcR7V8c7Iq75svGAO4tAFVDbiU8Us/dsrwKMd23zWMKZzvh
FPkKYCSfeHfWjgCpGlCzVERnrE+j26wc4w6/hIDmrZsScQmVfiWD/2ZJ5TFp73VHVcSKgIX4x2Jg
syoFbyCcYMR8xGiFesWb2MUEQnTb8viUZS4UVxM7N9n3KATa/GU2/rLob1iEhOp/ZIfSLJbHS31W
yJs7YGowIz6mIiZir5GmuN8u6CL1qWqeZ4ADIKvdokPRv9kRgQ421RzYYTvd1Eg9z5SvwFUYn+sK
1Knv/CMtrT3slFSeICv3+Dtrw3dh37WVQbZd4v3afGPXCctgg9lq961+yKf+hvjws6nSHVkAdXeV
aSKADmqWP3hky7sXAvPtRwFGdG3Vxhdv4Sp7AKFpkXhCFGc9wzp2RnWH7F4CquMONeQZKs+BBRQa
QIjsyvbtpoXr1LPHR3OBvoVqQsMmQlJRv+LXrzJvOgmBw9rYnuDU0W80amydZMhUmHaSd9f0L47X
NwcvpgWkxOm416ODTlroFIHZaGURAR9cZtnw9HHp+Lf38d3MgmI23g0tFgXUuwaTsMfTR6BjeUd7
uyXs1l4ORbn+5sU2GygDNSP/4TtgcjtZDrTKNShRv0K76Jf4k8qzWRvBIXucmbxlDDN4nTwZ6cRj
ecrJxqvku7IN8zns/KGxcyqlYyK+6C0d1w+iwhCkdLRI5LgkDe7Xh+sXM/pbEa3GuzgcOVoRy0JV
bVkI5Fx9o1DmayH1czI0h7tSqIL4Ba8HFd9n3o799NyJzvjkr9/eI/nKGfc5OxAVq5NieAE0PVYk
o+Y/lgrQzpWNK6sGiUQKQNeWZBo+C+YqAezxGDR2MgjWkDXONGn0zACDoTxApfqM+Krjo1dkstVQ
1IFx+3bGv+MmrMKahY5YS3b9cM7qOSGZrLfySCIoClbg5kpE5Pnu5nZnhFtL9J+P2n4DhBzroc+0
1Pd4ZLBMpcE80mPJcwW/o3h020z77Zom6v2qaCf5E2L4hXhjjbNoal+/oL8YWnZ4Pd29BsNuiV4M
Y2an+yVB1pevCkiC3Jc+2qkBlM76zn5CC6hdqk0z3pQKSkAcCQOYl01pvu2vjtHAyLL3RC3mxer1
goorSHU1DQO8GSBYZE0/oyoDWEStmpQ94UHVB+GK8DFh0zomrRKDhkFSNj8hGEW1mrcquNKZIni9
Krvq7SFy4xA/JYtC/h67rc4MHG+FmoIJLPAlJEabpkNVRIbHgB1hKQP13RZHxcTPyGSc9+rm+spa
FEflz76EhzJG25/JYHyfgZIFX1l/QI+B7ZK+EgmS7svobJtHrzNXWJcNEgB+72fRsaQc0LwBLisg
1AWLGLHT9UCY24tYNgmwJq5ySqNZE4hASHP/DT3YAS8kBsGNy/BYoKTERCWKsG6MRYjG6IvERbwj
kOwRGVefn7Nou6f9E9tYujz5kD8YDmxF2yvEtFv09SD5eQk1ziJINWks8JYyX7VsCUAsISucrjBX
5AmjNPww9gVTK0GUg0ujecbPAMPiGJQ89LMs/FuY/O9GUGNA/pT1VB0upffaaOkePl4yTiEhv5Y/
R0lkiUM4hFaSfRsQQwvej59yXa5y3+ZXCcwBM3mB4vTzTFcjs8LrIAq7SRzX/kNjCNRmsDJzMp5K
HhXXEcen2yvboqeONtNDR7KNgfl053vjXarGKRNvIgCJWoz7QXOQBr9s0we9/mOZ7buOYS3Rl5of
qvSvF8JPoyQkx3PW2YzVIxOS7Z/wx9x1tXmAghBdWPqsYRqhKWrZImmQhX/XbuwEAkX32GkTCW3S
oaJquGdOGY8sNssh9i0DDjraoqW1YNL1r7q35eLL8a8/UCUtS/Ff+5K2yJ89TnEOstTy382FlCiD
4IwG1P5vzNW36Q/JeXZoWGI72afd/Y6o6TLgGCK19WGMKVzfbMqkW8D8sy17Yuyozh9YoUuknWHl
oRIqSwX+bXDTCs8eClSVJGWHrWGuccD3DlThtQW7mbpa1/1BK6e5u4+6ZlO6Am7UQBpEEDukGZ5b
CX3+xqeB1pMLXcbWpEK3E/jTaN4b6eobvr8Ko11b78wnisabzuh7aDCZNqDf8iRbIB/hbOvIW6t7
u5q/OmS6NwhDE79XhSQcPYxGBP4dL53LgDaa0InICljYSxIpsApjnPITjbmonGkmhE/7TWc/1/Df
97bkGGoYHzMO580UGI/6zbVxV5m7nTcVr0kEGAxc81cGwEZcK6AWeQfZiNFKWaVp1yyhxuzZHnp9
OAhHGgnBxmgTWipwIE54z7f+ZevZxE1/brKcGFpmVbEqi1ZfKUFQrnriOn1H2y5Wk/M6SFMaV7Nn
+x+ZxRiObDLsIZ5fmEnN53DTBP2fbRWLlTO2a+aly3cMS79CaglKm8oHEyjNFkhuf3c7XjkmrEdb
nKBpypoL1OdUXQIal8+BUjIr/TUoWbFe6U/4FQoPUrowJRzxJZ77HWT2htknyei4seEvxImiK1Qz
bMSxg+etvYXBUqIfUHuCYN4nWcIx8pr0ZO70WxV1tud1LPojzulyJ86zPcyn5zJ+sXSLZId4bi0i
RWkFhd4aYCbioMDcVQ8cW2vxXXp0r2kkZKXXm5N18SmIR4wnMEfgJqCm76OYpH2HSRHAjq30Jzk4
y5dyGAp54RPK7qcsSEM0Xj4V4di/eUyiTtw7UVhhpeZFJpnANVVdq6PH8+teQYPFJgq1Cp9c46TI
YuAgX1172Nsyg8rcjdoji+x9nnwKd+TGrzN87CHIvWgH1bmYHQWoy8NC1rDlm/3WfSPfEU3sLEnT
M0Oxtv0bnR6PLs/8AdNUwGybogLBlX2bXvOSrQlwGDos4iLvygstU1ADxOAV0J7bZJU8sKBvuGxx
4LY3GfZ5d+uRIdMEW8iP6rajIenExB3nmc6p+Gk3LZ8esV7L7gBdQq9rFD8EZYSDOgr50iSHDSv7
YYGd1INpeE0WHCdEHSdg6Mkj7NTTJ2l1zvnDQAEWF+Wzvw5itZif/7MZ5RQa2+TTcAZ4FkTx8wvM
y0PQ5y49YC5d+y9UJRMgqpvMyNcR9pRaqLwQRA+5kU6LijJOKtXWAUsIiFdcA+rb4Zb2M3fNwIBn
kifdO9JroA2aGt1W/6Bj8srCldcp7pg5+4oEqZELNgLeFWPlUcELCh2Ph1OwmwQGbV/7LAb3avh2
0DGsM8Ssk3EXSNnGFPJm7mXzM8DBAn111k1nHqCiv7VNIjEUVfmFjfJwp4q8RP/ZWGzbbeMDAeXK
VXPrheYmwrXooFdfG89KPiXCnCBpRTpQNCAs6JLBA2Ve7tO/SsLrxcG6vYJtvpXo06h4HAO10B3y
Mhzv/g73ZjZtsk8PCUxuM9JVfkXZpOajG5bKpclPcQWEfILacK6Ffcjq3vUGHtK0jbO/HyUmHpcA
T+DssjsnPZnui9GlqT7n3k2DKxibibygTHFS7kW27yG2biDtr2dtsVjP9jaj9pCiHABVLcEJ2Rru
Cy0Q50IdKtp0wm/w+mDNa6hqA6Q8UhTHlLpBLzi80syiAGEso63O7w0/uDCb1ejjXGiUGOzisZOz
yUdQ3lShfIhoyseNzcumvOvsgkEMFCDdmnaMeN+Iiz68R4PtSDwI5eGcdrhj1J9ZnDBA+7mBFk8L
Atjivics454GIP30tOvBpL2jWEMEYCP2d8ojBzgHX4MtzebG+DOTSKBZzY2gPUREH6dvP1D9/1pL
NylW37iKMrchBRsfLbuztgk8NfPhmSHy+0/VJ4GUXi3zuFcd70fvhqb+2euRlV/ByxntvloWwzSr
oyD1Gmjg3QlvaClXxfhEITBXKzScOgP47lVhkcmM1ZKE1/mkhyRN7n983akhm0qlb2pt7wfr/jXh
GSj1eipOZ1dDTRqdY3VcKCK+Als4Jy/iQkGZv2c2xl/FG49squ1PgUgJAuwUbTTSanJkjbcjHtFe
bHHPtrjn/PLbuU5LifVA6XOJRMUEMKpD/+s8MdsEyUSabznSux4I0whzk4OLalK51vkXv66/rNcH
XNiivZ43wF8qP9jFDHFSwtTPV7wXop3JUXTfjh1PSrqFvITcy5c4uZHIucQrklUCG1RJxdGhYFtf
OLa/Pv/Tb2Uv9rd2TWFQQHf1JsiDCcDlkLqcL8Zn8DKtoebwNzD0FInJrOUSDYXJxpdOxwpPybdN
5xeNKynnW1gksdliXWXADW3wvMNvggmHIcGGjH6AzT6lZV+sZiCOFc/ZBwAOp8iYaXa6SNsON//h
zU3tmbiB8rmyl7R/Taaul4+9jsYC6VesD/c6uNmqPNdf7LbBS0plhLWgYFQHfj8Z1v+JEAf0RBRD
KSX9Jy38ioN6lBFDdX4mxoa9BG2r2jPFdqFm9pgBZCmNdQsSrEl3fqdIm7rUEvUckd/JuVSBUKqH
8RMTPb0YouVBAm+njsX4Ogsh32oVlftKqn+NjsyNVrB2mqtk1s7RCunqF0PO47u3DmClBHA/8Itq
MOMuJc4szkYysi2xsKo2jb3fOYEn8lo7l1iqufu3tTP5Y7E89bmPYnyAiE+2Bb1o7hVP2ZWE7r1x
AHMkOcq1S4l7M51QhSkWYs5zN16UNxvSfCdXzG9MpIgl8Ov9QAezKNZ0aBkgLswy7URRLwR+tlzd
edwwVPdW6OhSM2BiVVktjKlc3+mC0ZQYDvKfdnHRPGGnhnd3VK8LbCK7UmtNGj8v6t99BgaTHFQu
3DTH276ezlVh/6OLWq+/IC/JGG0oUQnhLYlcOcirv634HUMlXUR0q5Go+ev03tk+LBs5NCMRDAxF
g6HVOK91KtljbBFugEoMCR7pltuCPnP+EcEn7YrFnMP+Uf6j3IqiotfxMBKFSYP3bZYXWFvNFRk3
HWXAGlSi5h6S0VAopZL439XgKUqEPs4HrhNaaMVWu1vfzgJRjgeMhIVNHBZPqphvN+hcLpWSMoJV
+1U+hI948SJrUNIuy/aIkGYBdBoSe4fPBIxFhmpn/OpW3CHlCNYfNHSIlBzOdb7ytwbI0Oga6zls
5qYgLWQupkuBEzmrEJdf6roaPlN9Jr8IM50f4dfJyCU+8LBy3rQP6dgCaU1OxT5M4PflMlhAXufg
M1dKhHDuOVWyyP+LimkJQQ0lMcSSEokCmsUdC+xNLLiwYIPDqyRE/NgSM5qoI02yebZL62uTKZPA
gjoYnH1KHE5c25VIVlyt5AvbglLRlReG+0gKxwHJBjV41kjliTunGSNz3o3tw+EpKEHEq27x3nVL
DnzgJql7CaO3s5C6onezR9Am4gUbDpDl+57ApNMULDGWAYmM9X2IVOykmv8rdDTxyVdM6R9umWW/
hykO5/RhbErUPipg8GgU7hF2uEZqMz8aT6Vd7Q3cudhqQHM+7NLXPWXG9KRWk3LWjI9waUGNA8Td
W/Te1IauI0Gg+tlhJnTuoh3AKqHsSNac29LP3s1EHiWLo/LmVdhT8AXstH5mfHiVHgc/GxV6KztD
dtheOF/LOgTv2YNHiXOr1aQUoUxlShkqdbc/LkAJru/9TuxolAYWfCiF7ukKyz0+g3YY/n6zIBxh
uxBkAorP6CDGSlclW3Q9uLUoyJpQ+8t1iyshDOUsc1l2v3Ci9TW7YDvF9REf2t8sjnzND9HxM2EG
rSZ+SyJKwiluVrSQUvfUlF7KgmfAPzI822fd4QV9HJB2DnLjYOF3imFVpoi+uDCX5it6EGNi4w/3
hL4qMd0hC8OJTNZygDvgbWf3bk7yMryvt8rTKNXwPoMsqJrxAgA9li57iCjXPoViW6OQcJ/pn0mr
ObElxs8pGu7cgTdOVmMdBgfSIBinqF4hQru7yeR029h4Gl9rXcQg1YR5tft0sDvWKJDLOWAlCaSi
87DCSToI9u1wYdiZMqNAw4r56cPMLOSu+uYn1bgnq93LmejUllvqSNkRhpfVOLN4KpRcEbRK2tS/
VWQCvJMUeF+F3JYt5FwtehxSKzwMaknrjSlTEXb462COx1MIk2r9VkcQrW0kWAW+A+l2DFV9M+8f
vwap6FR6POXTACFbJNnwpARhpMsq+KmFRO3ypmaUh3ZZRc18Ld5MBIzyG1Qosx9Q8ECL3vA/BUu+
N1QWsuRGkQkI5Rx6VWNcBX15M3jCttCFagebIZqW/NovV+eu1bx4ohBf6qFA1O8vO4CY5016Zo+x
dn4NLxZL5dP8ErQD837LRNGqoMa3Gfgk0/ppHs9BVGF27A3rkWc6+2nqXBBQ2TpAY52Hm8POgdar
bz/xoPluX8YObfHlpiPfqmDxDPZv3EMkkuquXGCjqb6oyqPjq4V/yQwkcCXLGrD3YTug65bJoJXW
Lam0uz0f6iQpZFIhfowIziitdoQDj2kvqxU/Z0orZ1IJNkSu1gq8UmGvyFpeqyRISbBLRaz+2csE
EUlHNvraIMWW+Dux9Q45AlYaNY/v6WdNtj05e8u3pKeQ95Cgyp3FHTn3Hm/Ule6A+YB7XZQSiQmL
jiusMulWrHxwaQuki1e+MoG81D/eYc5V5gXRd5hgY8Ay+lXseuhTk3iB7YIGkyWE7DAgkMdSCWvt
Fi93GO22PgvAAhOMb7LM1mnwzXIqtlq6gcOlFGlPjMG0zH/ALwrmFqyETtjeZE37gDo+pcIsbjfk
fLs6l9sYi2GfgA3pJVPLHUFv/uKTVaB9JAcHXHkEPO/sDp4GE+Hnxsh1XikCiCXnYCw6G+rmV0kc
LC0eoG1EEZ5NVKlIDgXKZAUZdeNYQs8BfOc4hFmDtelmGgpduhOKBNF47I4wmhZ69dWU7D+pwW++
cy4tDoWzcEAyanuy7FMAf1r4FJmARdEb0ZA9eMsvkP9iX+rj/3UBcB/RZaQhAQsw0g6QUeI8gC2p
mbaSvKdKPBGbbnWlbDAKLEK/hadCwnUjViieJC7y7x1POpwVQKGWMPl3zRBZ4JuY0FBrcdfSn1PZ
7GXTcdnjlX8LkUI3bmbFag8BI6+Y0Q==
`protect end_protected
