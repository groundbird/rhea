`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GmVL5Sl5gxFpdB9Lj7KiiQs7sVvYp5JHeq2kQKbnQluhfdt8SIxbtqM3cMLEvUxiFjYBCPS2T66P
XDshh+DUng==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C0kONuOU+Hm6HdZ8IZLQ3HPlu+EpLCFOD4o6Eq7QbK4PERBZwUVS8Zwt2O4ORrdZ2nBA2KWC+9Ul
LMqAXPsRGXmnKsoYy8uRK6ifc+e4Qtanf5WWKrNKJdpMbKFNYHNG83YDfpSPVGkYLqe6M49aKFzV
vd9oLvJCw1bMkfxIdOE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ElEZxFNRqufO873T623/AiSRqGlRND6cKuuQ4q0SW8uFwmJMx8uAq5I3U24hspmmfYHAu7F61RJN
2ovr0swIoysQjSIX4M6HabuyUJoGNsaPD0BbO6gK1UDWXCDLi4JleCzHFPWT4pmwPLh6OFesfbPt
+0k3EWUdQrEKLBQn8q+Ydf538KqIJDA0x2iqvgtK1ELmQAvE6UXuXgSPHUhBtyyF8SBqsiPoseNl
IMW47u6ykVRVBE9iwlh+UCtpDbM1FPG/6sl9S6oqw96AqPiURaEF3u9E5q+0+vmYqVNEEfPLHs7e
gz8yjmSh47OS4YtHHy5dfleQ6KDRIckhry0oAg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P+5/IWiZIjLHpIQ7IOxh5G53wIdfJHldUuZtbc7L32yf+zQHa6Z9UTVD0DfCFaWKFQItQnaUDn9I
+nT4CcWu+LkF5R6B9QMw7EpACOPpRZx/3HlT+q0fX+fScNxuvu01pDfrieflOPQkzckw6eeDUrdq
/3mdGxZ6uOae74lUxHs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mZx9yTmc0odU4Z1GutLHA92gsWbuEtiSo58aioobVs/5+efy8QUXExNFrLoCL1V9TNBcOiyZhijX
UM+Dgv2Q8/GHa1kmT2f8vnXHuER5esRPSQcYPnBWB4HT4POjtc0ERVQuxiGY6s0ZLFJHkRhDDV+C
CPyoDBka7680qtny5flwsz4D0dBgwhr1xiBoectSB9xjEFwYknn4UEvmuGacKwEDtQyYpLMS31Q4
jKhLMNKUJBNqn/xjfCYyM4sb83Dve7VSpRGn3fDka4zc/SUN34QNlBp81lrsRShbvAQRy16JOHSo
VLKwlhB0va+1zeOvmuuF2Z6BIPHvZyFD1ejNYg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9216)
`protect data_block
KsVYqvdCdpxYmqfzYVpo2YNIslk3GHC8DOPqRdQ14LDPemfGXmSjaHlvT6C/vc5fiPnWn27In2AU
bipYZhAMdT1LpvgjtbfgRVmQM5ehNSa5AsQaLUPPJV7CodGazcDVcRHA3F92PDxfeQLbmiC2ObKN
caFN/bZ0X9NVw+pQaL4bVSvVUHMje0K6ooKNjXen9L2CV+7XZkpXL1jXWMFDgHORpsRziRgvv8j4
72Y1pIMmbO2MsPEm7EzG8tOZ3hvlc1gLcj23eNIxYB4PrpW0L4Ei+tSmIzn8NHzLe+Z6+6waSpYS
q2EUNtFLBITCX/R1teDOeKIVgihTF/AdhOWeEw1JvbOSIJ+gTVqk0j0sOTY7QswEHc0657gZS06c
B1ZJ/p6S+86FTHMYfCJRzFLiWSxTsYdIbSXeSuj6S8Q5YioN1wsv78J0Fnp8RRVkB0Jta//2dsBN
t6UKVYBF0Tj8kyxpbX8pEJBQvCtTaDZ35N9srn516ComdvWeokK9wsOVYxMYZH5yMtf7ybnIwo6W
sGVOO9bPDn1Au6rFaSamQpGSvLLdoNevQriaNWLfR1UkUjpMcMe6HbvJOZPTCgN8rsVRsqFeAYRh
UC1Aze7PY5z9pr27sKNYGCZoQS/GLk/QsnziYo8s32Si2gORhVe0+eMz/ysyTPFcPESa7a32THuM
RBFyJ1SYc971Im/Hb7lcXh07Vfl8zz5Vjtzc4f6PDrItr+6kbI3mW3KrSFV9w0rWjfwqjZzHQaJ5
Kb/ArOX3bwBkB/pkb5tPIZD7bpKQptHd5cerBdTNcvrpPYgZtmbTmORQ2RDIsfdBhfudBEZk9OIA
M+TjVe+8IZmidCs8d8yNs8UjjcOzlEw2JU6Pygbk59iV/Aza6Da+Di1993VvBhlP4IAUCrjuY8Ot
VPZgddHWljZN4hRE/DS/dRw1UGZaUejo9AcVNfwgenf6q7BrZn1rsi5uuJdhbXgQV2d49By6JQLt
tWa+YyLtBu/NrtJoMyAxeVFWOwCxPMfk7kV8frTGwN5u7cNEdORo9zRNruaQ8hpSJ7yXRm/jurWu
zClEq9g2R+DPFoXls5ZxU0m4wIPmsmcovPBzB4FaxC1EaT5fIM723HHw3u7Eg8VDbrZeUPuIs5fa
AYviMjKPmHw7AYDTVHkVHB6kMi9mci+kRJbHzLlVoYbJNrI3IhkVsDvIcWKMMQlys+H64SOt9Mf0
XllQEdWhWROLGHNyCjkf26JB0ufwASkouBYriJQEP1Fn1Cqk/aXSzvEL3fogJPqZMbZVrhvU5+2z
mvMiTxANAZyL3Dbzya/23T8tXWumO2cRgt0lp8Qs+0X+/vRKyGUxy15puhle1tseS0rjJpXdfBVC
k5vbFnpmsXfz4+9LUEKMXH0aGL6z4AsHGwbtkDsJPBMWXLD/B9HJJSD5TOQ2Dh1Pf5Ldkhtsc5Qf
09ZdIxkKj8bbHGyfA3o2cuaz6ok366fLnebge20QhbjrXNtrk4luTMwOHCEg/ZdhL7SY1jh+By/L
mPXlq5dWrvlwseRUQM51grxK/BF/U0QrUPoPDvdWxt5O1XWtKLfjd5sSA1Oy91GI55486Z0TvpxL
0o6M6LJwE3Vbg1usHxkNw73U4OhH7gyAyDnN+yasuSklDYJqTuD/yjZr/fuq6VcOb2r6IOpeztHp
G8NKMTNY+qJn5g+LWIagrUT1qkLJfip35xKfkhYVPLI/jB0YLzsHA17lIpxI7Glq/nBD9kZsdtzK
2u8c5sag5zKbBYV4XB0KbKgw9HYkjcEJlv/U7sqqIjngKyhmSse9tvgb1R6j5ZdL+7CJ+dE2quiC
tRowDE05LmvaZZevU12tQXDZlC7P71A4kkgD4gvjoq+VH2x9CFHUPNcxBqgL3wghgDYVJxOtZn5P
9ed/U5lp2mnSFFJK4zggRYTkgRwEorTUNAGq285K4CmWanS/lZURmODCUojS0I6jn/tgpf9qwsPV
kECHhxsUpMsa5f5j66/wlj3gk2XwY0aYtXrtgOR7EOvmFX90zkFOsO9jc55+sP8K2qR79h5Ylkdb
Vr9d4CqL30u/wfFX6WuyXGBNiKn3etT8BD6DA7fOqr0afLmmKOIRhnD27jiVzUF15G2NYqHclyvJ
j+7clawGOnipm+26HYMM38uAz/mvSCqnnT6re7zlJYUpkVyq7p7RgRqa+Sj8lq+CEh+pwH1L2MSA
coYxcFlmBi7wfo0J01RbBHvHSX4Ga76HKQA0bp2prFwATyazTqEuBW+bP5ESxvE0HzyQHwO+1fdB
aKF1f2Vux6EDvLRbCzKY7WkUGKf5V+IzI/v2V8ffvA30EPTSz2C4s3m8h5Ui8LPoqPPZzBneCpI0
um/z4rB/pQN0nuX4nsy3zxjx6hrBb8UxK6jxidb/jhzGSkpAFJhQ9bQJJSNjWJ41mPlsm5GjNVmz
6OoKcD4OxaK6Uk7bv6JtYVwbkkRLrB0Y8COgpWhHVvBJmsIgLJmawd3HvOABgy0Q2CG5rZHyLkRo
MhJEvcJ3ThS4dBreeA31W0rniPR/TdNE4gYPRKqM60ivRpnzUXqacbWJSyqavZjKdlkfcO4FDD4c
bhSZN9dJx+23iAKCcO/PHYGpeDhjoqoaBb1FLyrdvZa4+Wg+W85qTwXInJ2XY6TVBKcxN0IcG2Ap
azR5heHBf4E3uVYooFP0QO5OIxq7hU6CKfXGGzKyMz+Y6DPAgifzhyqXpYgJECJtdNIdfJy3TZVP
DK5h2Vl10T+xFhj9dNpb0HOn++iXGVl5/FD83LzQjIUdKHbeo39LN50s8sn7I2xebgXW7M3h2X+R
BBCiIKsIIV6Bh6kcpfdIkmipkqtvMgUx9CkpYtwmmafUaHPir8mp8mEI5WKJHHG+yrLTHXLDte7C
NVcleNbIK49UDDH7XIWmDcV12Jdf4z345bXYuKyOgkPBZ24hMxKA4o0AltpabeS3hYBcWwAvEfhQ
tgIWaVeH3sVQBkaI374hhUt0iZT8rX3OC1tM/1d4qtmXldc/r1UbDnv+8ht55fM+7qe/DIPbuGPQ
eHbGBElNAtIVlon5aQsJjK6IVRJrspx5MIYW5QslR2kxb45KFY6aV6iosVE3CsiQu8oqfrCbvjsI
xlmBgKBDrrk/e6Dr74QCC141eYUY3MGmZc/u5yeJfgN4VpAfmGzQimrUzB+HEX0SklZFp98I8AEo
OgA2mMfLG275VagvuaCoNvd34IAcHWEekEzBNNG1QZYD+A259+Nc9umIe20L+odpyyZoQXU9PbLL
SNkiLQgJjqbwYam6qPPwuTscqttC1uVQN6ryheZlY4NBHjLG0d3pGiYoZJDpclSLIfz/uQypgiyr
oA6l/4i31CWX5mwktTzGZaB4mk5nQGvBRFZaEoX79Mj7CmGBQeQQD0IwvJeKeYzZTyXIedAcSovJ
3hI6Wg+/PYj4fQ23qlL/wfidVPt982exCVsSoxbRYY3KK9xZNyu23EP0WJot8/1idp8TfqV+SvJF
15jowiZHf6WRw74w/dg7fyTHkuXtz665ixvvOihuOjbafXi+mDsbzG+dykLKkoTahihFrPllfexJ
17Iw2D52fD35QmPLRMAnRtUvKSHMoYZSsjjsqb8Pc0+kK3FLJdW3audVJx2m0XJm4eS1NomIYGBs
qBZ5M4Sqn47Y0l6gaZHObGmH7TE8Iiu6++0fqnVRCrpAnz6vFXXm5JJQVP7hPHzq8f6cIAhIFsf4
kBpxtM1ja/X7qmHcvrJuzuoVVkCaTq81ptsoDZGuATu/ix0plLDCbbVnSKV8Gq6ENnKXoTMKK/XG
TW85tfNzA2hqhLm5GFwdXHI9DJdhcIDXu1cgqKYoI9kQkeklQ9YYZYZenN2N8O8uIWSqAUY7gscI
jHf4CkIDAq5egU1Vsw+shNAheHeWUlx0Ws+To9CVxuv0od7xy5XitJaESEJL4bukRlrfEv448Dr8
iG9srqocKkPHQys5hCxxccAJT3yLDFSd3hpwlqzbNr/4z1GyO1dlCiR6xeJGmnG7FrWUOwPnxtzz
vHBMsobUk2TlQmwjTckSrmHDSUkH367sheVOxxKGTIo910GA6YsQa8Uoy7WLGEiuu2TadRvw+AAn
xqTFTevV6K3IuWzcw2k6RQCZqQKQCROH/dfwlVeLb6ujMXhlOVI6URGK78ltyMvwqwHWFIM2kONl
+nx0qUUubaG9Gv65sbQTg6/Qfsu6FWBb7YjkKaI7pAGXwsquqn5ioykW1+Q7RhoiiCjvYNP5WSEX
knYLRt42IplEA/vv67bRU3zVmh3zFXtkCaEO5OUlXhvDxZpDMyH52SlLUOUrNITHg51e2bfAbh+8
bx2jTDvsUjAEEku/L8ImY6ZesAYqXfJYYCWVe9ulIUB/IsnTuXMDo6EHqRF0fId9TpDeb9SmENVw
85+BX35uJqFjWwKnwgcCTspJscGO+1cIZo4BsEfJROCyCBiCSWu+d87FeAgo4mjPSu3NYVRW0Qiz
HE7UF5fdvCH+v0kJ2TPiMLyHwvqq6nk8gGJ0IVEtJvcKMZSvZHJhlaMVlaJykQ/WcJjgvU3XK8qd
NNwyfjKMux6Zl4Ct1ZIDsaNBMWW+u/5a16E5U2GCYmo2mFZle39uyQXXZrT7/NrgDfOGpNtehGQ0
rp9rhfkVbETY+2qsEEyy8P8/GZHUQobUP1ohebNkfJ0hz6RzEJ717XPI6aI0l1EuIpBVlE5wkglG
3R4skl6W0IH4E+wu+lzuTV/rg//mtFbkEFLNGZVZgsih3n9nobpWjjo026flUgAsMaOqcMpcV3A1
6DJT8Y4vfD4f8RhEE7voya0v7xdRwUuUh2bGRblk9daxvudSo+r6kJiOD+FR9RlrGHbbkSrK4HR1
CgU0TJXbJLWvKFzAYra8BIYyuJxTIF5CLV06l8gUPctV5mRS0FLj03ykx+h5x4Mqd1ZpIyFcgbYN
VTlSpKbAwWsFpFOWP213olvLN/B5HOd6WUeJ8au/DCRRVKRKchAULGeSoXKT8V3vAlaMMO0YQlp9
53nzO7S448dH5mMpzf3HXGV/1hsfeIy3MLXq2ByDDhxdLEMo8BcJ4rTowePojhUtmN/DViIVitc/
smjMB8f5UmLZC1zydYIdCgBA7KJldU521s1vffcLVEBb6eSks/YSdZF0jtaCWIrvGoeeu84hBAkX
4qFZ9Xtu3qMQVXFHPstZ9/tnA/h62rnKlyoZuB9NoCzmltT3t/ayz7cV6YyhhNl9bkVGhSoliZ0a
cjRt9WAfMZw4Lb4SMUq//y11xXwtVdc1va+/d2Ftz7EPOCUHDqwHFp+GneGNdYLJDthFRTidRJ4Z
Uc8s8bX7fsJu6xmnTck+a9hCySDi1Oy6jFMJC7mDb0P+YUHLZPxFFQ7sZ+oDBKBLMDVER4L1BbmO
Gqik5cXXeyTOZTrBG5sY4Ppm07fmqOsImlGVG9b+gAwTQokpZa7tK2ZVcKUn8v25vnJ/TbkBogCy
XxcjxveI1a+G1PbTip1TZry6EnO4mzCP7A92AVQACRJc3NjLhvZXi/De+s0A9LwjM9RRSyF8Emq+
HtvYV4Q2OPgWWr/RmQ5HD5nTaI/ArJHKIaOGLhcMC1ThkhwaU11ggp1UVchCVaxqBPr/5S0GAQdd
deEpanrCPNcok7bIYTB0QOwdegQpk1aw9Fic6GqKChDtwgCpBpaRFKDCtnrewPzVYEpYDZb7AdIi
I3XtBgbY9ieFL+HURBdhCjjrPi0Wv+oePYD9w2mqvmiAGgpcYytOdOvryxQaz6eKnr4v9pu0QQ3M
d2nxEuAB+qhzv9iOVJpTed8x3WQjlspK9mEPqyEclt/0tgceGpzwBxC/G7NVJMnK37+2D2AIZN0z
m9l8b9I/PYWyROdGjX26JmRddCANBvBpUBLRbj0P7uCs2RlRLS2M4rufjJ0OBYv0AoBxyk4z5pDW
rxvVVk162ghGJA9VOjWlSRmQ9OPJIzCGP/nGRK9vYt5ODbgYL2ii4MKcu+kvNPhhGVKhy8g3EYi4
ohK0Z3XEcAO5B7XCkfQsVDqDHiUa1HPixSx2SfzTR2qFuAv7BEsPM6uzzeI/LtiSxHm+h4XCDSdJ
vN3EuGB3+2q9j8w0Rvkbk01ZaGA75704LU4Tct8jM1Xjw9TpbG2oMcKDZSQzYZzqVv4H8ygXhdrF
AlelpvU+/6m4XhWWa6byZl9xLTMFrWX434TuHAi3Ubps+CuN15GEgHacvMJJoT2QXRq8u2ipaItT
YVWhE8L1jq07e4TrpoqoqwYSg6rNuLInr87wiEwxE/qe6aPTiz9zzF+v/LPFv1pKNrlJvhoVMLeO
8ynLlL+JyBF5u3nAkdPyNJUIhRJO38o9QloXdkwdRkzB4IFPUqvCddX/IbWvrMfYwFCh+tOGrwKV
+bSEzdIr/QEQALkMp5YusdTJybP1vzP8/x7ggNSOz+Q+GA+BKP0aMsYyAHcNVFT2pR0kHoJ2Ft3p
zdt4HMsT+vw3TmvpJuA0nSywZNbJPAzcvcFNQxkTdn0d9P2zXfswlU0p4aUvrrh/rlb6N9ogqZ+Z
8fNWxoi4upmc0VVkKWjuNoh7JoMw3lTCZu5UYPS8H04X0ZxGExdMfMfVrd5kYNCISl5JU6lGtroO
nVD/xs7PzWVHACYwY+gJkY4h79XHVLhdSovOFDnhciYu1bBu/XBnogFDwVMiohmwIxzbDVm5Mn4+
JHj3ApegTPvHWOsiTolhW6f/vTk5GDM9MuKVGq64obygxf889N++qEQ59vfnQGpAwUQfM2ZpkXxA
O/VAjDVOUl9S8e199iQkPb5o4CHSTb1hHrhelz2NgzAz+I+C8Y+PQCIESFtIFXudEDF2BCkLsWSi
8fzZ/1cmh1IsEFkUpa6lS66vj6EF1EiSkm5gGkjc8NbzYoSSzGOwwAsdL8SVuOvbowyef/29dZ53
ea5tBmB7yX1QAb2VVx9fqQpYt2bVhpMo1mWwytV3++PcuhC3TUoSAvwN3Pw92pycjsSThcVgEKWz
Zqr01aBt9Bkm23G0XxI3LtxNK/G3xacpY/oK2Hm3vIHEevb4dhToWooPk5+KVEtPYBmyf+yBjx4N
kPP6HSD2xJArEgR24XjQz7h86YIAOnmVv5rJoXs1laHQDx2yJvlEc73w8u3rJxF4SbwOJ32I/NTp
BkLYeEyhCrtK74DX4fi/Cl6OQLGFad31a3P4/4PsYWmqgpzwue/i4tqy3t16aSqd3eH7oXWKLC3Q
GW4uCm2SPQjpDvuaxMfjasYPnEbU7QELW6boZ3h5eL65OO5eY94r/fXY2xsyoqB/x6pHEJB6gxMP
vpBB4KZLLdH2Bg9yd3X/8LlxyARPF4xIVbYX5cxGNGljuT8Ui/W6deIOV7kL4ntYVMFmQDGXZTaX
Xlx/lFXwPltyTm1HLyOIUc/0bx8bz63N+kz6mxkDYh7tmNDALBaI7Ay8ipXGtqwOYyECoJEB0/DZ
lPgNLCNWvPoVhz5CSRMhjuRTRjXGdMK+A5ORssoHNRLDHFnl1cNOsXARe2xRWUPXWXlx2VIYgp7c
xfjmw3SCrK7O4F7cfUq4E4L66Y4X9F4KnoVK2e14RMz1FLatRRRyL/ytsS6uMlDGHmmoU0bMOH7h
wjCNYEqfavYSCNEenAmrh0o6Hs0MvMgHeTUG5qJHU0SomqOL7mDKWCrxf4erATXTGnj1wZSt9LBH
udCKqc46jGGdt5U+laSQIxrdF8JMmJAcJQSPx7Y8c5JFQRuV5klZMo+/lSreqCWZoSn/3MEIJ/el
jXzMW7kD7anP8yFqKyTMeM62GUbqqgDgC7L9rnWLDmpA4NvC3JPIjbMEuQTREVkBiWHEZHfmELbX
v712ole9nx5hA2TQCFdZLx7w+g7Tw4jRrfVjvf5RM/bNG8nPHiwB7Ei6WUo0vkhfuRg/hKsYFaoI
o/f3L6OxKyZ0NIn9SBR0rFB/R+CHtQIgRzNL4UsmGxZi3v0o+r4IlRVEjpP9htbkhYvq50oZpzPT
OSaiSiW9CmzdF5oWJjOOfrTmytJ6s0cp2y0UZO/ZLAyNaKAOip95mWKl+9Yr6iRjCy5heNg/iLjz
QZnnc3zLrmJw+YzV1DtLVWY1tp/x2bCbtZGStyOB1YZ17gf3xPDR3eFiF5AlRypdSt6bchapESQ6
5i1/0bJA9Wo94xKpY3y9u+LqoPyA1NghHsfh9hACCBjEJVvxIQSaIdYMRZaaqC8OxXjEoFo4hkrf
N87K0W0QvRyfue0iHHpQIKu2dIQzYBQ8xr1GrIteBHczLVYxZOk1mA0zwNf0LJ94VYFh8eAflEOA
50peR0IpTOCTUD1AVYOuYeLXJk5nOnIMqQHk1qi4mHt6wpuu26KDQp3qdyFM3f7CHMyxvB81ySUt
//APHUfTtKWz5ETybQgx+ux2U+iVy6fuCB+DUqtbgO3eJURM6n5yYHArbnqd6Y9wipMb+5JwZ4bD
cPL1V/aOxWQeGkE/stt19wcC2Id4Xh0Aas456zlbzjaDhljWnrG3WPlsfIBGhqB48dumj275fTfm
82Rq8pXr+iv7QzxxGusqlDlNTwUWhW9z4pgE24hULxvORt9CpEM5TcwJLb2kqLvvxQ2RypmPiaHH
9N6BjpYM4obhqxKFsLC3z4M3bcWqNeWkhB5TjK1DZsUEgTDdOG6ob8RrFQPqKJqIZg698/DDOqa/
xwEkEoCJoR+3aQisiJINpKn6h2ZYfD+blAB/nVwXAYhNYDrpiw0g86Z6tqv/7d/d8xWYXb6D9joU
wHfWLf7H0bOK1mcH3pEUaX/NyBUn84gjNAs51hBlBhjUJ7U0Qbi3V5yEhS5lpuFg7NCO5dsZXD7i
+ESVFcXOxJ7nW1K71K+s7bGpE6MoDHo5pXFk6wALezQOXu+3LaQSF0+CrA/QadH+pVolB4pwUHyB
zdl5TLejsi5R3jFZpXIOx1t5z9e//xMYuiMPYcyRPc0afQJPCbieJJdTwtlgovw3RxYcf/uxRjGA
/qYyif32E72JtqB1B0k/1Rutou8A5LFtygzeunOzi92oHcmnd1ZsmDDuLIqQATENjPgk9UXcdrtw
aHm3ejSQO4RiX3fFmVCYDZeQ80cFLDx9U4EzREtJhDdL4Ig9YvniSP4khAYb7KkhJGwcjZrTy1UP
kLeJxBMTa7po58gnyEkOreNFhu9/PhMYjNwc5ldi12H2FBd096XH9irHxR3N0G6V3zUeMvTSjgbL
OkdYj8ZSF7bruVRaCEvaPGD43Mw2tWo6Eqzy+Je3sNOUb+2YhbDbqZNn+TghqqechTqiel/54ADx
cOW8wxaxgmtUJ16Vb8SoeoYbbGvQVAxKW2DcburMI1XZxafceSf4CMVPN8fHHp9ehHLzjemf/Frg
lBK4f19X69idSR7J2SASwmer/tjLclifsPvC/5/4lVZBUzZWcTKYasOJpcQBf5cn8oOWynxdYMDJ
ZFD9O0xo9ylbTvlycnKiu0N0uCWTxojHOjtVsPbTU+x9dNAM18e3MWvHaZZ25/WuvIbxA4OuxKaU
p4N6AlddodMNny9AyTn7vXOzU2X/hR4qduF+rdce7VkrvinDIATG0GBN8HcibP6STQ4kQVUTaEfS
oapOxRSi7gaBQk7IRSRPxyj7Ii8HlPhrqE9lTIi5q9cImSNDVyDwM9cLWNBha9dzWQTNyBFLOrgc
NLVgUs/MeyEdfKLVaGSdYdg3vn/6540aDtrtCpV6lTidEh9sO/4TlG36IE0j74rnJ5+PdDJG+p8R
9hnIlL0V4bcm8f/rTLza9gzhO4+efxRa8CXJdA33hqouBWD3kgAzL8PapVU9kPt2TytoOISgEJOU
Wd9Qm7hRdLX7Yh494oFtSuSugMHlba8vJ6/sHv8I2V5Wk4UAsmwFAQIPBfTpUgE36iCgtadjwe9U
EBZl/u1BZLkuLzJK59aZO9UyPlT3e47b30r9VxvUWNYm55uZI6CN+eGDWHMz86n6sJBA+YtoYPIi
Eia+0hl1AT54ZjW5IUg5DRHiv5Mv0TKZ3wdGMFHo6rrgZBrKMxBrUWL+py/DX8C42mV0los3v+X3
EB3vEpjRsg4Yf77Pm2Rv4RgsJfor9xs1Qrvb1yoc1yhnIxSYNpKO+F6+MM7Ifb9bcZRh+nRnfn/X
r3EH2VxOuzRcicQ2OK2ta8KtZ2rEWteICsdlKoux88NLpYAWDetGyAopbHGPIV/FAh7GFre87EmT
JfiSI/tO9Cf3cWlROm7faCg2p4i8nnZ7UDbeR7N0EEC5LlglUoGBbWqSsZO9b8HKxtMbS2sg7cxe
TXCJZXj8UXDixQEtNWpgFEtMBJkgcVZTBMjLDnYSkC2b/PYn/IPXw13JvlvToagwbT6Z75mmQKla
SDStSTddaaGeIrnVqnKCDBNVYxOxRvworKQcB0YFkwElmRZc/egxHZOOE3xS20iHLG/8X1EEJudj
xZJhTBkRRMXT2WYNGoGn1zczFeDjkmtqgnIyKOh49XLsJ/9tC0EwAMLrDoQs51Eoi+YzSGMR7EYk
h0NIeDhGAVHbKBCchZqXS4vV8bPRMYQDkFJEwc2nwly47YtORPHyGsCjVWsGBxRZwSNqolAnIoYj
+EYR4D0nSyNtCdA4CLJZNDNjqABqq195kXq77E1cMYGNx2Vn6jpncr7wK5DuAvuv/GHtQQWFN1F0
NxKBnD1+b3jPfFjYO/XdZVAenHV4wSzwM3RSHOSawfGbdNI393l4lhMZcOKx4ctatb71GHpqdYKv
gY5/CcybVMYpDUZD9ZPIIu4DdVl7VOSuQRylonZYdOMHU1Q6ccuw+VgjSGu8Ts0E5zN5v2U8J+mU
2AEYMi4a3d5FFvOp/4srVC/kvsvzRQ2i2NBoX/WgxLSFHnCKCJYQ+Efirwvfjq3fgR6TkwUZ4CiT
K0jq4XH7zynqHsNAlnv5oyiYi2NpRhZrjuDKf3lD6f2Cwpx1z23KRFlbLcpp5eUHap0q8fUl2b4r
zyP54LYWf5hxOlXrDyLpOYUJMpz7NvTdghy+SLtSEkRwn+vb+gcm5CtFVO3uISpsTToet9JBgDkf
5p/YGM9gjM4xrWMGu1md/KvjSW7Ojnlza2a1XI0uHSzpfX5TBgXOkJ3azj1fY2aIunNUWm8+OPiX
0P1A3xmsua3FZ0IEvYdBcl90Y3pgPWDQOnFD5ZIvsE5czrDI/JX9G3sMKnLHQkzcPeZRyiSGEdaK
vhqM7b8w+06dlUWP43RHRQ7uqVVKql8GRr7CTuVrl/jY75U0/lTcwEWmQadRIlt3NKwY+f8BgS0t
eNd7pDE4fzKsRV46DsHt0Lj0sCCUQrHpK9Kqt1I/GqZNHfgtSZOEoObTGPAbnf22LGRS4pM9y31x
XjffSH84sjhXtFT97rvcJq7DJkhimsFuJOO7zbO1eMFZiFP/cbyl5CsB3Fdv9SM65dhhdgPdXhk/
oMOFVjT3siT2JkCVJjMlUzc61+11YG82E8m+9PXozNgBJACjr5GHjRTPP6EOWgOL07Y/m4CuYoVI
OjfDrOTont73ze7X0I15VFYrbc9QSxfYW+9KJd6kIi740lPO8Ham1UdMD6wvMYChxDG5d2W7i636
2KTu5R8m0XNYaRFKcLfKA1Ws2Q09oBWaQLKcVMVDegNwVJ1Set8bmpXMjc0EDFwqBawcbGCtreya
nUa7L86pmjsZcn1n6BADsbXutGsoPaY1FEofWY+AcZX4tGenPi49+UVO7t/33PO8so+sWZLC6cUY
IdKTSoi6J11km7N1cSdZlp1xqjx5MNG2g9yyqCofz2eErKPg2Acf6+Dh7IhB7O7YcxLI217XNHg5
zH004aN3FPs9oziyryo3M5FiJVdfSYESeo02e5x8dGnYaYJrLhM0RUB6V/bwhrjsi/2H2ia1v6hv
lYGZQDCZ/0tME8jHTCs/OGrx7eHAajUU4KA80zy1rpQGry5WL6HrZJzcDioygjAj7/ETAe78u4lH
tLAVdYoiaBuCUaHhoIMqPXzDKmhWFW7FTZ3kzsxLGztHm2WFfrCGEr/WxwO0YrBtZugSH5WVKTbV
lY1V+2aUc6kXCtGPOy3F4Sts/88TAmKSaVlGvq+9wMsRu8kRTWsqgFrXX4+7x9BUUP4GOBBHutCT
7d49V0Wc8mKTRzNRKSfCYdqUmICYg0pqBbgxPgzJjn+afLAwgDrBsR5Zpcr6U8sEKVCRozbe/O6d
UXzDCwG0kx4TIF7UyqMB04WaM9GAlwywBejAVMDvFG7E+SlKrLTSxXzLnuDP3XIPMxN6r1HIX5eZ
FlYbwk7z8c2DE3ub0oad7WaW2LAn6TpP/L+Nk3DAmfAk5qU6ELyi
`protect end_protected
