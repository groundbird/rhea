`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VSnujw2zIGakDZtn+Isu9FyJeHx7Pz8U2bDtI3TDO63118cT4lX4GS/uUF69tsNeIYdtqQWMa9Sr
G3SXfw8DeA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M+UNyhXCe1hknfqmZ0Dmh/RIXszbZSHisHMiBCqJB9Z6PJMcE60LpusT5tCtdf6W5KhXoY6v3h0Q
amycXsXtaQyVn6ZnxhICH/rj0VMpqktxgfErAHe+0hyFYgUz5xFWC27RAbPLw2oMiGOks4VVe0nF
ELLVNDS4U3svrFtI1nY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EXfXHlFt7UAG9nwAKAdyJgyFpGU7WG54+x2bp9UMkt5mRjtv+A15WGAITbQK79Q0NpyxscIazDIp
vrfAF1mbrMzzg3wngBLvsc8GDIVElgZ5A1A7PZB13VyoO5H7qo5OK/xanPESIxFNfkTQ92ENENe/
cHToIJ61p/3gAmJwuKg1t40skfoLrJOHVpqOYl5HKIzxaER2xHKnqMJN/lpDHDCT88bOl/rJ4NJ3
WiwQGwMkfdvzwbZrx8nOTHC++BtESrmxKPgt+QxjXnApACHr/aBzgYaELqyFCZ04Q8WVJbFdr2KP
s4/cbGZOkZSUXsiLPz1es9PBaSw1IU/uypt48g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sfBofOCMECSFGZnGCAwAX+n91KylIDX7mACGkt6LCBWJJZ2SGnoXy46k7Av0mlNF3mrPNm04mCs9
E5ee0TCpjDlIvv+QfgLVAFJMBsgo7QXoBn4JKb47gO0arxdCt+aacglAC8RfEHuQpTEbFWvSfMbW
IpX5Gq4FkV+pMLRH/ZM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pnUMY1e51hghM3aJ40NgTx2kb6S+CLun1HjPAkgMG63GP+mGipqD7mGB0G10Hk7/A0Ugl+/rgah/
XvEvJcUwMwQxSULkpuDHQq842d5l7WIG4Hnoy5kcct0yo2yv9n06RCq+ViCMoQQzrk10ZMyK6s3A
TPYi5n5PVQ2n9lNCr5MAu4eUDBTCPsIHBXJ4jT6eZQfmnWTwYq6I+zxac3R39Sm4tqnWpQQlz/20
XwUylcTkjZNZEU2nMuV7hJWZ/XixLw7DwlEWIiC4upQAYZvOLS9jtf05SChws2EOjQKFSC1uMPNM
UqA9RSRhhG9miyhCMlWOO/EIBgNXxjDOgs2VMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6208)
`protect data_block
lbLQ/X2y1BhIjtpsI6iSYCpHQBZ34lzTrsvwmUQgWfFogGL/suwU49hY+ePkcOA8x5QCSs8taRiz
wnHIYcM8qrN7+dceV0oVg/UcjbgKbUwAb1kquwpXY8Zw1ETHI76fTgBS6VmJgLnU47LR1WWEGaTV
YwXAvG+Tkqd3P0dflKgsqc6mLEfv6EbhjyoOqe0Fehg/M9AtaQDtztchLRea1SvvWSTsO1CV5yzb
9CiZv95tnw+jHJLWfg8cGMkpqgYKnHVfWQKMNlKYpRVL5jVeD6kHvntlfUU3G5bYqM6qXEnfK8kH
BScsN/uEDWJ3a3vpDStdHeoU6hrR9giU5HTCRKPahBRC83LOcGOVm+LK2FxV5y2UIKfqlAQsPshx
FpW/GXpCSj2ws23Hmssf1yjqm9EnOZrrTyRsWM3vIkED5AZsNZHDB3H5vHkxhq8p9dtzF0Y8sDxZ
VJYTcbg0H6gRF4z//tJBkGEAerKQQXYR7IforXgVb4dYmSLmJx8kBzo77WcUGZT2B+PDQRPBbQau
+CC1VjeFzZkw+KSN9i2fv8CLvgwm+vgItCqdkL7Vm8ww3l3BuRPeiye+OWgFxkZ+OznNnrLRExgU
nyLQt5y8JrxCADxVc5rMBygQA6QadDPaQoCSsCF3v0wmVgSPfSiXmKnXgu8yM8KiHyyh/ZnpWp3r
klLL8MLYmoqw/9EVLhjamdIqt5CyrVZoIljeWcXY91vdfDBBUqHoHkd7GDxJVF+T6dMcdyxf20aF
VQdR9JXYahmleiknCSxpOfXkLPfUkoPOpO+DqRL5QZDuIsPcFDjlOYTMaJ1goDwaAnQX8IZt9GQq
zQDMfQBjLqYoi8m5fqmdEzThSrrNfPEpsZ7cprMSjofehCuYvXe4Fqysq0YctifKjCL22iJQQiWL
xJCm25mPMXElfs1xic0NBf2c7PENm8l/l/iBa16YLAjxbbVhMYqaelc9sHm8EkBlgnzFVBrKCCca
TLwHdvMWHpFo2vVYTwXj62L0xvcMvoq2LNOM82gP24lD1RwLCKC4EeGyBtdijpIQxvY3f0oaqBg1
g4oXoKqXt3lLDEzI2OAOMNUi3CHH3RZQVoIta/CpM9Nl/ujw5+/+IEPdnbl/rBodzZn1yTMphskl
MLmOoMQ27zj83+pmneHGyMl99ie/Qo61rxz081DsuVWaW9s18d/tmB2JCII2/5pE+2VbbVQyE1av
31YNm/qaT7ZNIy/DRs6TJiCaKu3FULEpiyLg9ZTLn4IK4wvdQj5Q1HvuSBiG5iEX6bF2b+4lM19n
m2Z209QTlBEKkjpDH4BM0xlhSb9OA2M5Cgf2ggZ9zPh75BsDD/rGrZ33I/GuzNw/cFIfV7FQr9Ct
WFtiqGz5h20m1gGVEbCet/VS+yFh+pTJBwqX4d+mIdjhtiyo+aY/gvlmfqijFUeSC1NJL6jr/ia5
m7oEXh3Fm4sbIc/EnYQO0kG2SHWcQsFNiiOOnUeWIaQxiPMMrzaJu1AuUcsGmq93g6NV2RopAKQT
r5huc1exbksfsH+NQnwPcErL3bOW2H9XNjIAX4PiyYr/e604kQz8pMKQ/ZINL339BHmOhJFfJVeh
MSTlFDgbVttveiv9XMMAh0NJEQNb1YuI2qqvsxUfmbtUqMHDrRa/4Ez4yYbGbpyPNQ18v11E25e0
1KHab2tDMwUCN8IkjFI+FKLzNXCXVnb7Qsor0c9IKMAo+oyvI49CSzbp0iRdxNcsYe+HeCkHC3Zt
qTS77hag6bh2d05JqKj5fA03awjMXkvwObFAicMoLKpU/+7ztjQSH2R/URDHblO+vL1YuXavrF65
BnDQpOpm0bgMqLZbLzK7sMAZEb2SiTGatWXCfe6c/MJhNTFAg8JngAcrr9J1q3qnni4D5hkZouqZ
7dplEm616f9NvR5qulHo2iebY7jWbIKBIoV8VPglwA4d00xuZElHza1Wqau1LE/COcj8gIptw5lm
GjDhdX9HzeWzvTnuTo0B6INiEmFoLJeZ9TQvw3J/BPIAQVEck6FFrcV2jhUKq1/U6/AqVZ6jqRUI
VKsdQCcP6PGI4dJNafVy47yMkYMZaqhUVMfEE/i2IBNgeZUfqql3Z/7DkAQutL+4KYsDWvWNTsfY
T3lFGyLoLy1Ntdiy31+Sx3D1qyqdpIt60jT+4FKEhHcPRJGu0p9hrTSVI9huagwF6nwz45VYY/C4
Sc2Vu8tNIK4d0HfPUyepKzGW6RuTwIPDSMxcqgRv6x6BIOppilo46pfAVEwh8wqoH0STCW6E2b5f
hpODtw/R1tM9M+9T4MqO/LXmm76P/ssc7lvK8SePgOaLUU2OjYhqN6eTwkAp1/oD+xWJlt3Xjuqk
zI6FOBqewBhS8Zr6iLqpWxZwZH8RwNt+K73QTj+hqFDRzvDbsjkmj1sVP643smwG+uASq7SAIUTv
ozAAc/WgTUPEu/TIiPEufXe05T8r+DuXl8XHspM1EmzjkKjqwoRwq74s+uuwKZJRoVi1r1FGXE+h
doPYaERkxtu5XZGHCR0JfI3bZU4mj/woEfbldcIvYhY9LsoqQlNnWIpD1WUAhOhhM/ghZEw5hcZ6
dTQBoVF96ibnIwC291EeSA462NbSvJosq9x39/EOwNy3QRKOznjd5ylX8FoF7j14j7iULr7T5H+8
pHTCfz2LCWFROtthw4hxgO5OGqK7wiW3OeZxDH0waOA7ZSStV+GnBg5x2PBGhfd/FrFIHdw3jaR2
1jKpiuUXCXmn+iPnCWfJqYgek1t72qKE6MAN2OwdM0TqWVqhVHHcBK9ra1g4XtycCCM1zRA34qF3
HKWhth3L6aqYGFbIdulCZ2TGl07noSu3S8zjdBK0XtRBqzPVlzDJi6PFiHrsyl5nkFF8kVQ+kqI3
1lS8PCcrMLmM3D3XSUzUQX5nGjqc7xSJINNguRaVjs/Ynkp9FYHNob3dOxZSL1au8DFJwHkdId24
KMAXk8uFpeu3Ioc7Xv+8OT9mS21+7+Q7+RGiZv+bBzp1R88wTpsecLSEd2LHQ+iRYsTm+7rUKaNW
O6DMFPBP+/jvhwjz6EJQz/ho1HR9x5ykmBcX3EoTuLqpDmxtbMFZMALCB+sYNQJ3ZYjFIexM7nJh
+8XGDZbVxtjqaQo8+x3EJleojCOdv5BiV+0VqkWZcKgt5LQKou3wy5t72n7ajiAAx8PukBwVXm02
QX4RCufLGJrNmV8HEnCNzf/mm7ATZH56zTP0KWwOkvg/teuw+dp7TDu4ltrE6a8ILd17b+LuhT+u
aHOb0qy9tOVNMTOmOUK+CuBfdJkijnkcZ/FUBaLwy9bf/PlG/nSzF/4kKCWgD/pi/BouIATm6QAe
b2WXotwwm2vjs2EPpx+ACkArQAggtv+ZXQhtwHexe4AXwEyFOGMXoWtw/3mBnSAedsGtoNutAxtC
owsQRkDwvwNqC47i9YL99Zc1VBzyrvG+VhzDkeyOZkcKSB+Fa+AQprYuH8ixYDZdWExfplIBmdXt
an+aiDjvkSGtzfgveXQv44IAtHBIlRxESugIO3TrhwhmepNTvOpE0+z91oG2ygj62CHeYkWE1BH6
Jf+IO6KYZnEmPANc36NaqmtpqcymoBxbNK0rkQuEAAqDatKq/644KFyp82CKXQrrLSmtTRK6ZaJw
SYOROuxQguea3obfXbSHSDzc7l0XExtuiLJetAmDkIsOzwYAI50czRCf8Vcxs6P9x4Wzsol7Tn4K
RJ+3kVV+GIf2BG7Mf8+snWdM6QDNxiFq4USpT7L/I05rMqy4OPtOpYBZjtOKjg5aEzQ1LgAb9jqZ
1h728rVJ1A+wA1KchW02nCuTSCHh3GdWCCIat7ouTpREA+S8b34sPKVqaA28nNwvu4cNquTHZviv
b+tzDqPQToG7PDF25lZacIX3nt0xdlyVmRI0Ji1yjOHOqEF42tPlDBVIXKxvYkBp1ExC1W3ElYgV
IWnYAdZGBZ06YeelmP+8E/u5DSNnenLxpA2ifdxessQd9QgMLGEYaCD93ViCgowAoGAUd/f/Dmry
I2SFEDK8iEtSieKbeZnx9TpB0O5rwBQPjti6yYat3Vtmlp3gITa4S/IqST6Xqf39YvUiRX2RdOkM
JQLKAT/v0b6x9UCeAYWAoAA0I4UZRwnn/sm4mN3IFE4D3WYj1k2Vk4hoJOXwoRpRT/fkSX37sKZ3
Il1ql0rdsiObHcM+lQAQ5+oZRyiKsRjMbf3KZgUbwwlDW0fzurEnKGGyDDGZq7+IZqChwZbFK2R1
UG/R3WLGNRjHo1lMoV4U4BU2z3Vd0eQIZ1s6pwIWhU/FOfWuAhX/lDFYccfYMvH+yXb85fdinNc3
Mz0G4f5tTz12qYLjxdwAubO6riY2Tsqa6FnjWnI84Vkk1IOtGX5vsR7oer7HRR6CgTrqG5UmoBJF
ED/9xVhgI6bIYTyRAxAtpUEKyvGILmq92nZ7VhHM7Uv7NTsRcMdhf0aoYel5avN1FvsiT6yEmzyj
iGZpM3nvB2An4B5UZFK3A5yc5+b0gZUpt+ghy4TseFia2pz5t4dLS630RmlxmHX1HelBwFirpMi6
+nJPAvN/jwtPj+BWqJveU7RffcfQ5mX9/yGjp0kzOASAOfTYX1D5g8/kmRsreDrWsaSHvOwGsy+G
qaY+y03mBwQgqtspe+1eiaC4JlxDf99QMnSsgG/gkz2IwtKXuUpbg8mGeqSHkcrISKQ8wpUT7Gfh
QifuzDeg6fiExWfkrlDvaJmTU5VNxRmKsM4ycaNZbGlEl5M5flCTsK9AxEqaQja4vhtLVyIGJbwC
km4q/3qzVkwXoe64sI5Mf6PZ44nF/djZzq+eDZ724T8Q+JVqjwUBuI2/ue2IS2E0cRl4m/RL6oiv
OJ0iDash+O/U2BZVSY4UG3/jszRcdmvcBUYQ0ZlbAudPFtjPMA+xdaNJunFNiftByYF7uBn52Mrs
GSAz9a4Gg7UkG8nST6ISHDVlAERCBvEMRlxyrOvt14tNtNXD27i0iE+BBj0acKf47eazsn5AjnKj
ms2FWnsIKp5lyNHHELUCzuM/7y3ep1hjfopfXk9MYuKGaoToQ3A6e6tZaHMZXbuFY4OUZqiJezpz
klI+PnvqFgNVrD1Kh7JPv5Um1zeCu32nHgl91GTQ05JVT037elcQxf4498iJ8Kx0xKipUPHo14M6
qvGmPmdk2l5dtU8JzoIMxv0RkpfqE7fcfbBUA6JW+GPj/HKJYqUxMZtgMnhtmxu23vs0SQKjS3IF
FcSfhsbvka8fqQVUDNaJDUsHmbjRzPOhmwjBbQSD54Yw5c+zCgqGWXCGXt6JsYSO1MJqybarNxv8
69Y+E8VlVd0Y3bWyRQCytxRL0wq+bcz3o/uuHHc9lUbyDJR97JFfNQBXdFcoSm1nEF3loM5hh64D
z4MfhBPg44DqdSgbMEN9unv+f52djMexsOl4nDaWJYKpIJ76MqJvSp5cW7EgHEsVFo1U5q/nJ1g3
tE2jgLOxaan5T5bd36suRNyGwosJyj+1TzsOsT64amZTEFxct4v6iB37tBi00DoFAHn04BoT3GDs
067s7L7k8lHOqjYARd5dD+n5kykhTLwjEbfmiBvawQFlddS7MDF4TF7WQRWE1yfne6lcsFpOW+6p
NzikrpMS04ziQkiwR+d6RsdxK5+sKXTYidrxVWYoiFHvU6jC6MpiMFo+7JmjgTI4I+el+qKOPp2k
yHUtI7Lyy3KKNjUWK7sOFfySQMbyQIaQg6UJwSW73defm2zZB5oDTW1/+UrYvw6Jg7gTGw2+g4f4
woImLctOl1+vcd5JY1JOK9QHRoqcTDHcJjFNP1LuIdDPsQ7Da0165d5GKvQoVDSQbOVgIvxqfsY3
Ky0gz6E+FH5okVMymOo2Ap23S4j7xXVn7RDFK3aMsEma+7vZeiDbcHJD6cvVwHZkHxde3u82weHo
fPSx81zfG3wi8dE94OfDUJlrsU9e3BCLkuH9GM9OrzsfHAmy9CiWBClo2XZuMy/+3cgyqnuDTmwh
OJc7Y3zawKaqK+9RyMFMjRZzu9267RFylORyVvbXaj3OyFNE4Ept6PwUgIZY0WWSbAn1BL8Oq3kY
dXxIyO9XQcGLT+NQt9925ueds3rBGeXfyaaWzBGZlJ+oAwbDnUrNcDrpzZd4hrZLYOzFFn4BS36e
ZrJCeO7B3GQeBfupRsuZIxP6g6+ur45hcicorr+glFU4s3H/UrurwMuRJdUvrfx4GnRfXIOo2pEh
ZNgdqAdE+HnsWnDbqlAraotC97T5raFvQTQFEquqf319BPtYJ6EEAZkOnzGuojDJ3oW2ZX94GCXr
bYPoMBYG3b0JtfNhoEIm2irsfZDXIfS0z55YymIIDJsw0KdYyHQzDCKJDDpOOOgkHl9bJENo8ZoQ
ym9EkzoE+GpctDy5icnztUTFnQ1XUJKWclsH4ea49P3mDeS4jnEh+Ikl1TN2XD31cbayT9uMkmY3
MVnOf255jf0w20NtPqa6HWrfPaODcREfH5P2+PSM4L3z3Es1HfhDbMom91yvSE5T6/smR/nPINor
pzKL1e4qVo7I17zHRrwtKRZQVUEop0G9/5dPslY11239Uuc1KVeUE9oTFn9NqWvevHlxo5gsuH2J
P3f0RytQmN7AuZpbdV01MtZMwzVv6B+JzDyDx1vQda4o7bFhsp/Ij8FEx0LZEFgSwcyL/EyNNlED
IgBLUGzeK47vZ79sscXvRwl9qDFebLIBJnqThVqmVW2ZC/aYXv9/xzSYFd8SzlKdf8vv4wxeDLR+
ZZaO7Tmm9KH8RJ6/Y6FxQRG2HQvTufkZXJINBQUsodaP64AqW6MJjnFVkLhbRiOlChBzyEz8zKCD
YfUoDHrYVFvKPHCH/Sdj4rSODdOA/JoO2KhIENwfstesiA4zGlBPsnUhsR5icjAF8hsSjEPVcbGG
VDq0jKdjrXyDdYDMtAOOFd6hkPUVmTMJrlWPB6ndZd0g/4gwAI0ccN+joQ9+KsnVqZSPqC2uZm1S
0/OVe375CgWKYWNl03jStcUs7eqeIalBp26ubJcPAgFQ3Jgp8rFAqGtowVOpRmsqJEnvw3pT/s2A
HvtxrTbwqf6YxC6XMi5JfoV6W+Snk3+eStos3QYmtimTbq91XTPQ5kXiPFc/98nG+uDVzPM1xm4L
DmnaUbfcWUg8yGDgMvPMIsaxWVabXMrSUXp06pvZDoXICJDmzwoujbzmVrwHbKw5qC3H693AT1c3
9Ku0hdMnOI9zsNxGQd8sGI7e2r2Y/xQ8p0CI0h7UcLGV9bh6awmcBMp4tKH24xnF7P5nzpJIaxwF
zR3t+XBDcRkfO9g4s3F8bZj5haV+GYN9SySHkVK/Y+EvNeQJjOrNv+Tfyx3VrP4dQvCIPRH+8H92
m6vE5lajuWBRnUCQ2HQqHlXqB80ODrgRA2kb76HKEp499aCJpuby+KgROPQBHRDVO5QxTWDLwBul
ywPuZ4dtxgApYpastDhjuWNsYz0pBUYBOHxTtFG7En5WDZNCJrrm5scOiQ4U4I9HKeU+fPsuAkpq
t6NJ1MzKe6PEBGHE8ZLQ2V/Sn6d9Aekj/4/Va+Me+K7krbWTpDHnQlN/xxAEvbcLFoDBj90KxV0u
zwei1Q/hy6qBhyhFi+fMTIOISZlElKeeTFw93wHsYU+ICqes4RsYepgtsP5pDKbClHfjHxzkVpJL
fKPjvvGOzRm+Hch4NWznBv99ElGpDJ7ddh2y1x8Ap0k53xoUkHR4zGrHstE8rHnvPOJ5feB8i45y
hl25nzLEsK2j6BS1eU68htV2D0w5VJergAue9sXNzPjaYNGZmiQNbtMQgy5MPX3B6HTNYOjKyH1w
0yMluA4HkhBMPeyFuiwrzqeGouEID+cbU2tnXfdjCxgxzy88LMeHlqI5tJ7+M/+axDdKi84xzdOD
eLfqyRpAt3t2WxZe/znvoYEuBUH6WQNmodXaLHQA5ilV1sO+YxYyXRMS+hOmd1PDU8wmAwjIJLq4
WMHItw/ucFmkxJnjdh24+JOghtIS26/RUEoQeJyW0ioNnFn0Xprmo25c2G5ZwVAGqVLVmj84Oduq
5sQnGa70kqHfH1XyzaMkm/XqqtavaCujT7qouq4BnCQyl8+zVFP8BWuQ+GCoyhM+cG6SKJL9sHZO
v9GnoiTduvYdwf3WqWJAkBCw7g5kIQPzPzUkP2Mrv2eAraXpyfALq4GfT8UjAQYym9Pjm6p9vO3p
hpzfLhqjn3t8PODjz+BJqAYMugXsAV/XfxKbCfeYu89WCJ91DeRib08ctB8fR7UkgGZQ7w==
`protect end_protected
