`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DuzNy6f0NkOJ6/FSahDHFcZ3UIBBtJ1dC6i60XqkuiCKG1h5jPafjynD0gsAgjHBJyJztvj9cCCe
DPAYjFjuqw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bMGu7Zdbg7xPlLPfXaZyuBNHOqNxwyqlaVWFR3DSNXQjtUcWtEm5dkYTFapNmnG9/g5UESv2JmIr
M4mYFfZ+mRv7/m5cS37QpsJLxIW8+4IUJtTOQ6TRiGHMUW8w0JLmxR0wyW7so1zbTBe30wUBTRkX
3W4W2z2g6b2RLv31U68=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iYsSbM/mWJYdCNMV6E0Q1MS8BQnAlQJNvJnQ2V+GaSGizdlmoXGpVejHAlB6Bi0shtixscLEO1tJ
uJD6oU5q5GhIgZ9FMIkwyWx7X3TrPvKGviRwsfr4bM/QT7jPGODJvx5ETplpC2DbI68QcWidm3xr
Qmc920KXWTcwB4/b4O3ojt3o24y0ueD1ylUJ5FOK5uPBtc6nskMVj/VUdr6ijs0RVL1vH0+5ymkb
ORjRE5echNRHc/EkdpWtCQrRRN36q0BcPbdQetxcmJcAgCdHeje1c8jN0P+SG6Y0V6UxpdcI2Ecw
VPN9Ytc3EMZLGDRAOc/ysuBqoyHmdILh4nbSVA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q+DSMk+pOahPieoRh6F0j6iTBoUQXHtFaCR6Y65HT+xn+KqVeWFbpyfcE8ObaImPDeX9L+65rrBk
WRQx1bpAHHihqW+ZJKeYvmiaNF+1q8o71MhMNBGlK7V+XFwW/wZEpPh/sfmNki8aTAjTEYEg1qs0
CSrlpiVU8yM3zwbNpC0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
seBuNz8aIOOmtHLHswzR6AKXBiZ94zKuAHMxaqnvt7DQiyaxTqW2ak5CyFvltaITJqRdWOfx6mU+
oj4hXDv/zGutEPHt+cDjd5fufZPKMtCwGVHy5bqxM0u4L9M1VTFfIYfb4Htlt4YhpHRcrc6admYK
LEECXj3iMK9MUSuoMIrsYYGb4cw6NBFH9zBnpgXgyiwpaj4NlfNZraGgVaDQPc3Lrr6cy1Uj+pyk
FyzKZ9GLPnzFSTAmYWth7N9JKAo4GEVx36CNskUiaE+PaffmyNYSfYWkiwZ1fr4Z3JjHo0NIFtpp
cuSH4ZGqQ3I5ZP+YTliyXyWekZGqxPmONH9xeg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15200)
`protect data_block
aLYyVPojVqCud8VfkehNjMFTNe/2pjcMnRTxiFwoCQBqazzG9J7Yp4JwBfLDGhDeJxgwIUi3YcKW
1TBc4ReGraX9aZw8fuGd2EYdTjQHZVz3uAd8B1XvCVai2pxAdFivFmy1JVhbGume20NrUgDLqOXz
qmSd2g/aWL4pZGVgvGgWXJD8TNfliyryC2F8zvDw20k67nD2gYfy1muN9MjizT/8Ka53XYMoVj/9
tni20y1C35lyvVAdpqDh/P9z7TcyGylF3M69m8uiFwyFJfwWvLpjJlHq7XzxKH67En9y5TmtPB+3
UOtXux1HDNf/2X3KSB+0RvCzQ97mpWIEmklz8YzgjiNL6IX+ntDHJhATPEeew0M1HtBbpetjz7Xk
3SC4iWjIfgXn2hhZszEzOw3mahTkiL6gTQbthnDxBcykwIuqk1chwfwjZgbX2iqNi8cq1tlJFodZ
7MQ04YG3HtkOQ7gexgVIw0ZG78KySJ2K5yagJbIHoJ3g2jnSDIZcE0xgycY9Vt5V4DM3idbfO143
0GViKWoFh80EKUmsSPdylcbi3/xG8JTod/QTVzoKtHDh6P+re6fjdXsBI1Gp8M32PoP7PunokEew
zlbMFH1DfJnOoqeDORupn/3nD5orzErB9v9vp88tzZAlnRushhU1A34JZsi/ZMBigvDa2qcbnwze
uRfbjgyOFpn5/VkctN5kaAZBG/QFTNI7Vu2xxIJQcKAsczVqAy0PCL2lgtZtJGlj6OIf0O5Lq91R
EGb94wz2eUuMETvjuXP06gAWL6t6g/G0ry9Br7KySMSJ1HpQbrrY3p1GIaZ6SywzTEjk/0kASQ9d
fmew0TejyzjXnybTY6Kj4sLZdp09rwQTmxO76JiKa4NV3ufEvyXWWGv4m3OIaGi9zbMLy1E2zpgw
VLMA9Z5xkqVY0zbYE89zMXwdSegZWBDegpggQlVT5bOehUDl1YT+9q25hRo0II0p8TgqttP4nSRQ
D9hqJuJfGKPFppabgVvky/Lh72X4PQwBMViSNQM9n5L5hdypH86BgrQz2gCuFXVic7Y1u23UjTz3
FlvvMfGrh/83hin2CtBr+ImA7/P8/PamE0ito57Woi/qmlV0vRvAPv5mAykfLg86X1MRVXhEt0H5
a4JB4LVf/cH3VEQwu5kKDp2LRAAaemjAzy1fbSGTq4/z5H+ZYKraoQWl2TFDKCCoKPAgLdJYUjDd
GnZDM3Kxm5+RvJY4EVU9cgeEcz04UTcbGp4dbKFYyQm00acUKYhuMbINc4CgT/SrLZSn+8arZHvo
o9/gwbAeEPJ8IJH+MEl+kOTz/U3dn3FZGzb3PXLiJ/fOQls5wJyj7TmcQjqx+0a8BwpOsTM1ha4x
Cdb2Otx1j1+PjePFkTYDZDmAaWe34QJymApuSjSQjP2kwQEGcfPDAo1P010OdESreMyninbhzaTP
NOXIQ0rAETuN6XR/Br2B1OyQXlZLKStKgnnjX5nYLbRJR0dPdTsz5RSzpFOp2v4qTKS+9KPYtfoL
XmXxwsd1jN05uPjwoZ8v6deenOGxB0D1NjBML6yoRZIgwwy/yWt8ksTS8ZbfbFrUeRubFCA6DxcT
ZxxSepNA1MY/jyr+d7/V+M08bEgMm1HvpW4tLtU/kNxVAAEWVc+IU4Wls5d4XNILfBSUlmGiOnDV
+fHlIqYaOOuWqM4eGyK7xe8SIYRjLZPfUhcekjODfeSXIv6zUpk1pchWHjdohO9UNgrZMyXZg0i2
TQUuxpM+n7omoWxGAKX2pKLGvWm8piS7CmryKWdw7/Z9TH+e4EzGqimfrXTSx+lyZ4vQF+yrj1og
0fkBbZjnpWGre0kjeiaJAs8HFVyjKt6FymO5qVI5S3AjiuJ11Cc4C08ArkjEM7vNHwuV7YbRvIcl
rNYj/O5e79dVrWCENVpJ/a5ORAGw4m+Y25+NY3joVxdlc+jICgAWoFT7tzT93Dypy91jxYG+mdbi
sQW3GvZoGlISAVSH0UkpuTm9qaCjy7CoCsm2WMg/4CKyOi4uk83K4NMWsXYoF9i0JAsqdFklsDmE
0MZD0Fk38DtHb9bPDB/NKM+VbYZNTKVhRcmhZeERAhCe+E5x2x+sV0F+/k+f0wbTb4RvCf/o7IeH
f0N9rPDth7qa1zrmhFeYSWaJoxkILbjFNvVIhdAK1TUZP6V7voC6q7oNHswEdo3g7tdlp5yElWWz
/ftDmm9Oufz3/rWkHBxsGMMijF/71g3edrXDKZ8ceExbS8DkQD3sMZNBMC51wm9Q5/nZF4K3DS4v
DOJVSpNawVcHuPiaKEeXILGT5J8IU48KZA0pb0qIc/w73Ijs689qTMeVGvQm2beAH2fo6CKiNF3e
k1D1c747QM3XBViu+vZnjxFFmC+ToOV+YqFVrleHWkOjfySo9hHyc+fsjmovgpqcpjyuBVRbrkXO
Q8ADDNSKNShRhj5nenfGGnie+p1AibAotcYU6OZXCKZIVUCKNgc0r2spZWGyaKDXe636GK9umHpo
k3DelfZdBZbR5shUqZSakWe34Foqfc2kHKCWyKfOTUjjz1G1U7xg9OjTqr/3EsSLZwoQzP1tCgcE
6FiNELXhQxafmnuef/CBlRTa/fRjXJR5glQJGa0lxXNKrY0d25RU9s7GfcfNEyaiGMW7bCz3ArzW
bmBXr/zUWz2KxYOJ691nb+/PqOns/lRUnYM2TC5x9y+2TfxpfGmQEip9qq4zCZY9PamaXmwwTcqu
tfHgFCSW6+sEp2qrTpb3JsghRDFfH4zccf4ZtOXKGSViZSpzDdFKtlQeg/Lpz4CmFZhBMxa+vZse
yd81wcbaHtw0P1AJoC0z10aRdWrmm3LGsaAM7AGqxyOP73RtVl24vYjTHlCxLGIYCRtCrIwfoWq2
dubPb/Sh9XsyWE/dJzXavyapodsBjQJtzENNOMr7jFfL5QVi2EpQdZBRsSOEF/0DF/jtw34Brz80
zNL7Dn+JWi/pQd7VWhDC9pTHUa95bTxqLXbcs8O3uj394y0ZIlm/vq+IhM6sOXe86OK/L8YZbend
vuPDbk5GN/6oOMH8Dn8C4tqP1JzUtrNRJwGvcJGQXX3Gtbpdyac+wCDGlcy18pHoI9nNtEk1v9EU
UyKUNbk7iw3LIuBkPrLpvuOTtTsqkegdHUu1+Gw45xHas83FmB4FhRCKhL+c0vuae2UzuWV7UTKl
sV5j+BundiYPfRmiY13uPvYGmXUsbcuZoCELOo3wLkhH+dSW6oMftqz76VWJ+xsJZVvFsicSrXgK
AclROKzAn5jvk81xQ6ZVsgpPhTRty5u0/n+U/ayanqpQYvMVid7eP2vQKChMbYJnalsLEMXyfeGR
FcaWhnVdFmI/NHxkpWPomebMAKFJF59UnaXWaesmWMIdqrnqjuWbmsAqWY9qs2Srgv+5ynGBE1th
PMH7MRfybxaiHFYMMw0GErsLuEQhBhiJ1ffr/YBaFSkdBWSRMqDvH4H4EpCOTEAqDA2s5kaPD2n2
RQqhle1S7MVeAHrm4BcJqYQEeQOtAlKqB23zQCV/1IBcVIhOWHWvLkfCkIKgbOHMoWVcVxRghBSF
z5Qz+CTUUz+qEm3WpDMDExyGuZNhXMsuRFDSV1SaakywSbe8za2PkgO3P/ezuk8nnlG8WN2dzIC6
/Y7Tz2ndQ7RdrhfeQ69eEKjIvQkU4o2kh+S/q0jVbGHiZVP6ETeSeKMcNeqectPNoAvfYgudU9TL
OGl2zMBGPnk/wsurAUaSlaJPpFXgV22+ckn1PHH6AZgVzcSoKpwrjeqBcY0uurUP+pvKrneaXhRj
cYshRPbr3HfHz7vbowvIqN1IZsVGm8N3qopgeuT96fymex6QvyUgb3D8I2QzFELrr9nKlvBWIpzt
jcq7mf0VXGeQLuz9HcMJ8jKKzAXtSCiACwPqzFmLgvlBsi+Y1BU46CYePS7+tNPss6ubf0X8bI1E
I+kIYUcvZgUijU+fKBsrRn24lTdH6Q0zuZRsJAXC0B+qAB8B2KKmMiIfJXeoww0fpY6n51HpedRd
9Lfs2HGKY3RJULREdDRhkS9vzG1WZRe8UIwzWvzLTem2IiADVWZYrzjp9DWUmwasllsoBZlSFNWS
zHa8JnprvCuK1tIBuyU8d94S8cSDNuRf56b8PkdniJN0gopHV1dHucG+caRNYnVI/qpOG6BDMsV4
b6KgSpNWEMEVE8BvfoLcMdsK694x9n4LvIhN1L2kRlqLOBgD9ezHCn85mU4+Aj2f8LJ6r5NwaVfK
cDdsaWI6pjEOe+fxoBxFNH4FtqNNMhw+X4wgl/jS7QrP7ujby0859Be9MjAmIJLqIco3uaOWlKi4
IFwpQMl9BJRMvqBEMuWpHHHQ8nZFm+vel6gK6d5Ak8A1jEVk+YEWq+Y2D2IUwyqOR58Wbx4I0vij
jlXWdieTa4kprXRGVLbjwyUjpCJ0wxkRQX04Hx4P1/wjX8MEn4XPFd7ig0mgxAItNxISFQ+730W9
uxHe0z8W3W5LSJLWkSsX1nZzE/ZJJiQsyP9SS+BbU3UQIZ958TObWx3fNrXyNOWkO7CfuUCQxtA7
/aLDEuBdV7sY0EgpCN7AGKS/8n6ZNpny7wmSwgjWbBguz1KBLmn4jKIDENKe2y9+jQia54Akmc6a
wmtJXclUmRG3nsk7Alhb77I5EBldAsshUZ1gei8AanZ4kY5JITtLgn4/EX7V1O62LwT9hdmRJu8O
wdVkVeiTresGJFVnLeoYZEA3/fVG3Jp373MWzf9UfPKPyntNB518+lx0AmyUhGRhNikOjVXNHKDQ
uZIXYVxsCR6Mgv2gPKSuWFy58kZzPu2C6avk/l3BVxn6iTdDcFlsYmf6i2XZprim4qyTaLtESaho
/1mGFQWp3U8+MJrEqQS0CbOa8a+9HkPEaKoPZni3KW0epOtqxHR0CAr9yRc+1TvudjjcY/S6aO7E
Kv4dxGwNpnOl07eARB8b3rVXhS7lfk267cPCy1OCZu4Te0yW5O9n7Q04krHCIOtLKNsL7hW+KpFX
Ki6vDuxWm5VB37yFwotyxKH20cihelPkWJj1Vagj2vxYQToaHqStZp4ntZ0TWoCZCphg6aeiYW+Z
WhMNMo+gae4hgSEESUU0ylDHEbs6RlHsMCFpxilMPI1KGsHoukF6MkjDL1xISB5YEja+2PJzjkWc
y4OEaV9jus+pWYBHUx0jtUtwF9ZFjo6SPW8l9trmoYBgO5721LbK/1jR/8rMcBqOFFt2zgghD/5N
AbByxCrKpSKtHv4uoUvec3/f4LZ44XVSmGUR3BxORRAweXPQz48/GNSEclFtezYgdTECnzz+avhI
58Cfdj6FG8J7mxThhk50mvJRPHsmPTHHvessbs5Q/on5tyVUVFb0n6Lk4PpJNDs7kGFoP6fz51Sm
x9pwTLspl0E7dslKXMKKPhC9Ro0/XlcxQyZVkvNSeaXCO1L9LoDnFmtWz0zLKeGjCs13zkeDLzHU
D5nVMnVc/bON2Ae8qTRlEZpxbd/4R6vjefbuSUHB14HMvBc+viC9N6yMr3mdllo0ubvD0I43uNCO
iHFvh0LUgEELAAPxZ845izr31xh1vA+Rt+wldCkhNhlIka5G+8R9sWZIbWKRB46H1u8GXOKormGL
g+W061LEsxlmQ1aDTVTOZaFkvPS4m+nYQPP7iVdYc9BxNtN+lBoRyGq1tiZwxRy3T9sJ500ouUT+
3qQ5fvhZJy0rW8Vqg7ztkdr2v6xR5+9wYpaK6iUKdREIJ/ZgvAYXaq/jbruejAPeD8Jbal5rkaR4
7Gzd/USlrIITrxqJf8c8Vm6m5mpSvi9GAL34sBzP+L2PinqWyXQz3r4BgwWNNmMW+fnRh5Daxdwr
YN9LNcKM8+AJ5NC7KquDCmm0kUGFPwiPsK1I/0aAOqxab24YmUCDmDkxSB2cnDW8w/jA23TkLxCS
sTWiuCgb9BxXaOkhzhigk68rULZ8VRC85a0b56+dbOp2sbDU0R2uX0SQk8AslfDHQCXhoz63AbjU
iLKk4DtR8CSKl5smrDT/+1xpMWWX75oWwlqQomRl3mfBk48A9VSA/o7PDFDRNkuLvhfFaJmfsEgX
vifr0X8hnb9c83A7aBugRcnZbuDoolfljHFjCiVU7P+sjjdQ1mxNstJKvHic8zjGF+7PCdVGcvuY
uS0Ju8JMb2KZf8+C36PTT6ovJ1vdhcA//yRyvtsds1GfZvEOs5PzaOx5ZcPQaOKFHTRvkCFV2lRg
IVxQGDp0lZd7GR+jJo34ViivWOF3KTAeu+zp3W1R3rt41XBndJPpwm46kvchP0yXVrcHTdKIS9Lm
XOskKEzkX8CgE5e9qqLQiIaEv6z67cs9XLlQvJ7kQIO9x3HaYhsjT1M+QgyhYHsSpK9q4lnXKjxn
GtSIb7Qj91xPRlx7svDR54fZwvnPYRLBakCBpzIMmUdnL5SQ67DJ0U2+SZWcW7y9pnwAcXsgytLt
XF04NB7gi2SRY0MLLClRkXi+sQDtuwtaGpvj+3bQNrrGBhivcxOuCJQWl3xaCRWRmo475hEyI6nk
lJdIEF1JcjJt2XOItcYS+v8yBHQs3yQtvuG5JeYs4Mx/XWuCTcwVq2h7TdlRJl1ZjupGVcdmGYlw
Zik4K/sOcHOn97vo0nFDIHkXLasEltbzYMs0Qwmccs6o8Xdccws9hxhQWF9eRJJmT2Rr6o+v7abI
ZSa+WmirNuxHCeoJjVeVNpng3UJ5AiG5Ycyb3sXbV2M037Cr0+golDpZkDOWxTDB7kUs4Y3JY0zz
RRyJ2DtYEIwjyXqgicUBov1OJf62Pt6H2l/MCzAgweByi0mqIHOiPDy3ybI8TYzzo8bddBiF8BVf
r5kWjlnOTw6unktToYs9wX6X55NCzm+i0v9cBCYYY3mJypxJczbs8k2cB80WJv2wu0bJwNEU3wwD
i4+brXKa3ZJMtWgyad/jexcTNpHZcoiqExUYNqBrzbmpL1Gkdgn+XfWruqCo5ZSX5db3S/cg+81u
7dp8ou6xSnKnL2wF4etTSC5I6Ozjxj6vDPiwyMzzbVqCkPEZY2Lqn7K0GViLhlh8VCMC+2Y/0deD
ZtPv3/qBvBtFC1IcjaIk/xD8mqL+xuMytTtg/n6h3S6rPwGEWh4ebH7Fow8dmAf/fRBYlb9VLDJb
AsVibG8SunPmJtlm8YDaj/xy5XkwhZ8HCAz1ADSic6E7UsOQWvMYbYoC+zjp7P9wcM09hpAPxT8A
IIWHL72tgt98H0omUWafdPoKwnoC/j+ki0HIpS8wTygx/g3uLuDoutpFj7wBJ9h0G5MYzfcZwgEG
s7N5EUQ7tLvPQpH6PJUye/4EBG1eXiAlG7UdVKg5ALIXl26Li+6oldATIb7VnjH0PkIaqsWhP+Zo
ECcSrKGu5DUQTbQ2k/v+tZ3O4BI82xoje0H1KXqECAK6nOIG9o8ddaZSzk+O05ythbQkzaxUMmBu
/drI6ar5sm+aIhCP8UQX/oN6y1r4lkvO6QANuCZ+v3TvtlAntKlWTxYgHBfk2orPGTR3Y3HUmv+b
1Ru0o6pMUBPqiEFWwdR9gh47w5sz2Mh/wCmdl2rnsaDRe4TfQ/I0buvowq6GOxwrmRgsNtYNX7GE
1S2HnjNvAhbnY/ABdreiRxN8vyQiP68ce33cMbPZVK0bLsGDt96DXjpP0fOeW+iYhh7ZFU1wGxLy
Rn3OW6VkE9Gr3N2U2RZBYuIXumiZ4coZp7PahtDgJIVQZ57sdRVqQgFgwxG072cSY5uNzQv8ibqk
M0HdeUKTxd7GoHuYTSSw2YD1AxpVJZkbM3zqbTMHplo+U2w9L+EdfZR7GYSQmdHxP8IoVxoKa3sh
EBS29mGb7G2UBGP6PDI0WArbJ42vG3/a4YXkgtQmUvDwnGfFJIQzkl4mAXOHT7+SZsugMQe/2U0b
gikpVb57FGWRKQ936d6L7iwqhjDbL3bZCdeefUE4ot/BCJXXjN9osCmLcjzwG6ww7K9S2447tUC7
9C5Z8jSUJ7xgqrdBbl6FSOdtUU8Xcag8e2dKalUNugiCbAitrbAggeAS1U9LxwrUojOOhJZEuFq9
M294DuvmweUVTtIUitdFsG0HDwENxSoup9Jl9rsfRD/wFQfMUW7ppK4WmR8NrVI+zoWYUZTRgcD/
TY4pzpyA1tL1+YwSl/+YCUI1zAH09WhqSoAwlRiw7qvyv085awbk7eR3D3oTRrTlnSHguUJm+VRD
ErWcor1744YV2pxfakKbwYN+mkGm+tWnDRCpUAE5q6YfWIm7wnDu1C18FSIUXGe/xQkOySc722Ds
VJ9RonIP2rFuk9cBBfwhxc37+/iWasn1izTbmAsZlWY5chDLvDxsm4IDL/HR1UCbcmbKTJpIro2C
vNUQTS6Rgey50/w2H2jLJFduBJziHPPR63N8p4OWykZX/8QSSOzuwvPmakp9VzOZWJfyH3A29eCO
w4zJn8vNkYu19PsujM1E+JE2z2TxdBClPRD6zBMyvq7iZz2zaTMxlDhevOWazpbyKO7xgAupauqM
kqXVYooHJAkOH1KSmDfcaepBfv1kEGPREB2yGAXyIApYVG1MZkfYQ6hrQxkdoenLJw7I69gsNvZ0
S29O0m/+TuCClmwDP5LcYY5wmGFmA76lm42Y8KD5ikeVPwJqYIRU4QSgOT9Mt5WSA1XoiZq3JRuQ
pZawmpgPNo6BzxmQ9sy+H487cB61dyVUKNu1vGjsn9CDLv/hawJ6dgqkN33A//ylgViod/wuGiwX
LELUxc3LC5vSft1RAs4U6+2LGNZ0rxxlK4QsLyIXt4fgSrlbukrGcBEewuI3FGV17/ZKCGxaZnO5
MvUt6/NT0Bn6MF1IbMdOWIR2SZsdQLu8HhKEfSnKcpD8jAQvigS9kk8Ery1KjjC8VYC/9PNZRm8A
LNwm3uzuqWJJihoN21eq/UQwJ7J7aAKZZEQYUAx9LMZL5tGuHm3qhtosQk+HM4hS0w7nTVJtVR1U
6YP4/8NLJ4vUiDtUNd/2dtRNlvesqsE83bfjH0JZBKpqjZ2DkSk85TE+fESo+O1Ly/fcDTAiqyIU
yrlShc4dtXERHIkVZ3nZvSYdWIz+Fb9zLQ3vS3aVHn/VWa2wQAzbBj96UUGkEHkVzhiYTLnidk8S
OtaSCigs9UOtDbe07lGLGQ/DzDcGno+Ldz9bsIgHL2/uDUcNdFQwQvI7gsptPzj15whrKp2v6O0l
kTY76h8gialpdB5BNSnx8Z9R1NrqleOdguH7DdHcYmU0P8FQnWHhINCTk3OauliIBqnd3Rw/q1PA
eYexl+cNWgG96wIZj3jc/uOyzFsnXDe39tDaADKZoq8odmxkVfnDS+9tVntQkmmnJ7imm0t5olE3
03fdGqMM8MFuO4bJ9C8qzt7Qz+e10CePf4yVT5/KPNgf+4BjECEEF+riUKsHEw2INgtFztyBskUz
Vg3V+Sj2uKtUYIOQf0KMuuyT2sulEIVt4edkKw9GzTEkW6MG8YeOWjn1fhV0fPHJnVEymOWidHBi
dLmKwZcApgjZhx0TQYLekPZJTPZc8nOFHqNRqVXR0aFbaj3cDT+MzWbwkQUr08QRXsOtfPJKnkzQ
0bJ5LNCIE6w7Wu/0tkUKItuaCp5+DDkriWvvEcE7DuhFjbjEfgQG7PKwRhZTcsiqSUccOIJo455y
HW+Las5hCembmyuULMkKNILGA0rPbuDfFE+Z2wP44EgVFyjqgaYYdJTNh0+Tez3lvJSqFnHwv1kn
PHkaFv/DZoXYqaQ9Fw+iPu17rG+u4P07+B16SDg+GJPVoOElRnlb0abs2qipq7PszoGiUB1IdwpQ
Tew/hYmicirHrTiFBNoLl8c/9uc+iShEOhsieYDgueKYogmNx2OxZxBoCNIcJOj1ytRGGJByH3gf
Erern1UtLFZpGbleInt8kSQ5Tszgz16PuTH/INjMFYxUL1EUTTghOYzmpURHp19UbislhBqlwdtf
qG5HVL4vrhAD/zl9S/v9v8ZfoIUJyPFHhkO+j9vTEU0pD+j+2JtMzl1c+GsBU7Cmg3EynIlSFRRq
PAAQGsGZ+4DxKqdp6g4hJfiWMUKPI1hot2r2wszBixMkzO6yzrrrjYiw+CkywlLfsrNShGWP0VAz
G3csCR9QQ3W2kTmMtjryYfzG9EWOGwnQ3a0r2HJpkdrk9x/t8p3uYHZEJmyjRdlJVlBwAzsOzFPC
45xrNJylhvmtnEzC0wOj8/D+iwEMTz+443q6NCS1SNOdkXA8bsLSjnOHI1yFYA6NKLZi01W05Tke
UW058KVK4hLEI3D1yP8EyGMsFG3Ell3vEtVVNplENfhg8ygN/7KgQijY0KGqUkoesb+swDGSX3Mn
3zsdylxM04BzqVcP6bztC3wRUObjKKvQi3wxrglgRnFA6eUzYPUm8ZFF6roJkF3Kx1Ol1jii+5F8
HJhbtUZ+5Xz5c2FDb/bSwQ01tlbgQTlgEuFmyN/XP/ZxKm+dulCL7xroLO1rv2foMjpYMhw9x0DL
WbB4Z0V5x30UQWXj9JeJOd4wAp0iRnzN4Cf1WEuQ7RxYR89PZV+dRXg4J/UBdxz74lVyauuAvdH5
KbBikCuw+ZNn7qIc5/TZiTid+n+4kuvvuj4jsgvo+yNpbua6NQpAELw62USn45HicGcpF/v7IzCc
n2K4PpPycc5QK3wIPufZ8KzTl6IPMFMgxGw9Wv0P73tSe9ovfurLMERtGnm/+Ci5DiAO+/uh//MF
eXI4XKfBtgH0wHtm9YABdtUXHVyPjHjTzlcSASn0DWGR60O4nVHRBwYJjMZ/PfixRMzeIhssh8HJ
AbQcj9FhA8RT06zNd1rD6eqABLaZ+hsiu/cKDd+k0b5Pj0bxchHss1/PR93mdyfeh5FDZHYSmnbi
+L7C1kON//7toJeGzjqyD6/ENsWXz5EACAOpRLOFCg7mJNNP2HxtdqrmnXJ2paA79ubvK31mWLXw
dE1aZ+FKT7n3XA3RWMozOjvFlkoh8g61mioEy+3v9FIIzqg35iWKBL7qNeyG9TPym/iGCtvxvrGq
2yG44l+HCImzhk45t1+gEtC0nJwiU3ORlFbLaArJJn0l99BYuqsSEP2CdOPln2ihnNzM2j0jUK7q
TewpchjKZVk2niF5P2TCjqHTse+sFE5xn3xAKERaYuHpaJfL7UIZqWRMeSEZQOh0iJ9nghdiShFR
rx4bnnKM9pBUebAhF45XFC09Y32as4TP+24iGqdgxsRJZrWCGNd6If373mjW/L/sSk9NJSUAevms
xT9RUGd265copf+Y1zWvHvhF0Jo3Utpd8aYboQYbjZHiUKMkdDpMMvslvWNrs2tFMEIfnhd3u6P2
uvr6M1CmF+ZCt/TDbZXzccrrqenzHyyv6XkjfMYUAFrx5afvjXIvXUqlZ+TsbQoPSYt2bV+Zd05F
4n96AuysvqAFOrJ+LbdkDFJjkEpN2aVeWfOWkixV6YYDUDnin9euRAwlzfARZfuj98Yh63QgymUk
b5RremXlSrs2xUmVWiYrKLAiUxHHOft0rZw1RlXqW+JonPyBi6VuB5TxTw5gbQjZ2A8J6APzyYww
QjrnzP42jYqc1kVEJ23+P6GfYHXehXoHaXxIlzKzoGJnuO+BtNz2J4bkOwZnfsDmfjzd0nTEs+Pa
ljwcBFBoVCzbjMoUdlRPqQhWVwnhzNEUSaWVdSI4sVTTbJgzpE0nHa8MEyy96pMY4FIAbcOU9z3j
kpcg7+7X9UMKPOSyMeE2PhVG+pBZydQ3IRSX/bIKd2nPDHg0qU71+eqSLa6nCzENAk1/+r8lLcr8
QZWfvMQq4OraF1svLIcrSSf/qfxT/TUeho/ZmMyoMt20DAvsh9V3C2Ro1QSsdvKr2i9ZIecNV6JG
U/Aaiufxr1flAVx20mBagpwtlY8Xmyeo5Y3OouE9xnQAOOWtzjK4Qu7mtdCjl9yTzwwCbN00geJ0
smrYGOQ2AfHk0jriV1HLjYYWtWTaTgjXz8DVM+P9l8CgrPzM0eP6tqditSd/zePVzrs/fxEp1O3U
JbimO0rIA1s9u9KqqDU8QCDrmEm/tyeu01Ng8YFw7N2n2Ytq6xtVqQa2rAts2+jRQTDOvqMKDJ9R
ElgMO/KPe7Tqo4YaqQl9I1g8no/BJWsmzVRwoXutGJs9RVvmqycEWRKeHLOz6YlEAAXi6Iq9p5gX
y2JC6nfSLmOxmuSJQu57cALcan4XWgXJOjitSmlEYgedm/QLEmifOjAGDZtoqHLKOkAN4bnd3/bK
2b5hcWT6FasN1NaacLr02PeBxsH7oQloEFTL5Ume5cVoPyXrMIi2ndR+kS3Bw9mg/xHBfX616aMu
50q+yzykLNB3eapJVmginhuZPWtq+s0M19OsUpaGzAzoIA8usuala+jUa7pTwDkYUH7BM+60ku2f
DWJZWMCkgyv4Ubrsq3kH3nDIH5ooIlWKpmHcnU+xZTb55XH0ppFiqLR+6BR/NfHoPHpAWycwyegM
dIgvlPmU9tNfWy52NT9nmoDU/DkZN6lNU9Qo2TgUs1+igF6FdcoQMTabiuHiWR+J2Rz9pHz94sm1
dw2TrTPjAhu+M5nUhegqNoWJsoXU7nJGFC8zmeXk7hYEAyuidj1bccYHsP+RUunl/1QZDUcIzm5u
O9DEwu7mLW+06SVhR14XfWHOtoAnSdrhYV89CNnwCQSrr95VLCoQ4pa/+jsZskJVEjPxBHgAK6tV
bngH0lU6lAAzULih5j/6/CJwXxxTNQJLxn8U+IW/GHff7T8mlOsqBzHCdJxL5OgQ+TjAHKcEcwKr
ihcFPM2dyFllzlKIMgjuL/K+6917TuFCXGrj2N9VXjfc690cMS/uG4g+fDJ3dxPOVEFaWyMlMFQT
S5CFaPeYnOVV0wymob8Ls6G/syuuDnqr4KqVgkbL2rrADACBv1yqu23t/1F2IdJmqVMYrBYi13Z9
z4Hx+e4NE9QExIyHote8vv0KRuxpji0Uk56BjyeYIJ2ZyzgprGR4kIgL22tq7dYFP2AZYmdJ3r6n
xdKqBO1A341hxMUtV9+boHG7Ejx7huRZc2YpiblS1QRDgGn4WqbTWCQj79O3NegcXbGmcRbwHM/Q
bHpIShryQ3pqQnHa3AVPVmEmherUBpvxejzOyCvoNkkBO5nv+F1IoDslcI+F02NlQlB66jjBjqax
Yo3MLC5WUQgbaJWYxAYFBwOmSGqknTpVmZqHcIdQW6GME7w8XS+AEJAZFa1jCz/etZTj/54u8Bzs
fX7cMWNY4PWMa/V0UaDTCui2DIXc+y0V4DRAPlSBicgd1oBs0Kv543+Ar3uORGl9p9KlAe86DQHs
ubiSxJnfk3OVRqtt9KAGOJFwWSbE/CM5EGDALa+5MEecluQShCq/MO/1CG0rBAR+nhcoCH+yjfiL
QYq+gZJexLVl54FPLQMeyMDoDH5d+TQewJ1/ZGXltsE58fy+OmA09CG8UHm5KOOyiVg5UqO5zDzz
+NH2K58hKdXqPwunCZx4a4AC5qSzWH2BCSpGaTqvY5nPM30yMB9W44BSipckhXf0UvZvVmGyEbR5
NquarRCCH7vVH9qSGUk0qiIumHBcpB+qROOEzS55w6J5VnT2s+iD/d0pU4ljAT7vDIdMZye85EyP
7LpMr+pbxiOTuFlC/hvbZae1houqgeaFXwAx8jQe5N7wQAtzS+3oh8s67ikAfFhJqgvBAZ0+Qybd
yWHkedYpfScG+4vKFjuWwyNRXvLYgmPdMPYw3o54wBVHpEjs7yZ4EOTw2RpvAvOvSKeC+O1GNY3r
2Ykr4wQxY3hl0DhVOxOIt3n4CFeBY9NipYPEDeocqRVLK9A/Wyzc1jYMzeZ8Yl2+hyG8glltWhBr
Lz3MFmYrscf8P3o9J6TfMnOm5kFAEY6vDyuGOraLKnuLNsh9GgpMyKomOhR65U5owlkeg/q8xEiJ
GVPyPc03uTAJ+Z1aIgAK6ibmhKhZaHwg8yURCtvaPjs+l6Qx8yJ5keHYFVmqlaK0u0jOsPk1O0Ob
oDLX/El+nfvhgsSdEAH0cHqFeXc3yh2KIJs8TAZkOUGiRz2m9QKBFm8XX9yEzWQfNMGfMu0Axt09
oTAFyG6PcvFOMUuF3ihytORhWDmHZ5KVb64MbtSYCldUpZU3chlz/tCSA3p6YQFReffFVYwldHPc
rQaQtwfda4rwywMD70QEhdHK9sxxPRPRvUHWtl+fQu/3Xv86wlaXhgZiNpWfUCGnn+LAS5fWv8R0
flSHS1MxEqXaIL3CC2/9iJBcAdR9zIYd8NxK9WIgnRiaQJrgY3/wpeMr9D3hokvUMTI1msw6Ht7D
hxu4xZyg9lOg4hz889b78ysHKypkXFKl4qnGKsQxsDYHP5IlZ+wQ5sgN8o/ncXqCetIRI0eMkY7o
YjfA+7pq6LCnB1gYjQNgRZsO37VhF9wcBLq7zIxkwi9BpakaTFq8CV8X35yvyXYmVZIpzu+fV1eL
3938iqCNqnqCzIEg5BLs+1wgS35NjlKHnAD3vHuvkrpEF28S1N76zfo8P+BxGO4whS4hAN9OhhCN
ly+qEVXQ6ttqPMJv6bWQzXluj8lZoCjxwB+BiWB6M+El1WC98FkX86Oml6xfwKLup1NMbHou0qiv
IWDMANWdPa7ePEGJXRsJ2EX/xB6Eflr1xrbumldoRwWKnVXrmVtDXl2nJd/WfY8sM8+dFEfmBdtA
KVg+NrZJLe7VnmbiVviwdfTKzmr89gdcttejjELFlE3CTOUsy3In590HXyZmLa6E8LLfp2m0B+q5
q4UuDIPvU1P6YPaw6z9HyuDORDHO84TPWjJCh5Cz/yMSx6DGQgAnuA/g8j+fneWwV26lzfBCB5K9
pGIvW4YMR4XDS0TVCyZ5iygH7QOZtOe2dLjIa8lcurA7lMrQkIelku3aiv/aPuhlKtWfzxqgQoWB
lw8jxyfxn6vBsEDxYaM+i8rUZQxTZ70rIOWsgiiyM28LUcbHZVuCgie1TOW+safmYW0RCqS8s//u
FB1FSiKwg/MmzlpuJCbYI7KJZxCIpIHvuHOCif8R382KOuPGlC7F9bcabw9n4GE2cTOq3BGmkJxM
R3BMnp550vDFSy5VAjDRWSBdB/YUxrvSMe1sBuykBFwOZ3Cbg280oam9f4kjDDGnTYijXj7BEBpT
+pZjzvSucfXfLUydI8G4zDWB1HRzUPluNu4do0fDRhNpK5ZRyuH9laBQlVbnxVSDuN0HHu1aoyqM
m1WfYO3TkTJ48tk6uJpe6f714q+SVtLc5YuyUs7r/aCrHd89+NOjRit/MX2/NCkqziciM4vzfg5V
rye+bOjTV/eUYhH44RTVdnk6tKG2co7/FNyTZfcN3G9B9mFqJnVHfJxGEAR2KM/5ImMkJtrHnXPF
/fgKFzOiWCSf6pFO0O5tAl5vhe2rPlpcsouxjSg6PAO4CDIWestI6P5NLVldC0pTSrI+44W/4la+
2co+pynvh8h0TTc0/Nd8jGAqDNnnn/yduHXtEmLuVBswIMcxGgqoJ70KM5PCpo3tUPeucqVVRV2e
djbfVZIShVeff5cRlY8kXdhe7JIU2Vb6D4vsgSHkayIvjosvELncPiIDBWOK+Say48GPmT1a09aN
w/oKiRyr6f4vH1NXz/py3Ko/D2rd5w7gE8lCany8hsneMptJ72EByr7r5jPhDI+FrpFaOWcXhWya
clb43cacPcQMJzsWCPy3w+xtp2WSjQInGLXO+IyaheqpWp60JdZKnAcBwvwdPXpr3v+jZ8bqWtUh
+hQn0BYaeAFxBQfhBCHOdXTkOs0C0H9dXZ8EeLSbFw8NfCiSQxDsxtHdTzJVAB4/LZefiDeguGpW
iRRGB1Pj17SzoS2kEmIsKo9nns7+SV5ARiJBVyIPiZKiS+4yw+gRy04r1u1kGMPTQ1tuwizqU00C
vHPnu2zla4nQkmTU2DtFeXVniuMErxnLyD2ohVe5UDjLOGFbrlk+spKjw2tKCpBvrPd0Q6yz0C7E
JYdSdX8ypB6nUtrzwVHw2YLO4q+/8MMntIfgEJEUNUIpgtvx1CiVMoVEAPjspin48lz8p9+X/BB/
U1w0Uwr+B9f0wNad+j+QGdjUru6U5kJ5MeYqql4BRXyvCPymKUBj96ptWJphXKME8jK/u+BkVimm
KtwFuG7cVHXg0MYKBNdeFK4DPpQd+st7Jv9MBpUapCdGI5NrdvFC/yTIeAHwmiJ3xHlVsz2bZXBa
uuTwAmbbxt+oaK0KgoCbwvPA++mhAa/umK7Zw6OGqsyCiLy1o/rDptq0abqIvPAAebA+0iIda1y/
MuS0Hd4CCI4fhekzLVv2op6CY57oy1tGWfU0zF5hNK8zoAAUneKEz00I7qAIMt0RURdBbSOD9EMm
ZkorVS+AzA4Yp7ZrwQ/X38J6ZbRt2Wv4R2F+H8U50k5im7SI+39D6gdfWBDUCSkFp4TiS7zDBcS4
dDinxr01lHUf86KIWuDt5T4Htqo3osgEDwaA7/qpLJ/z8w02Ts9zejpbKtnCZHW/2ZkB9BvMWW2q
nfwK3Xe9g+jqDBGRuh7NP7oaWo27OAfkaKTtW/2wWpN/ShP2+6n3ar0f9k0b4/of3L5c+XDTddwE
KYf7mqwSxTgrksOY0d2LElOxM4QpRLQ4qLq7mTjANj+tY+wyUc2VNrwETqu0bbspfX31VSD3DYkP
VqKexWn8x6Oa8XoZ56i0f635wMseuZGCSzHibNuIUYRsXpBYfcfVPZ4/gO3YemrjuGxiXN9RogSP
6jlfLbQCy/iguxG3+CElkRcCfBjskLHZLBx6o08M2LLSSjwVOn+5NEHWKKYCHdYIl9/fswILj+fQ
nMnVpYtRyTUOvtNqfUkDSnisP0EtLyW5msB4i8mJlBnZsGsNQGlZV8uxh0QSKfOLY3gI+PUAIp9T
whHwtosYnEVJYGWCbSMEovnUSQ2uGW/mjfH92uAIIGQM3WGS/IsmL/pXTcGuJLcfOFp06476HiTP
MTH0/m4HRCskbuX04U8ZyXiCS0ddJE8aI5Ial5jQdMmrxCxjHtB/cP+FZV0Jr5rJTg9JvPHH6QHD
vgdnZhFkOz0VICqxGmbcq1ZfPmGstjkbTwmgM42UAaNUMkw4BgY4MzR2YwRDocMArpqFbFZuhwjj
96wZtXpQX6Ju+FEaNd1LYvJ1ZeL3LIGxhuAsWt/zZbzlmRsN8E9YANAq1cFeGhK+HVcvEvKWKi6K
p9tDc3VfaketWkwn4ErGjFBNZwKb3Lh2l9du2U87d2d/RHFP48uOUJcaFeYlg9nzDkjWv+0oQA5n
XV+mqUBOtBqrQBCpV7/3UbkUp8i66bH6TCoZZ88TzkDf+xXnGUCitvyCuEq/19hbBPL1zmXNgXCC
p1+l7gGVKmXLSvPaj78V4Vs+n3F0iRbVSzLLlt2FvOFJvX+iZ082/UE70XEGFez5FQ45THhlYBIk
PMeDzcKmv1gsEKya97KXtMC8lpIZn/OKLMDne6GsKAX/QnCCCTH6zmVVU/nJgRkWO0JTIqcsTUaM
xJmGG2NxDw3QVJL8RqiZkiUOur3tqFdbqI489capkPi8s2fai4F+yfFyPW6lIs/a6uNgVfaa9uL/
spfU9IxdZOavW6Ldmfk2gnoDW6v+0T/2WMaUqX1wevffU1MsLLqv7m2JmLco+SAm74kDeiM18W0H
rtVG1oVV8k4xR7fsvQSgFtLY+xs7F5i+LTbdqaPWctGm2cFLSR05Gm+HR/RJqW/fFilV11kQtBOK
e+L8mmBEeH4qHhTaTPpWzDk6/VrFcwMMZTyAGo7EGxO11oqxcxXuW1/ubjqsKdf0kGXlQvCx9yrA
uij346jYta05HSzHkzZ3hv25YY1OubxN5reTMAFxOHlyePXU+ldzSjZyBOYSasdAFuElsYea76so
kox7k+ELfN/A7vJQn3sMN4WT2rEjhBPDCOJVTzbtyUIOtrsQ6g8JwnNY8Q+gGaJqI99hYLo2xIKz
97OQCqLtXQjtQ8zLlIGy1KEfKAzK4rws8oqS/1Zq1SuM9zgoS/fiFB2wZ0YEIQ1VMdfTz7Eyi7NC
xl1Ko0+CP8Gd9mvEK2ZH7uwCsZ6TNnXaRiQwKiTS7nYlRw1ZvXyhgrl1MvveojbHelGvwi6qO1B9
ZP9wo5scvSXlHeeRMteBSMXfmYggGPrSxipVvE5dwjMxWOlcr87G9UGeFh9BKwzAwDg+8nrJYB5E
jnozLFHtZeuU7vadGZvUf80Rcjvi2I0+9LzkYlPyTdpC29Jqw5yuCiIFEIzXno9wi6xf4AXT63is
MKBnkMWgFcN+SffQrmr/Wc2ZhufG6dcjH7H5HMF9dvlr8XLvi0tTIReKL+BdsUKj6bo4WpfwnHEK
i+6ry1s9lMgv3BxaRfLiUBGNHGsK4doVkE5Q3auAAmVGAI0DBsm+1AC9gJy01IsWpvuOwusPUfw1
GfrpxAqSrSDz7QmJc/coAL1qPSUfFgvZH/cQfHM98kvQEEj+/bcI/rFNEy7fJeMF2K7wL5pnAwib
mA3/13lIVgXvoxREllAuWopTcqvI82liLMPv1O7XDqp98qN1RTJknEp/vSpUeXCn9vDK4NC14rqg
LN2T5HsV4KSL9wL2IX5F5L6FSYBQDoRaJo3R6nXcxqCOz/MUJ0kc5BRreQhsQoJHlGWTCEtfynZp
91VJYEx/oONIu7tEd0hRRz5hc3j101Ap6ndhVNp/3L7UVYiYEWctQAZtIjCRPB9PyMW86Bm6UDJS
BICdDxfe/VM88PpDjNVa+nEVCz/NlvV904ht6Tmk9iUYPh6kufW22tlw7AYKDPKFsniwa1LPZnDa
+pol+GurSiAPUDCFJCZ6v+A2OLChT82yGGsMf5P/AajVCYSAkCQTJqsLEkN5mHL9FKonwy5D5vzZ
atIN3CBDo0LEQVg3sqhKCLai+XxdCXsNbnv8Yow1lInHnPGhXNPyFLtzMmxJ74vW85r3lu9GvxTO
eQnVFa2IKwdGrwx5G40D3HNfy79vpatho1ozE7n44cE7i/+CAvlLdVdi2CtspEGMJ8G3RONFjHNo
5exVM+dPhU8XQzF9VdVfAkbnAF1YsBsBP2mLYcWey+qMdtqJdzobCEefx7xfq5rBLLMPq5Tg+ny8
bJQq3lGK5sdkMMCfI9m+uFl/3cYhcdFNHmMkg/gPHL9n2XU2o7GeZILcIkFuIZU7gtW4UBKaTPLJ
0OVQ/5/Tz3G8tohfUelGa1mKd9ShxOQ7fMzdML/MuEQirTAXk7G5CYjpm8UkQNKV3Ym5bYdNvER1
7fzY4Zt2znqr+W3LuCtNbAxW5Tg/tGF0qJlNWNjzOMOswFgYE6weZdXqZcQtdB2AjmG9Iao5YaCV
5zdPbuXbUkhkhFBozU9MJOTq6wA2iqvO31B5oaGJoB7CB3G+aSMa8T6rBIMDj4UoFfKWz0+yGG0E
vSkoB/GdFt3+TkqskDQ5wHL+TbFAUInlar7T6rozdYoXrn6seNwEA/KcVCxe9/xPHSSu7stg+8Zc
pFzffjT26qmVkbYJ8KMKqwWfYHg1HFThO2wjLftpwXdx9aQtuyfa59Yb5sdcrogqFZH3F+7v0dkd
jm2xx8trCxaAikx3//ThkYyk4nNh591WUnoUeTlV3EsOxwKqxpupP4mNjtwIBfwugOQitBrQGi6P
uFS0XaZEDHKrNV1J7J2ijOb5n8SVNPD0Kw2F+I9CNn1ouEuegid5d2y0+xRH8YwbExizgtif/jH6
51Xz4wBerx45NHxsKk2u3jvsmvg2Nl70paCvSyxwFoycrd6mlF/tOAoH5giLfH+AodKI0TtJ/ICn
A9SDoa1/Q3OAzNDTbsgcKiS685sg99bf2mf+rslovxa+XCBmbrKBx39qTF73zwncpOCkPBq6VTEo
608AAzRewZOlSYzCsHq8HBnHh8ZmrdIdGrljXIizt+6eNQSi4B4CofezK8prK3WqdBAsXCFwzdvq
Jb3+DRodV3gtCUkDZCPf6lxq0SuB0eySJPuJI7LCtp13q/kydQUxEx25a9hCxfgd5gRYT5L3rQ61
NegZKLIff0zhJ1z74Bk+FUNP5Sy119EN1FKvnDU0VJjDmJ2s0F61/d7H1XqVevt6mNLkbugo9BsG
kyEufU+koYAuXg9uRoESEivnd0HZIp8CTQzWdk9e3Rpru1zk1IWF7GDr9KEZpf476OMMen5z6dr1
gCQguO5DOlcBpDAGaIMpI+KCVi3HySQrIPyIr7TO8qP7coZAy9wNqmL+Pl2VAuJ6lsnDKLp9GPdE
1lmLHqOFTsm0OPZJsL6wQdG2oeB/VjJT9I+uxpDcqNDJCypVBtI=
`protect end_protected
