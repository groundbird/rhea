`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Q5VtxaZ7x+67gumd7w1hJk5K+v1u3dnw2Mv8Pr+CuTjw4wvmzBA/El6il50AzfmEeOjfqil1Aaqo
VyLP+Ligwg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F8pCNBi8VU90gIFSHWBIQXe5QffySfqMtCSDkF4kQokrVP4TGXtSNDRw+2IQHMkjkFZces4X4hjr
7AFbM9cUO3a3demvh4Q/KSoOzr9cIyyPNeOIRCJ+MhP08hqxsffldMUZzfwNJhtsXiTmuVYfaVkY
j7X78dqS74tpGsMpYzc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AmetBhyP9Mk4dMMHeGgpcxMlUr3cOZdeu7ZMly6iix99Ij9bzxRdYgNV89ndVK0fiGU6ThkdJsaR
tcwQPZp8ZJ+u1CFcdABfZxeA21NFHwaSsu7OPC1GJsorv+iX797RLwk3cZKTqIduIsiI5Lns/zLv
YkegPjSYqSbcoY/3n5FjXyr0jZx+SS0L9FPulL7DQIerzebTfMzCNu4hSdzSv2g37z1m1PnEJH0i
A9aXlVwyXGxokbkVcMIhcR+Xh1Of9ABUzeEr7IIF6KyWCLLzGK6Ot23p1/EBb+eGrddaBivAN+vi
m2zYhTZCcap1wF9cnCUv6Z5rwpDiSfj8OvVEsQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RObJWenWkU1dBg0RvZbXykmzEao5a4IWyxHig2HdkxB07VeqxGGAoTsZQn0qiRKigyvzCKWRo/p4
5JVbxOzw9FXnkzFfIKc5ZaJLHhcPKz09vSITf3oCHxJoHUv7SmNArnLtdlI2AS8VIaFTgWyOk6k6
uv2GVmcn145sfnjAs8M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tXjJcEGUPH8T8tOjn3zLpzKi901VLzA8059Vk8++7OWYHam/3sPiRjwGXKiSvnL/PTFL5Un6HCLL
aL3hXd8uWOwW3ng5/lG3fjTMhHDJHGYaxrB2/53Ul2cjJ3PoZ1lLXnbY0ad2LljnFikmZavKYrdp
YHtiJAJWhMPO8slFVpFUOySKlpttDbAhaNfT3/v+OVfy3N0CIIx8lNdhwPDJtXhjI28I7sAgZc8d
r/DlrZyPRH8UVLho256cbM19dP1me7SxK7Q2RtsKmKmdVBjgUiaLQkPCKaUojmFCvl+kxVm2tADC
sh9yQ3u3SbuR2YwtjJS7VwnClCyVz8Qo5Hi4Yw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16336)
`protect data_block
liw5otRmDyY/4I/DNVjh65qP18UOqstKtoLQeyA5WrjYIpwYeaGtwdOTWkzjmodsoHcn2JxQGGWV
421Q1yyDw7iX9wZGOrciLq6BJMXEym3ZitI0bT2HFSk4zpjRsv8bb0+gpAtN7u2axTgDZ3CN4HWa
/TRTe2snrV6vJf+en8Tbo+gVVDQtTYC7fShjFZ7ZvjiT2+J+RMIe/8nQx9vOoUNojQcbdXycS5N5
qBRLcdo7ZrZxtsuDv9ME3KTzZ+xNYz8E3F3bcTC75FEnqahPoeVJPSUEhubWOvsd1fpHnl1Xj3op
8bZurwBfXjl8DL1+vBmiFe0wFrmgIIDwoKmVx4FchcnBve/TS7ltnWkblw/kmT/UcDT/AC75ad5/
wLgSgD3785cj24uBGGqn1KGoW5znaTkTdSeUyCjMprjkPTuzo6adoXTE5o6fxzZTu8lwaBGrVI4M
Cu2U1d/4LRePnV9BlziIkIqqsOxhWNTEsp8gBPNvZ6L7nOMY73eZeqAFqzGhwbZhGOXDoXjzA5qI
Rt0k2t4J+zmj7ouSWQf4LSdkPKqAZwxa8QQR6mswXB0Ea7X0hGAo9Aqw4fVKOfFwM9ZkPV1u2Rur
xmo3RHqTiIrEfm1xfnBTYE7Cgnt0X1tjhKavnF6V6R+ocz+T8b4BGpS1ieZpsZxmWS7bjkaGExDX
p+OSCOw2awEIvtC7wx4RQhHqVizPCZ+JThbV/V9EjM7xVcPuwcL21W1SXZUHdCCLSsyPiL459cNJ
EUrnx82eszqVZpC2JWShaXu7kxWqFiJgj7ewVvZSOUMjWfbOEEnt05LlurRpKIbo48kqrHEYWcbh
b0mPG07IfZb3hNT3Mj5iMS/3GR5d16vYxAQcV4ou6WbM4yL5YTTI1VTV3EOm5r64w6H+Rf458g4E
dmhzpAJl/4USupFcBfE4CUGKr6n0zfQYqAiDfsvb4XD3RQQHhSatNEPwAj7F8E651i0Yn7CjQLOU
fxZ6TynlZ2d3vC8SHrgUNS03sDK4BDnr+IbNDG0QuKw/VzEK4uH+VH1KtT0CaTZB+0wI32xuL+h5
RpbNwL+oEYYdECKwpy/Py7pdjkbP0KR1a3+dgyMzjHjoLdBeIY6gb9ESaOM9L4U5WaPJzB7Ld1VI
I6xHsFTeU9AXq+W5phxbxS9IzbIU++FwSE789NU8NzBlQ0JGcxPOoN8sJ5JjiVCa9Fkp9TQPYj92
n6U17/akCD5WjnnPOTso+jWW4bctkFLS+ab2Dg0i6afPh5OY80mRnDFi1aViFrr88EHlAnXy3VY8
mAzlG6lPA7rPBUbUJuvDkbW+qdYcxm+dOjHhbcfHdBlIu/2ZWIrtd42UhQi53ChR3ZJvt5h4JnqP
dPwaFAZkLKaqn38hYSm9B8RaoxpNiNJ8hvksciLysWfxZuVyTcYEo0yiin2BEXT3pUFZebotLLth
6wRacyG8iBKgMEVyWBLj+KHDY+h1lpcbARBIvfPOlpbOXyzGve6kL5ozjxsvzQpsuhr8EdH32G0M
wX+1VxwZxMYkeLRTxRetbFkcijIVIjr8DQ49ObqIuKFkk3kFrfx3guKnI6X23O4BzpaLJqKCEK4j
8WcIeSBho4AHLPuz+WBi/0HbK9F2Gq30jKH65o7xP7obQwy61m0egvtePmKEiv6qnKCGzMOxqo9e
U3U72LzZjqCr5Qlp9CbNA6WrOh6JN360xH5j93TZjAc3K8HbNz597aMWm3jpDbTcL7Hx6GjsHhz1
1juh/In1s3u1x0Tck+CFxoOCuSneXGV5qUOSWOaBAwYHghsUKtX4oxPyyx106QX/oFu0f6S/KlqX
ZyqCTFmZPSk1RwXk/CtXqB2jXq3KA2wcDRS2x78UVbSlU4256GhhPQZQEN2DljE2ekSJxZTqT09T
beQZoA9TEqrbNN4nO1uyhMvQQxYAYxh/O8eVu5EEWlhvZBBPkoUUGguQLwosFiRBiZR7ydHnXaK8
ZksjFAfcQUZMIBtgW8n7BANBDS0IWIFC5F0d+bpYWdAPKHQoDEaYzN9yqs66qK07lq6vHVXGsrvr
bvAza9t/yqb4tRzl0Kkkx68aoNGisI5ooz5F7lnhXUcd7DVm2Q8HlGH2k8pjMqSsERKjlL+Nbbcw
b+rK/PNucqbQkFGL0DB7EExWsUV6JlMYAGWbtrF2/5spOwqmbcQsgeLdKRULtp8PeeVACAeodUV7
NPZYFTyxrC17Y5aSfyzV7sCqS2lI/bMrmdFxe7lu0UUYeuaUvKUBXO8lFMxujYOgJMcK/6rEnhfJ
pmV3hQ+6qpg1OEsztcXduIH19HLNFRZEg0YGdboX1n5lGJ1tCsFy0bPUEQDvaueKX2fgqUBWBegB
k7LDp1SrZWnLOjlImbkPgWLk0I4pHR74Cz4KDGOBAY0VBhU/QKY0bltWZMEuXzggrtsglJbvICkb
20lcxcD/2s4+5h3KI5jcf7m4TcEmFu6Ec93fkLNezOAzDqfaOldTMzz7i884NfmNt9Q7Cx8/WLwt
5SMNtiIKdQw2KQqX/fY3D/jJsygTTXMpknLdbrb75awUJVj8TLiuH7+oT6ObtNIYkd1EDEpFiffv
SrdIafNfMIoXyXnz21PIdn1joUxssZ4qoGxR/cIruM/WDnaHXvpqEpmd3J/TjA0MCk+wLUpSCq9Y
8FrktLPZE7vgLUJPOpGQjHWlTCRwDUFXCI11zuX6ky9ci2QZpXZUKJ/2mZtRtHT9UegbH4OUSy5C
v0NoEpFSUF++wZLZ1UkF4lD4BGoAC7LDSfKnLpZFZiv4tZM4ZGpu8sAKkMoJYmg8CzVwkDbZX96Z
KefL36ikkEV5BpK5YFG98O3ctV50tbjag1G9S00SYgiM8X7foO/0iGe1xCM6yfhns64aaVus0Lkz
w+OugLRg5bCcjJCBjYgBhJBPHbwQv/E9kyGz9UnNymN4aHpUPtEOovOwZpcVmPwT6KUS4/vkCtYE
tfYaGXCLxDOJgYZQaueSzbJXTXZDK0xvkb8b5ObIoV42ehbiMpxA4Dt03Lir4RBBxOs3HvT1+xK3
BaoBvwWheSmABcfLUEkKXDX4msgNO+8QHrzs9AqGULTcbx90otSUvq5xys9sZwnj68AgoRDuKkJI
WV2Qmr0DbD3tR/z+Ctaagd1T1p9mAl64QcZiUW0/GyQ1AD98S1NPlwW3MYBWIWHO77pSm9cCj6kK
3YntW9v51nY+u7seJZBC+usy7Fca0QUJIa8h12ws56W81OkUFBFk6/T9r1Vde8kaH4VG7B9TXLsg
IJoTvyUagIVLGNnyfA/IUa6xyYi1cHBrUo5m6uRHzGlPcmZVm/qDpgEl49FWmEYm7NpSmAFaWiLU
It8V20/EpDCwN4hSHtg8dyNYQWfdzu4ynnLrHOD1A7krTLETe0MH6t0NFKPbGpNxKREsZPJ9tLV2
XLW9RMge8J7Rbhe6Iu51KLLzQ8AY8jnawPdt1XStZ9QgsANRzAIiOhFXlG5evkEtgynfMVAIMtH2
iBuysRayq2MYK5+F9glLqX1+7dLWGmmcrgzXEpKxXh2lwkc9t2aE03/DDYPOAD7CnsxDdaBB3/BH
q5cXbTaZIo4H2Loltt28wTMXl3YD4Mqcp0crQrdowlmc1KttRCBpqLGESWt3vG5NIrBW1TvJgq5H
YwR+LGWoxVM/4Aj8IV8ykItKmB3cQ7Y+y7Wd+YzsogEOldb36fJCcC5vKETNG9A/pwKOX97lqzXC
dO4t07TDw3dEjImMRvEXoOKc0W6IZDMVFVIt9yeowfzE785vLjfovWcwk9/NTmlPMAAQIgex18zi
wpM8TAqs53fJAqLry3Iq9tb3gFJHzC7RfWpYjdKcRWsw/nkdcnGohf1EzMHgdantLCnWWOWLtVcr
lvoI0scD1oTsPA7Ix+jbLuN5kdFeN0o6Xvt04oT+uhXAAr6+SSCv9hxMqTdFuqf6T7Dt5XZ3sfwa
8Sg8vYFauWTrm6ZF0+afDMIclvg5VagaEFg8oTXvt3di/ZpUXXFYnBqAzujPMZ7vdXe07npmW6HB
CxFPimKdfV/KNAj5PgxA7dFvuFp2iBSsx76ndWbsHyAIhs9ZvkTuaTYKa6Bu8UOldcgvoXYtl5qa
Yo1g7BLLNpTT874+hp4ObQowVOM+vgjm2SkZ/PTB5laFm0AAQwIm3+cMw6VFNnUf5EIAz6eP2yoq
InkUJzqAbBeZqLPH0xhK2Uq4lcMz2o7KFwpSjQ8fqgiNcbxVOjE9Xb55STeDl2qP4dOsSpE4kU11
IXPP0JUWJTCss6vi5Ac7TMYLAhe2lMgOvhCkk7ng+N2Jwcw8rx2bX/crzOoUFTg/B1QvPyZD717p
HjwfjL3dZDkuR+z43EzBSmYo4T8ZO+hBSWUCZlgMJNOFimXXR2IfWMJdjf/0UBD/1F+tP7tX/Wcf
z/PzYTWRxPomo8NFj0qYgn7dEkfMOynoGw6nZvalpzBXMH5I/s7xyP+qXHSb9YzF5g9/B/oDTG7R
KJhEOuRh0PP/DhW2c788WYugB5W3i2MPS67Iu9EYRKLm3JMnnZiLhWSW+HePQcLPBwHIlytXtSCk
u19xyLvzrPwgXsoX1ag5BEroDFVFlWsCkOMiejvzTXWxzEl0fnSMlG6lPe4zLsnVeiERSQAgmCQp
89gFiNIGtSqeUVFZi5kmzPD7f3TVpqBzyeK7WO/JAX6+PE1+79cwm9xX3DUAO1ZsrA1H+26gry4f
TLc8mQRe6nrkGR32oPoDoEDxHZBkDZnbRD+/5YENw1gXFe6F5kcULK2nTjFLjsJleTDVQoVj+uSz
ULK9CbfO9R1wFoqe+O5aenI4nH6esfcItbuBYnY/wiYbBqhbzBf31RyKvlTl7jgR55GLAGK2XhuP
zbzS5emmtGCbBbOEPBIWgnD2Ys+ZGYbboqvHE5mxqlVsncrtUSbqogVYjN0mru5wPLKp0pJyLqP6
L3BNPY+pCC9hplrOKjKQRK60H+wzmSbSdWU+fDvhvFsrIydkl6BiLGx2RUYM/ftr2WVFTzkb7jyM
DLojr3dWlrvxEcC39PL4+bp/Go2aKDIBTPIE4+eXrBE7PzQQaSufZlko8B6L3rkZdp+P4eg2cRDs
7obYmuLBANQwoad/5Aby4YXKfdkzM0YOiPtIKQxjZ9STsT3QeyGOIcJ2wXViXzqxw2NwG9lczKP/
2RvaN8n5nMMJXHos775gcvI0R+9t3JByEVRvFefgI7EsOVa2JZFJP6RA5FJ54ec78jL096MSy7X5
f+7clReFI1GB5Vankt4+33ZaWVvnU6O3p81tFAF0dw4dpuqcTx6aMS/G4ymCgOTbcBakLHM0W/UD
YyLApnSMedIZyFAdAh2IJd1zXfmUHHgnWVpgIN6mkOJOYCaeat0icykMgkAR++aGFrgrW7IKQEQO
bjw0M3E8QWqekQfkrO+ULrTLLuDPJ9+Qs7EPTKz3ExLtFk+50THZ3n/7DnrdKCXlvzpoK5uPVzMi
3cuxGGaApZPf0U9aPT9E7L0Cmc1uboHfHBdrEb6A9zYUjIgGMG0amLqYL+76Ej4rwqQyzMtI4zLO
KjBP2TwqNrGMEB2RzJd04DrkJHL3WitY3K4gLewLwG6PYQf1tTwVSNS2XdRsBL3of88Qd8tSLQx5
bxBx/xvHkaCpvQo8EOMnRBzyLNwuISVHdlehGxrBb1dgWjmg2hha/dFh3J3ArJFJaJNTUizZc5Nu
gOPdxE20aCwGEpFlD+H0FWn3DdcDMoqza70MV1u3JHWGr8h5uwnFJakm+l8DyNg2OjXKlhEquDuR
Z9eMQXRyANSFGpMKbY6CqHfIti/wKARsEf6Ei/+KK2VF1BxUdnHdzmOTIk/DC8iKnprM3xXeH7js
KO4hjAZ7+eUO7JW+SlgJY762oY9XgxiKpCa025phNhDK2yzkv6hBq0NhrgIZv4F4i0iHMV4RUPpH
qqBkL8QkbOG3pjVIKnDGeHIBdTp4ryu8NxRI99n4JP4Xss6YG4l9DTwop72rJO17b93ciYZasi0m
Iq1MEDR+/t4iMKOIW8G9pdNR7tJYS0uD2TvQXWIjajQVuSi6nspVN7Qg30RzFpoehYAOOFvUKqFy
6+P+q5XSCgMZUZBHZAEQlvOPLygLRX3CjUus/BkQwJNvn2rahcPAbsyQbEUfuvjCW9YA5BzeTrs3
BDKuDnybboQFXJV7XTkZwqUkgBlIIFXG31+A3wF3wETWm0CTCv80voAXUhmW7mxZMblsdgMMRqFr
UghMrB8kqslaO1skyCP2Gl3r0vPJSwKZYN/XIioCoBKIo7YhNbuwmoN1CGjrO0BXSWmI+JZQu51f
ckxZMFH2ZSlcCyM8XjD/aJWqD+BtAnUgfxeBGcx0RLNk09O79cMkHETGqYCpS+OhsDf+2DSZMOWj
Z6VmalC+qbGXV7cMZ3KwlfANpTLcxpzc9L92q78t7YFqTzIqVPvGV0MJOtdUP329+b8kWMboIzLj
fEGgXqp1ICHHthxm8a3NNWQkGW0m7FzSourg9AH2KzfPymoX4pJAGoMQRIvtgVq1487VsVocyQEX
DPNyo/ZtSgWFK2mhXFF6uRB4KHV8ivnpNUfaand8mwOA0I2IY5qFJ7IwWVJUC6b8bbigFtbiR5zV
HRoqFk28gDi8SJjBi7QyI370nDPZRSu1uKFeku60f7uO4pnUMSVJTIAc1Y/tYTajO9KqMobO7ZrW
xmYnNObdr082Sd5N93C4bhFSDrIBGMBbmlvOvj0ZEkRQAT1ZHZ54U73Quhr6cMSpE+u2pxFPdE1A
dhWyk6edDR/4TNfu5oxeK7FuAMpKbVgKzE8SnqTTG6oGex8aFMMqvpgD41+qvokYs+B4kv2T061b
cjaqyuBYHzChxKWPDtQR1JkOYhcdiZcL83VLvd8x91o0y+OucD5WOzg6wiAdRPlSPuZUe4UnFiis
zf8fto28HGPpSvpCEOnknb0VvZ/lyWwMi1Yok/HeMgFG4w0UbqfHBmfr+sqMhpRZ065TZmioueIV
vVdEwMJQtomBy6kp5qDB2BhhPR9Nwfm7S+RT4oGV29U6GRqMw6W/CSOyKk/nTr8Gk/9H1eGPfGPc
E09oT4bUzqfHc+jx2FINF9ht3YKaSnD1eWO38BTBr5NloKRl3hZvlZkkq0sMqbJIqc9/dOO8FnOa
x1HnBO0hBCzQrHOjo6ioiuRbOhjyDHYRp/mxdIXr61dWLgFlb8Oppe6MeVUgTMgaCwseRmtu78+N
gNGoBnKGzo9FY3i23tvzCNdTiEQ6prAJHNfJay+YEg1ivy+5EynkdMueorM7p93Pvck6A6KAuC37
AHNcgve0PtJS2rHuBd9ynyN31d1mN69PbYTlfpHSoIWu9xqZrJF2YDiHokAbCQFpTiBBqpeDSj5C
/l3In94YVloA6ddN1BYF0f2I2Vci0B4Udn7vbD0CzGRTZSKOVZsho703NlEpHREaSlT0sSUW581O
62shqJ4S9tDHDDfyLiZ0Mo6qvMU3Djt6szaZp1bBQs+AH63eeaoo+gLox0082XjWT+02z5OoRhPD
Vedgkto8ptWWw4fgKjqJPFag7iLHipFGdiwEJDqbLTeZY9MMKHHhnzYf/i27shpKNJUFRFNKEN86
ZE8HDu5yNBdWUYIZfCRqHietWtOSqCnp6nZ19AbEUbwvBX2Uf9dtijwU+VInKnTaEoldMGuXdypP
B/KbmnRVs619wZfvbWl+HJZAMpn037+ke6SuKQTcX8thEmFg4rAMDNMdgAn3pRZPih4byLXb6Vsq
1w3/4nViEgSpzbOJdEFNdHAiLnmZQo2ftoU3jrJjoQHcQi4npTWSn9T1/cucRD+tZDtbJ1T7Pwmo
25CokGXt6zq3KUbGprx5SYdC31y1TVJ8+mrD5ztAzQp/WKT0QdBL/RoxljA5U6rgqIqHa5LoyHyK
vo6PJ214UaDx/uOkf0zYq1dol9avr4LrcCCJoW8nUAPC861FbDIKIV99gu00Vf4cYIs7vAQF1QSt
cfCtBW17j50LhtkjgopCOTcn7NIk2qg3CKYxLB9ouLQGqx0HWRAtuBI8b/80SnN64CQweEMZ0mFT
aGRrCDrmAwdQdRLUNcihSkt3/7wqEUzUUdVabIdXRuDCtFcnh1M2OSwg6ALPihfXnH8U3YVJ0bk7
lH3SPQuo0VTOlCH2C0m1rlU9ZiYfcv9tLe12LLAK710VQLOwO3bex8ZHBWcWmpMYY9DkwbAx7NQv
afFsehQQojrwoawpvX+05pKg5+sD5F7fT9V6L01q4dj3wP7jhb9qd/hWZeU+K2C7vAH3PFZTmYQP
5X2HyflA4Alimaw8d7vJ44N3E5xz1n47fsrs07yNF+SE3TTNS3voR/rLpCH9IEcxf37RU/Vj9RbL
mBnj5R2r+5bGD8Tu+Snx2sNop5WWHnhnMwZTldSl3oGgOzMFWcWVxnnTFadOBN5rZP5X2/P49Kiv
Uih6mzZGnUoJ+PTgxpoqtKwdaUvkHxkklkIprV3q3YRJktKEJZqaKXN1b+1qsEfE/uy1CdF9GOIT
+rby7FBGVBKIzuCS2o68TovRoHZyIg4GTQb19BNB+7MsT1ahEezpHNNBep51UsPBbjn17TYBtNbx
UHNsHUzNxYel6cbl3Jk1YgMWysNirDhPxqArPHIvWoiIRC1aBTw3L72YYnqzurNBssnZyYDM0sjo
78PzG/9qTTim2VBCTx7gvxMv1Z4q2atWZv8VPaOJye51i5EOSgS0xgTxl9EQxjk5PR+vXhdUvjnw
w3FSNnl9qk7LGZI2JhlVhjS9qL4nAuMTy5nd3FfxlD3Ak+2lbyH9Fr15XmrlwMG5zZVYCDjqJPKh
z3o1l4PAVHKaG3gHLcsDpXci4/JGImTZ7Mzl55euTCuTlI3VFLRv1+tEDtdhGjjKNn7i98JYuO5+
GKnMjx3YQQnlzGQBbANEPaf2eSqGy/phomayYYN/B7sKAUqUJj5RuwqqgiUcD1wG9qQ0pNU4WV7r
1yzyjaO/8YH1HsGPFdPw/9iwaaT1cv/YRCJG5Q12XczB8O4lWyKT0W7m6mnN352aRSczHMxeswuh
Wn+6yRFdQjaeUicqUcUxrzcXia71OpkR+NJ5ptydvb4Ug3dYUxmmWfeyZoPMPaGluRWnLf3v2V0q
E5OlG7dMPpZz3x+x2DeC3HPsTZQdHnFhs+ORbwrWfDIgkK8/5AgVHCj0xcRdFWEP8v0xNogG04Dc
Aw+lBE1gQHXQiS9mON2tn4i6mIKphb6sIacYpYyAoRihc1fhQ3BpZXJ9t/NEEwM6A7yX2XmYZE8X
LRJ7gcsX27XwsfMF94aAFVmipIWbSklwNRwMGXz+F4Or05xyZIQdRsaycZBpXj9I92e8z8BR0rVq
jfBUeySjta1nBg8a4120zs/XygrC2apEvs/9DXknSYlA+G9++/otZxgHgO4wDwVROmO3+C/3EH1c
rHqk7N7kJK9SL3CtlyITDDYdkjAGFISz9ZnImRHD1HsuLFIJt/YcI+dLK6UTqiR01DZRhTjygFQA
f0nAfGiR5jA8iC9BXW9m1KPedKOjR7EkppHOSsRO8oefT/w7faPNgFL3VKdIO7dLcUPUUQ9xJC+l
4SVgLNoEPSn+/Doka5KPaTBf4Yrv47Z8oQ65iDOuxbK7OrGjjascXiWGUoDje/6KCecAiVNxmRAW
qRJ+tfBFYLDnuAmMtjG8St+ud1YU7gwfdFMKvJVWa28NhbdoYLq5MR16dQW8tsa0lWj40qYS6jza
mgGfdQFEzsg709NhL5PzU2buiNF4zjpySNOCr3uQpgS8YY3wVJUeAaYRSD1Y0ZyWAQRCo9JCAEvI
bb59F5oCrE/fP7h4jXB9WDxSaCWd4WHtVv2B9vmaERffQuwK3kn3KyU+CXHD9aSENiqh5VN1FLCt
6MivQaBImp3qchM5+aIQ3gWYPHckDdW7Gw6YunEF0wVZk8Wqr01X73ZSsisazAhs77mCvk1IAiaQ
m7om5H/dK7Amj91pAvTrEQTgxYs4MoQ67F34CZ530WViFrN+OiqigxwIl7jdbN6kyxFcgNFuGstM
yUYdbgjb/Umq9n/mgtvKS2HMi1UIoyc1zUOS7xklSHnVYVXw4UZF1czWDkksc98Tc/cY6RD+rVpU
VbmjLcV9nfE47hmhpU2t+VRF5UTQWNlXiLKpy5GDNUT/C2bklZ4Olc2y+j8n2SyoOrvaVDYBULgG
x7KwU0CbLLcxoh6UUbFlXntZQ8ramOSxV5Vvz0rDNt9RCx510v7K9P1fgj9rj0H1XEsrpQHt10VZ
AqtnSM2fnz74RhZQOY9XSvDQK8yWulwgjhhdiAwvAx0Hzho6u6yUL7Aia5s+ng0NzoWHDUyaDnIb
gXDe0z5cqdU7RvXF9v9LNvXBf+941/4BokyBQNlZXc0LjBSsJCDqpeufgJvx7tdsz7DKV9rS9WzM
KhjchzMTMnOQeLf6DSSIrZ0fcXPGXWwXlg6533FYgzrj7jlICmkSCq3qxvWtS89a1TjEcMXcZ8cB
/xNHaFCdcFoa4WnzxIL3TH+Hr6EZ+JV3k/XRoazsSLGhI9vuqW6KRUvDCoBL/548FgFh1Itxbrmd
cShe0sVbf+D6UuZldx30BWtwGPMxTEqh218frtKgesjIIj9WY7dvypAZPI0LaQpFdspnhqJpK0vK
om7qIHcN+sOxHpNqdUH32C6qtIAIn9cfAa9mUM6zEhKAwrtBJvMLlxuEvasFX9YEnnnJFrc206MX
hEiC5wKwqCEZBNbHUY4rNXEE1+Hrjhsvtl6T5XY1Eu5iKA67CwUo/6d3M3MAax5cbEF6yQ5YUsMN
/JXI3YfC+qsvLHIkszpRNgDwq8RxRQD3l4kpRxs1SP/vVx1klFk9mH83o6m4lpNukItsNAARW8rl
jFJq4nKzLXH2taJNpbwy0uZFptXh+NLtWRp6t6Z3pEYprsCM6py7RXPaRC2657TlzoeW/phCIi8R
TyChpJYrxYtSYWtsNaEqWsD9sn2unLB/zJnL66qVNJGGlkMFZhgi/gK2OH9s4AvO4uGH75KgZJ0O
Za1m72oLwtLPH8yCOC56Gim8DmLDNuhcpILaa0MsbvremIASDEEH/lhC/xo5CejJQkeKkaCqUtkx
7LC8UK46AVprk3DwB6GE0CTOR3+f/COZOYWwowmLCmiMsjhhntXGRXdu0bl13sBwzmo85upz8lFR
TveEnxCLN9Eiwj74DUmt7FgkTQ0X5sKuWDS3n/egVq+0S83yKqXM/rG32VJBzCRLnS8Ekf6FuVyi
2pR71VYp2XrtQKAltzZxFtZ8cyNGPHkiz+JXtxev1rf+D9ar/wJXRoWq0oagLT7cUi88vY/MzdD3
EMP8ObOa3s7TxZuyOtnbO9XDH3XBr9W1tT/aWaKbXTKICfDIOZKMhsrf6qwC1x6k+9R0z6eI9Xf0
pKLon7UX6/GuhAbY/zZ58AY8/YG/0zjbUWZZ3SjBUW0uWXT8SnkwqWswbA1HBSP5M9g2LcKFoIa8
7IpjbC2qSSk/wBPYrgS8F8e1ht9Pp80BE7mhbBgjGDYp8NrXsSFtgmAfTNjL4n0AUx4o6UbN3TR3
w4utBcXtP0GrYqZw/GT7seg3HxXSdhuG8sXHTT6q4APJuS8daWO2oqDbTNmNT4ZlilP6U46YW6xZ
7LnE7nI9xymK2uUPFGAmY3u0DKZjzh9TilDS2XjHvpB+FV36acdT9pd3a+uNNoMQP0lYYLSnTVQa
qmeTpcKmUc0wbfY1517PEZ1d7okiIM0jaok0MnAD4lKVqzxb06fipu4B4QSm2piC/OQSKPdCYiE7
Nzo9X5KT42MUXnwuZupwbXGOYpkrjM3AaUcRSKhHMR/qxtxpH09Uo2etQ+hFnhGhoA/En2+qkdYN
e7f0hUpC6mWJcn4SyFoKGEFlmjBYPHqKhB8VKmTyT8vX9FArMjoZyNqvEF9goXpUMWXM4kERA44d
as1mW2xRIzrhtY1eQYG2Fo7yWIrPUnTSbm5MPYeoq6/dvK9ce4e1JkDOv0LVJqlXfXqIyrQKuD0m
iPfWEux7c/RmxssV7HZOQRwd4kc8MXYDrwhkxpipI+ujbqWZfJcLEH4P8y5HD7Treu78ALsCIBqz
Eegnii9uh+NNhLhnaW/R2JkD+ITX0wJfbZCLeXZXPj7HUC243oiTS/Lmbdg+dpEoJ200S0xhNMS9
BrvgbebgW4nFlHSawwraw1GtgHlT9zeLQIUg9LnIyRwVCqJ8J9odlbzN0ORHDqZJQ4xoXIaNAq3U
dXb57+g2TC+KWb6WPCgQw6X4THQjodXuHmuxhWu1K8mMP63K8tDHiQZDJNYVB5ivykwbg2JQEMeT
j2nFl8UFzPq4mgpvUT9vn88NbTvON1celxoJxR0o4n8PlAKfHqf9G7B2m1FqUbuXahEdrbCUGMFj
EbgWszKeGiT9xoLPiFfTxLOSzNV4hm168JZrOSWVFq9dweM9/no0pRCxXRFZvU/AoCoJYJNli5ps
gfrxwPNe5NJsiNiJFqmu/XDcMgF9mwRct40eddkvNxcEg8o+tqZt4cli0O57gEXTIQIwwaD7Ju20
6DeO/xhD8D9rRVHvr8DP2Ed3LLwj2MnBOl0slah5EqzgaWkpjgA4/sWpZdRXrGbgw7Id5VmdXjbd
EJ1PF45eM3fUwx4aQqQd7F5ZRTEOrhc8smyzvdR1mvGsZ9huUCkhtYKcz3vAKG7dRloIBg8RQGIu
jJTys3xWONHJ1Y2gjhPDks0GwC0lvOQVD2MiaRTiCkyN1G7ee9RMBaeJO3fPLiuvkPfxH4KkCoZF
pKwaX+lsguociJdz6WvRizCdzLi21sQT0nuFQBVuR0PFuaXrgDxc58QmONVo+F33S/43G8PNFobS
4wcreMkw9UzFL1p6Tp0eIkRwr0ww3KN/GldBmMthWb1gKHoUBTtw7kyZSeNQe6irh0g9CH7GZV0P
frTkNA9hGlSvDuA5GujvEhOso2oikYytQ2rUUEA5hb13aoAEmUe7teDOlYreb8c1tRtOaWcfANoW
xkoizO/rycGaO793UHpT8D/cmnpX9DAn158A6rdGm96OFwiz7Yo5E7+DViWyTxiTjwZbXwE8WHlU
WDeLm9eOO4SKSqfFxv9OhlSiwKoLl9Foddu+EqdcT7BTo8q4B0kHNKQObz1irjz4CUnCiOAF8/mC
AlUrTtskuwv1dzUC+l19F9Py3xB51iHyxwWEt8QOmWujIOUVD3uAAKDSL3g2hz3eZJz7CzB2cKVZ
ubpys4axE6CFG7cOoHxMILX06jltDHe5D9MQdexzU/xy5oE79QkAs77vN5cKHc8yszoZVQVMucBs
XIQqe5rdGQLh/QgKPzKHFCJ2TobktfgzymdPufCqFv/a6qL/bk6OJCn4tmKikHAhHkpab+kJJTI6
7zuceQIUiVE2WOJXqwwPpEDpYFQbmtCyBZkFITF6DdhDanF3fPHbB2Q3F4WSCU8vaPUoEfVBQa5h
tAQJQQ97s69JOgx/WHqdjP6ysSp0MZuZgbLOVnTeV1J0Z8LOwy/vlgLnRF170Y7l7DyQ5eV/36Wz
VFNxbQw86AJwaxRmb9DBZIjILNf5LkOHBkBAjgKaTj947sVlaGF8/0A8uw3+0IIOEylLKqvE+jLe
SH2TOElLTXGeZbQWnyJqiTAhHAKpA+bQTIVtA2XNSsAVfrGPSMtWsvMXnFqaziDPfvblDUNgY3zk
9Tp1wFiMS2u9jO6VNt61YhMzHuoV9oXCTF6bjVOKBkQQJbKPfYinB/xFUmO5rQ7byFSIrG1GVITc
NVmQB8UxyOR82AAq4zpCBf2WbIXgzLXoRyago2AmFtv3PnUei4lzo961NFdNAFlZdt1FI1uquiag
Y/PmqcgMkMZHtWRUluUrXXD/2h+IPOGU3ANS6+7lZ/ezjvBwbhF893ngoqCBJM10exRjOG+fWNKS
aqgpCBWSxdIqXAyhJPwJZvqoDX2DX42wXORlc8xB0i4z6XfcH17tQpC+vZt5qAxICWHbFO4Norvh
XiIrl7uSNCa37zbIIzpVhT9svKafnFEZOD38ogEcrpjgJg0cdI9nEISWzx12f2p7u/4n2f+jhFxz
qk/6dIHGbDVYy3DlsHche8xTWiSIRGVaWdqrABQW8BQobOMjsDwuC3GMaRZTaPWowRyKYoNi/Gtb
FEypX680FGalURcNqQIQ/sJEv+6VNVBJr1i8Vz+goDZKP9A0fVKts8ZBLezTRM5BMKyH0xjmifQx
q8ON9/WxsTvOePl6rJGFg7pnYkFRn4TXsUHdrII5Dr3/t76nCo2oz7uf4zmuMEyR1Vr1OMJrU+Rk
FRRQfyO52oh5hPg5XkEi3jXdohmOWS3yADH4ZuDBn4H0jSYAtG8pBJzDhiC5+dfqHzjosIHKNmku
B+ezjupnV5F0jlR2QGeW+tNLa69IDRiTkVmV87IJGUkiBQWhEVPqSAXo0Ol2n4TJ0fJzr69d5R0j
iItb3VqlPChuWkwBWN764w6U7iasDlDUKRZVsqt5j6UQRf+pkRG31Ch0Kbh/1iHTwrQyIGCh1cAK
WksnLb3tfIiMX4tQSA/AX5Wyz2BLo0ND52QRI112AlRACUBbXzdN2zpfv50DfUesDJf2J5mg2X2h
fOfQJflSnzev+MfROqn5sF3pNCk9MMqvJk7ANBUJifWTa/U3ZPkPGHP2xEV0Ic8HphUUj7JgktbM
59c4Wt/DhBX+C5waEAJB/EKyNB8lBIBHjk7d99qS9b0M1BLd8U/l6tYkolq9NhQaeqBwyn6EVbca
8nDCzWVqELw4HFTtbtLwWPup3x5RSCWDfsiAp0TkQ8hDyp2iEz1I5tAV87dp/+61XXy+vDoMhPYn
C7057mUTdUC1+7pOJcTI9aCBmHOKm/hu+79Q1tmmUXjxkB3QLWzjTxgnX7WavN9MoyufzUj7/Efh
7VwCU81H2fv/vaetbOp0uNEyNBnij7kmHmmT6bOW6Oe0+KZFZvUN2r7ji4TNX9rW19As/s4WZf2L
pAuXCdGOT6csChlJNViN+NPyXQRN/cHX9WEpNdh2IswcGpg82dwNNQbgEYbl4N9kU5owLHerGQbK
DR9SFw5hQKK6myj9FjXiLOs7k0lrTwfzz+goRHN1nPsHmJkD8ZrYZGH5Jb5Xa/0oQEzqbUR9n1zI
gWKTrv0Y0CMOrHAaTtGMIvz564dH6u0e02boWn8oBESN3S4jkHltx4+nSgOBlkBweNzk0r463TYP
tXvibjseNCOnzwIkgKXfVzBPI+hVSSGx8C712yJInCiR+F7PtaUpaA/WZusoEaOk0cHeVGVPgQK6
NbXO9x7MCOtH/x/BQrVZGVA0asRGxNvraYrUBUbrszH4+7+T6dhZwO46BGL7+PKC/7jWrZPMScd0
ZLgaDuRBzSfAXda/9nUE4i9iCvQWVrNPGfIdz4NoRs2nWWeeIfnebO+3YOoyvY4GQZcZL3aEeC1E
6n2Zb8F06TBI1KtgyUsJWV2zoji13wsazv6J/F/iYyMhbwKxkDtibHm70Rtb+zAiFb3X1ELkar3l
oWuI+yUGStHXbIzVaaCZZF5ke58LTRsUaSMuDYTOlKxEtNIwojelNgu/k2kvvKnqBKlwTWMbWB4o
qhUkGVDB/jONFFA/EiquDnQX5cU70OtVLwYfVBNTl6cLFttK9V+EaWY8m5348LqmEjc1YAvUKtSN
bK5U+kI5XjEPVl9HaJXu2DtNeXFT/hzyQA5KmuBmzgGrPOwGtsygjj4Gio+RzeZWxGCdaQvqkPQ+
8ASmm4TC6Fzc4T5ashnCJCkIQCmtX9pr2nKUQKuF5UZIQSyotsZqSVmZNg6lAd5q/SbfmFqI5/J6
1mr7P29hqhkDEWrzyz7qpEoYGKeWCZapisepFu3wrg36HKCw26bxSQyWiSeNFSofnt7u+aR13vAz
yiyByZfS5BDhOdtENQ3ZCfkFx4fuoUEIiuXf5okdYGe02qV3P4YiWk+9ECa/9fiqn9PSP2L4Rs9J
LEV69L/SlbolCb3XVvsgUnMHkLr+eh8WpPa1w3a2BOOwSBI1up+eaonact2cJ1qPB1JGcBQkYRkv
VSPn63hoSRYUwk+1J94+LpHKuG9b2mr0uMQgTJhzRXPTwAWx66ATH0HQKtWa5OhMp8yLA6zV2ObO
VvDtg6pZeA+0vYFbPjg1B+/FGHGvJv8tdqDhNGrRS/fyKJ1gBsrdD/DEih6VqT0cztr0t5VPd1e3
dmSn9ymZUhImhH7Ar5XtBVx8kbMQAAwDPPqI2fw6nJW82UMG/7xmZeCcdHXAXiX7avFdokyPYkPZ
Bni1NSUIhxhxd5lcaR15W7eNCZF9AnfHU/3gT9/a1bE5xcS1NdE4yVgE+VEchwx+FU9WblAklQIz
872UjC4fdlf32aCogBMD5icBj7fCCsBI8elih9UTcfMS8u8ivLm53N3l1bRO5xT2S5NZZ7FB15G3
ckL540WKRVI6I6AF1SWrOTaqoLDNQVwJpb6fhH6DtnhjEn7XynCsmZpQme9G2cq4XkSZYdmrJv4y
iG4Z0VftK0BGJPiS6i3MMNcf4VqERQoI+7eoSwj4a1qRG87erq7CHr2q730S463eB68DRpujIDpv
IMB4aTsTVu8zsf6h0bbtG9V2w4D6ufga1SaAjte/dHugV7O5jysNlGKP+Z68jA01XkRe5EuZJEb/
xcquAuQDQxTidlvNvRhbLAdcb5xJdJbKYkPGcTyhdakxPOGRfks8LaiGs4799VD4Kq6zjbrUyIoU
E9lxPmcfpKUOKoEXTj2AjA9lSG83SsstgYuRWgIn65Cw/CnwUkCZGi/KMQRAQ214hqFxCe1SQ6y2
4Gd6nNNkLEjA0HSjgLiztN06HYiFuhKpXPIJXNHfs8R6hGCwzljybS4qoME9//UGvGn9W6NgoWnP
z32SfTY/QSNmeeFUDI40tkxJit+0C2X55/LYKVsgKQvohZm0hFFoD9EUcv9yuInlybdHWUwV73PV
zjCf/4byq6V1FsLCTDE02/3Fr0E5MT92gfGjUuVe8g+verMxj0Bkb9mjwp4CxHsdUW+N2mlR51ev
Ln8MxsGDcsrzqigqEqnn6IMB9KVk9sDpAtu22s1T7QZEKVQxetzSZr+xYpLVEPOh3h23oLDGjZ7+
ZrFqfn+A7Lu4hZR5SFEI88xLyYLoXO2+ApIVQaKnctP4WwQQ75YynQ23ZNc77efr9wE1UtdGNSnH
qznXMoLelKp2ZVf1FVrvRp5mvJfqO2NPnV1vY+LNqF3rWm2vYHKeie6Nnthci97GR2w3pVY0eTco
a533lz+qdoNztlLbZq+x4hjiWO98F7syFL7iwiHmANqzrdyoMtIWD2Q92OBFbI0JJNOHU4UViSpE
3V0RUvZVzzKBoP8RzQD+sYNckmcNUfDXkACmMiLUnw23StpcPk88BYJQL2k5n86z1Zr6df6LXSxP
PbRQlUpJ9VLPp7W/we6Hb/+M29LK2w+L7z4dRor1oG+AZtxg47zLznJpByMAk6n9E3g+hYEoL54O
OlSch2dqe3saHJyrZ41ieLq1IpjLPZbn5uvtPACllIoqoVshIxlpvFclL5rCVuJE8Bd3peg4tXR9
hk8jVPwt1y8L41oOUUtkBCMpeK9LeIMjZLqTGIzEGMa9gvNTWE4ZesJQ4gE1Gb0th4+mWn3BAqEN
b/fquGuD6bLsxYs8dBkhE0J+nF/MZKdFoKEtKfFF/hIkQk5hUqGjxSqLQgQpg746S0atW8WoaWZQ
PGZNoFNcKAxfIIfphF626Fa6WrRfkHC35LtsKqe/2Ed9KbabIEqlmLOK8HGgJitnwRK3fs90+gla
4LGnd3SaGx0ZoiVaMI+vGfm98jfNyg+PZVg/U3r/7M45OSdkIIYttopw+dwopdzSx8qsKD7Z9Aeh
iAfyHNfsOjnjR3j4qiTW9VKnf1Q7cQBgiRsYTKC96FfaqjxpItbUez+pyZnaesQJ5J9wL/gfBUrp
B9+DljyBKK3JA/zX+VSHro1tcOTPt7BIr1BZ8WaDFDnB8K70wDODtwHU3N3AGdMoBZAnstdqz8Vu
w6gzpmg/joL/0+WgdS7luHg9gg+bmxTjUliuoLWAoZde88vo7AzhfIqw9wmnEvcfTc1TbDTvMzfo
+D44DY8xAQGoc7leLl/NspWpy6io4GMRhz1QkUaeRIg5naYHqCvd0LSMXDhCLQndJ9A4944ByzMN
w1L/UCiVRpmmX+rIHPPZoWazQM0sFoIWyYHmR9zmY2EU+luD1msprO9lrhBFhylxy/xUqAzAVzWb
akIkpkmPSCZvlkimK4MGkL9y/2SemdaC9mSAfM/JYkO0JmE5vkcKntUxPRKgZP9p1XtSrcbQl6Tk
ugU4zZylL1t6e6/U5tiLpSAJfvbmbhe6H4O7yZQ9PnVYfHmB7jt7XjvjdeBrLtxZQrICg9N5eJja
iD18qeCfdXwuoIdzjQzuvAtObzcVfHHUi28HhNhxbwo/UkiAA9/Z3GY5SKA/JMZqkYMyB7xsR5N0
0xhKqnVG7QqQaln8vohvqhdbPZDecZ2mOgqax1GwHjtEh2ha2RXV7weFlJgCZvEl16b3IhVAXxVS
+MpMg0jl4o0IOesDR8FrVriPAAepT1j3WxavKTFOjvs7gDvNhLCX2j5HTU9H0dp+2moNvUNljgBG
EDB1+aYGDZDpyg+DFFAbMaJ0+zVWUASqMUYsqc9wIm7Ym6wcEN4N65S3Yp9GwhHSUve01tZ6q8dW
Y1e0AE/8T9O6Dmo/GvdY42Cs2gNdFHTUMn1qqnxdlXpGminJDcBNqAWEiYiahSMmLfwae4VYFVfv
AFaPGjbj5k2aprYigdv1qM+yunGdswHfAz3ps+0sqFUHtfFHDaj/AgFn11fNpNYjsY3s/7/gz0Yr
3mJedB5sZ2t6qIAWGHPY5b7xixu2VzFkFlr004uBQKN5oz+mUwsl/TTQEAaOpNgz7jIJpDdexAoE
RxiW2mTcEzEje0+x0vydvAaKOmC80oJ+pai+uMay8snEQBMw9XPBssWmjqfuDoCK93Tz7DWF3ccz
R9xyA7X4Mn/j6Od4Kg1sEBbjh/wLGHVtK5nBhdnoQ+Y/hM7vaYbnfSdrBPWq3zjvk6odGYclYj+D
HwZBQsokCmQP7q204nrpb5xP5mLGOU0FbrF66+mOpoOQ4gsXS3i0bd8IDdgH1j1YojSscoyJafdv
z9lPJoUNYicFVClVIxUaaoeqCjSfq82DMhL0BxxXDOApEqx2M4eY6qS806m/XlsKK85foO9PCDaB
jVRcUZj2ivgRKkkUb6ih41iW7QsRdsucBzybc7l3/dEO+lLuCm2Ct+xvs5FfRAOMcTQoZaojFtCJ
o0JgoJVVo37guhIF1n9r1aIlNZ48yqjeITyCzGUhzBglvSGkaEViPeqXGQ8uBRBSdOqdqz0+W7lt
FnlZoxPsJO1QZkdTD4SbGipxP29qhkvay71MwiodX0fQmoiAyUJ/6EVbWr4zeHMX3m4RpOv9h8a0
dbw9+0Km4nfikC886BNgyOgwAlNxTtIbZut4vXwAu9RZA0ydTthH+e6xiDz5pQWBRVCm1eNxSP7G
G7YkVTqFIlw8TCokir0Jxv2C9iHoRwYmj94DIQWBPr+FbWcPAcb/cPhaWMSFtzjcKsCET3/RtkvO
rjgLgYU4E7zIWtYKLVknhfbahMw57f/y9A1MwNooPPkyZBgvq9b7fIJrD9JrJWD0yVsX5GJbhSPI
Nbe5qS0KgwTCpQu6NW8Yt8+8xI4cArrYVe6EsjCJ+iRAUXgdnGScYbeQ7wCrX9uuFKotsRHMBRGV
2MO49BzPThfongryaZEfTpyyAi7DtKHK4fKITU/MdNKDwwox1V0JIptmHTo9n2CjQkMPhwFzC8Sd
zoEcHdX0MAbsII529G/7HXoYuVbDqJcdjOVlwLRdRZlkaLDewiPeDc27B/kh6dUWqV3S7MoJwn7x
UxmYAtqKA+aEcCmT7ILQEjLS7XrJGoKie8GVmVqxosZFVKzQ0VSEQarGmYfLkdXLpm8tW2MmkFOA
quzo0I1tfHAqWO96oH5SCC6ELH0dcV7AjTG08y/FUbcxLq8UM5s+3zlmF5NPX9IZglkubzFKqZDa
t2EHvgX/aI68OURupvZxvco2F58dapE840DTFrRvwb82fUmu/3JgJO6lgBE+09vDWZpYe5vhIQgw
LF4sYYIIF9TPdkfOwXS2vXr5bomhNljaazXw4ySIHNzb1rsEXRy0z85Pg72i3daD+n/MdbFZmo2q
lOp/e1xpS9pVBJUA6GOYWS6buUP/Sy7MzmzYiI2NeuAcn7Cw94icp+rWDcGrFUsjsKfQqGYI1Q5U
vgkPE2vz1gjUtH3apUdDNglTXKW+VqIns7NL7ivIYRIuxXzmj3CoE36A/6HQlx14j7D8SZ62mqM0
7pRD2cwvBSzOhlzd6FjL8JDoqTR7fwnSkBtSQJ5Kr6vV09sf0s5zVpVoDmTa4jdyaYKQWg0jlQNy
1lw02ZKHApedYqX09OReEWKyjFYTOjEeqvfHgJ5Gu2kSsISc+Ol+dNlCIKhZmbBJWyuDi7bidO3x
Y1R/VKv/5EaORrm+GsQ6ye/OMsGcy/Jvr9cXjI6Is2HtDLQVmahuopDQJZCFSB4aeiRXOzjcqp6p
+ko/Qpr2ldAUM984sbJr5f49hT+HK/2oKUckPsfio7MuH5xdgu59x0Qwfe93bXLiESsmTRwVyu3v
0YUZoJVV/FXAEq/+an3OX/5P22RXDo/LUpDOWHKJy/ubilOAY+Min2STPuEJA+9pWThq5jE7bsO9
DADFD3wHl7lqmnC5A/q9z3GlZGx9JYSwnJLJU1pgnyGe/LlCxYT5XIzp+jWcc2rwig8tweTNStF+
q8bFfSpi+BKZCkr+kbDAdPVm0eeKkDr9pezx0nXwuIBwrEXknADHuHfiEv53hfJIjfe70UZ6t/Gx
edVlmM7n2FQbJKRR+cQ7hRgSvKrLN2z4tgwtIELrA4xmjZOj/uNSwR50qb09y56GSAhXipL4w8rO
+wimR+9zGB5EPkazDD1tdU8mrMWG850gO6Pp6/y8rjS2Xqc2KK3hfrzo8z/1EpRUpK6rKRszcAMG
weon1rGmZPiByys3UgBpvHX+xKO6Q1oJDWOc3xzKxTXGOPLIfKgQtnePpvpY8JHofWxBi18Cdelv
2oDTigbnAllsk3L/JEgfcg6j9eDo4I2P6aH7Vhdmmi56TZq00HstOwWRkq16gNSEvKkUY90lopJZ
sVeZZwvtAvYkq2+HmcCusPLq8RsgJHX+hkw9BCsxQqiID7IEzh+cGyyFKtKLJJIBG7MoFC0oOc0U
6G4AFOt4FjAgTvvZmz6maVVzOfy7fPbHAy21bMxuHMbEmGVp7qchnORceEK19FDwD3Y9Oosbn7av
Hhb+vDA8Y3na2wKtNNNZcTpBErA/Qgzu44ZvmZRGmxtpeftnzMTfpzlifICsbJOl9GBazdQ0dLew
yTXz3euy9e1qLm7AEj2WxyN+eZa2WxhhcWpXp8yjFofS7Z0U88kikUEZfBmjHeQ0XUbV1GH/4zH2
4j2JVVE/4XOStKVpFdpF7FLA0kaFNEl1El3d3D1ZntAHb6jJvAZtzngGIGCaCXkTPyQKFF1eXl/g
HbQ9olAKb/iESNO1cfFKtJ3C5RrrVYQx2MAAmy9xZGNs9tL1SwF+VJesoQfLWrrxVY3+M7J099H9
LgeAR00GwoFQzkyMMXhsaMuz69jEq/Bs4fF7aZDe3R3kRf7xLkHFDTu+eMS1Y1+681NCF7tU8uBf
iuc8rrpvCamn2j+Y/am5hz8VSlb68npGgYsyngK09/Kkkg==
`protect end_protected
