`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OGSt9kblZ9pH4yeXTZqFdUUjbkWMeXE1xzP6oE35JBV/rPpF9h4FUOD2xImtG1VL9HbpcaynL7e/
uR+fxedJdQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VnIHGfs7MtrCwsgP0SSHx+EdyLB3fpp3w0L9sTEfrKUUt8Z+gergcFAnPQDaLSg9EuaK47NRySgT
rVZEpefoF6zN/GlMk6MCd7WRBfoOaajswUtbm1DPKNnycnrTvIkJ69HJiZIsATBNzW4hydOUZQXJ
hQfQ8IEAika57B04NUs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GZSrufdtATcvMzNU0yK/fs6YNXJoa3aPn0V1jPSJ/7OMqFy4dnfsGS42i28Ou3JCAnWa/lmsNThy
AEFAHpGoA0BZCbdB5LK03+RdjZ6g2yd2kLr0Ms/72H22bRXDvrJIeRH3A+h5U57CdeuWdvzZKH0j
iTHtTZ/sJ95ZCD8TpDKNzWUQGAmNDealu7GUgAXO0kK9+AEmEBdiaN9wTnuaD1ZPuaDnNa7wXuEv
hVNVV19NQGpE6j0HWcRu03NZEHEEToVx6fg8wHsstyttB06QJywg9AM9I7pjQRgjZR4R5pX8sHx1
SyHyuW14GYWF9lOtrPBM4pciZiIMQmzG8ZnFnQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CNms9J6890AYhpBzMRDf+uQlf6RlKxq1MXGcWfHStSn6uKP1bNqzZdSyR/hBy1TI9xcwjUxD2bHu
1dFGc35deQ2nQ4DjPuH1v9C9Rd6mS01mO5nRsTBswfo7j7eO13tdbhibAOHJdzuFTyM5lfdJv0VP
AAgCt4kbqreZP+v8uis=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t3Ga7g/+2FOQvu9EAib4ZsLK+mIhGjyrM3anHccd7uYoKS0Wuc4p3+bg7flcYUJeYqZvDt97Lr6q
8lvwPQpiI623CRJV3hwCoJwLdMxb85Mw1FRj0wDK2qN9g7/9ApbEGX7FPqsC6UEijCfdvZQHGoFA
MAZIpVlhUroQ2IwEo/wvH+dHNKLmrIKQSh+Z4khw6k+j6kWwCr1Tu6+10HfVxO7tmS/u9605veHp
XY0o8Q8NYlr/86uGh+3hWwP83SSWsoqurK7RGE6GHXyEazh43ThJuIXAfT2SWz/R5jJGCzwIHwcl
vXcXet0UEH+gvacEEGLk1XNscWCI5LGwP+4d2w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4048)
`protect data_block
/oXjxcPJQ1S0E0wGEqYVYmGJBJSvv+6LNrE8M0TL4fsgWvIys0buVszjmTsrh6vStqHbBl49+Hl7
nlyqgykBOAGVi/MGTXjLH5TXXD1V7Odt1NJhkZQpNY9GFQVphDb0LGB4+eGIk2Ew88LlzJWyS+l+
PKRDLGjskhqguR8l2g1LcSb4oJsGObRoW9lOyi0yLQ+0+1xXlLPvgo5PLEx3A462o6lViVC2TP2H
3dwTEjIgrZkgy0T/VX2w/CxB09gfOvnsAmvdjPR4Y1clfn6KIwam+CieD4il8z5FJJB6A3frKsad
FhTqHVsGtRvWWjayYOoxWz6WPTpwK0+7vmyRyfq/Q4Acp8Y9zeIJnaMJ0vkgjPGyMcT7whw7FsfN
0I8AqmROnZfNp5AjZkl5nJHBITJy1/DmvXuW9KgBtPQctNMetdTbRbZUmdAs12TLpSMXR2oeTUrT
KZYyLLCt8vtvgg2v6XpoFSODivCVVTdeOoewTUJ/mm99UhaH5wKG3cmKXFLQKGIxJ3YglahwikZv
5ItDbC+6Kiv+OgzZDisWjJzsJz/OgO+G1Zy4iLrWkwo0v3OiNeFcZ/H5Y6y0307Jz0Bslw30nPu3
lJineHWm0615DrRtXaK7thXDBVJ5b6bpxUn56e3tbJhQVSWN/TCw0VzJUis0zvqZTPHHpDsjXn18
c0wT/KIQMwoqzgHkDpS/arv5lgwOB08HQTkcFAdOA67kXCdb0h8BKpU0xbaZ81Yky866Mh3PrS3B
ipgK6re/Fro4+uJWf2I7yG0dbOa7Psc6BbgmBZEv4+3cGhTYyJdSKDl6zukx81jBtYoU2mNO1SZL
KUC3OAqg+Ea+piXx9BEGpGIs4MocUHdwv/HQ/Ol4LM1dcCy4rF4aB0tG7waX6QtxdETaDj3UrU+g
WBz+ths+Cln2/ilpW8ThCvkngVS3kBEQLFxCg34+Ankd+e4ancOkQEFzgQz/Ql7PqbATuQ1CRKKz
Naw04c9R9h0dqbpl44ZWp5VqHAQQpmgeEaIwdvuOlh/TvGHPRp35CH7NRabwAdh7a8uNdpfE/71C
ZVD4mTch6HXyaEib/6SxNFytS1nkALl+va352OPt6luTYkNeZ3lf2sabP6NPcRgcbMq8wurO11pl
/3U8Bvj78KgqlA9bKIlWsl/dWxXoXjdKsjrnWUZMVnGCdhtzBWi6kCJYHDijNVySIRZ9H2nX7nKX
QCcexYXq/1/9FPKbbdfH95/vMrKjMIgELPImAlgh4afi0mlzURdAUPfDz1/Xy9uKvzP6ktrmyBrn
bA7HKAucX6gUM3cs243Mc77j/ITQtoxrZmkBJFOXno4PhGUP5K6Ajri/BkUP3UNtBhJ7xKHO4b1d
8nZoDmSAovdCXOUoRurS3QnYUFjhQFWFOWbr99/Jabp0SJUoSarOp9aME9USw8MGw1K+4HGeJPvH
ocI0+QkLXiELmMiKFyriv6Yw9Sp2JpdmzMbd8bv8/3Q/QryLFG74+IY5SP5sLzVSqdIzeBkck/Wv
+84ku0pVYCPW441vlPvLhr0qL8WBR1Nw8/q4pbLb//wAk+lI0WdYdbirAYtEzZ2QxJOYsESafyj+
ozvC4Dt+0IzbSyCfyOJFGEfX817vBOTGwCcZPfTRtDxuDU+JkPBjArblMNEvhT5XWcqfBCtMenqd
r5cIN9KMN/JrvsQ0myJm0FSF0d0X0P2aWNcG6kcIS51f3NWbq6cFlD/c+kxUJP01wvfBVoSuibZn
hZ+p/rEI2H8xaMtwDy7BUYehXgd2BHJD6vfeq47LLr24pFQMAHmuzpRzJAIYqx+2UMZDZbWhRz8i
f1CgvbzDR1sDxttNG9cqix5stJrDB5cKULOEdpXQuZq8upSe2WRgHPD2pVb+ypNxJwZsHA2NRPQC
AtDjrfOrSXvHvi/3MacrL3MGSKf3ylxoUTcyTBTMYqZonl/M6q+WbWW3BOOPplOhPSyH/1DGNfs5
g+7BX4UfkGQZ7d+bJ2LZE6rmrV2DP06JHujGrw6AJh/XZJxXOqXvhDgJ0ZItkHdBeJ9E99Z/swTC
nxFAvZNHv5BXuTOW5678h2X43HzlDfNpBDmUVxIPErKpss+hpLEBpGXhkSvTzNo1bPYdLbqmUmTh
8xru+mbBvsqqIjp8+xMRHwRh7A6I72RMd2OBUstK10Zf0/LyIFLr7P38gXvjXxieXt7UA8pbDJZi
mqAfpUZkB8SibHvmbPCNadY7Zim9h6y7SLArtga58ecwR+4nDql1c/LfntJP5+ktQmPvEHGRML/W
WTf1H9mbzxPTc8wT1h49FY9z3uKBtk15q3915GQQeqXpDW4kG0Jqm1ASiNGv3Fx43uh9YiglQF1s
Rz9IT2ewx/JuGNyyXVp+6SIs1/MDdZKcV6hydU87AtqbNwEbGvNKLudndZMu5N6yeXKtaFkyYD9X
fwGLpyl8JRW9kvFYAVt8XwLQJR7wEWDDYwN5LvL6Qj56EGoR1kcE1u+rTbZDQjblf04TYs3pHwY4
Shovo66Fk57mu438Ch+SSZ/7u3m9cwBMz6KjapPLPyyGZ7jwcZJoi7JRwc8qGBx+PF4Ol1H5ZMr+
d+BTNI+hv2/hBfpoagBeW/hXDWG768UzDJwCYgo2VEXACXxgCpghczByxYPa2OOZ9helkTC0NG0B
Coi2CotZe4tTqQdVL52dMMeOhKIIAUHgORYYCirjxC8ilrtBOLJTk3zUJHlOY4TyEJ4PDsgG1T3J
bodmjwbvAXQqMoAqCh5kDo3ZPRUh2pZprgiy3IVqb9pABKF5+q1KHhz2L1tCzb6+G2C60+jjm4SB
EDhdV6J6GnIlzgzCRgR3enni4idxEerVGADVJyIKfrkNOP8LAYZ3ErRWFvJP6grLZqwtmVEHjfTo
dc8zoK4itINX2HG3w0LjHTBbft655fQpJZIgUBJnfMGipOM445c73h52/qQ1ggnmo0ofJH8lP4+m
No1fqkXtEE83FrS0Ah8FQOmvJfffajfdFBmm48iaIHWqD8VBU4m7iQWKvUgFWsHCw0V8j3UQy/12
fLjZYcBUDad8Hh/3RezwShXO2FaVniLcUUqo7G9Q2toUsp151OKnoefJNoZHlakYenmdygXFFumb
J0Cti1BZ/DwZzzeQktNpwHhnF/lIUZ153nOSKlOooVQZtdCHsRU3WdmvSg17KzqM3ogbYJhZ4TJg
O5+97WRYANxWNHBpdx0DNAlAoqJ0JoC3eKR6/nrtrEjEKqWq37nNutJEl+JUrl/ep72QACJBsPPB
78tFsBZ8kb0DmrpmmcHX01hoZGv26cW31y/yYioe1aIozd9t0Hz/Uiw8i88PKwTZQmIxvJZiOrNt
gX2fVudxqbSfuG8texSdLwz3x+LJF/JM1jlQVg/CyY0V7HrC9lFycLNujGVozndqgqzUhuAP+E/o
yr5Evi10/92ruNNUXLq4o9vZk096MrG53GfPAK120BKk9ISD7DoYtOkuZiM5CB5DcmUSfoj47SuA
EFPMMRiQXi1bNYyd9WhlsTZqGQm0c9N1RDPEoskAJf9FqYtxUs3lIb+uSNDkTEM4PhxiNNR0AaKa
x3BrYIRirp8TOnWomgYntrCr2nkYg6Y/WP7IxGw6LXiAH4zcZBdRCQndjjiqYBQnEMU+oyz4YNRV
C/gikaQ1xTmHsRGG4BiFnmXmZSm6KqasjNkG8vHWfXrjMt+WZTc6ss5bw6purS9xZ3IxaVULPsmh
8XvvwMZ9jALr6hPzv5fjM9qRajr482ehqH7U6TXBHtG6cGcJkcZ9Z2m0iFsevN/hnR8WcWY2eYVx
eAU7sRM7Xd+u20Ekf+TOLOElguusU4aio+LginCIr/dppAcSWGUBEQIHjP7/r8Wg6lx+dclCl1hK
B59ta60rgwGYH8N0u2U7ktWDh8k2ShncJBvjzsSBf21VKloQfrXYEYwYyuSF7sUHPBuga7kMmdSD
jaQGOp1dH0uyrvg5flsKPhlCZHJRo1D1/afZBVI/cvUfl0CkITOb9lO2GPJiZMXhO7bWUUOKVdif
vDV8OXWUJv+VsSJ2NN0NXO9qcL+IM5nEGhdOBq4qO4yiaFU9VHPFDCntaXci4/d96UYzn+bmjZFV
6HmZ6OFBZp7UxmDc4h9f3a6F2WNObnwaSYhTB6rXYJ3+h7lUKq7JV5o3v1f5Pff3N9F1/467HCpL
JkU4gy6Lnp7x0xcPQLOfYHskB/r+NTTi4DMoO4leAyI4n4EM/6K5EmAlHCWd3WjkMHS6JEKR+s2b
hujInpKxIRYQmXynvddVVgKKHJJEx8iqF8WsKmkZ8hkrnoOQz0O4EeApOt0KOP9AIxa4udIynuQn
WBHayUSyvP6Tll0umGxITk2aWGAiswckFfSOakaFmCuV6U7ZuI8IWxWEqgF0h7YgIGsQpxRQmooh
UjDgq64AUd6KprLqIp9SVLJoVBHe//Bdl5DS4Yr3awwiqvdbhCk1Atm52T3/E023obzNrcajdfaU
Z6YwSyHnGQ2LE0zGHQnnluPp40zZXetne1z81CkvBDj6MvLNDkNk0x/agTE0WRBWCVVtIYzIWq5Q
/UOLBGG6sOO54y7lXESkoAacugoy5a21PtSHg8vUQpUMydluwNCSZoDnQKYE7FNnIVJXfW4O+UNi
4/0FnqhRE4wSc9nuu4nQwHctN8Jt/Yaklx9FzOol7OsX5TZC5/EcfXs2B/qsGr1PuEYSEPjSuOkS
58lx4sJYo5+qW7cu0dkYDCfQ8KKlP+GgzQMD6dCkbEb3VCAOblRfS0NTYlJcqa5JKyhBXlBgHt/w
5O/wXcKztN877Ep5CgpQENpw8qf4qChW7Uk4dC6kmWdyySQYkYY4AdCKqSLg9lp5dbElFlAwBQbi
QjmlqRAkcIM6lwjj1xObOSkraT+DAWf4cAS4CkOtpRy0O2/rTdJwl/RdvR2K1Q1OnKPbZFt6Qunf
gW2hHmWLehZXSTo/0VKvuCstr9rZAAHQQDrnSnjNz/yLzejAEQPtSRIjTOZXAtYyZDR5xvYjfUB6
UF3tc2F1tUDAngTvhTsexyCKXLtzw/y0hGYKMP9zAbmIZCoq0v5JP82jTnu+DN9I8zz1zz1RxBxt
4Q5sRfsdMlIxy26FVDivryYaXxh6sANh/m9avzvUYqya2ByfrvnEzOWNjalS0Nfao5sjzxdtSFEv
E52Avb2vmizJkuneY0G0GxEOGdem7RlJlgRUZqqOx7d5G5AHkl3WzktBTTGvRfQfjoymCfAQL4HI
qhwQAKAQucwxuKtkX6h/kyQgqbzN1/4Ya2Uf1bG1pJdXXxNhpXbPDj3yNJRy/mrtT/5A8upbINXZ
Rxf20bq46WV3RLmJr3oRoTZwuo3wVTu1htWUCodzgrjalFVn95OtN+j/14YO7T+v6x1N2gu7H/PV
WA==
`protect end_protected
