`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K/qcDtm5Pa1moPZ3EOIWrUiw79e9ekh3PpuLWHvJ5rMpNoPyyfBC2CK98DevPX+TMJpy6+Wrdyrs
1vcCHJTxfg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P+sC7/nd6RO96rQnaoAyihEzWRUrVFdJ1h7TI78j9eLqckFThAcR+hzaRe9bQ2A/aftfydiSRWZH
GI2jVMJwZdcHyxrA7JLlvX8lTpZqZiNEmfKGOlQA1+Sh5SMEaksQJYhXBYhDTps+JymKp2Zl3+k+
XBybapbKFpqDVSsmA9I=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PoP4iRxj9eiVMv/HXjXRiRxB1Duw/qi21FMWTL0KGf6dyCzibDiPmowv1LXU7lh6zj4qUWNrYsKB
3I7n7s4cxwMzJOh3KUAUv+I6mFoJ7jRKCKrvXFipymLf54OmUA71bFGQx4StOGd07Y5wzPfDlPW+
wi4lB5xL55b5P+raDfa7M27Kxc7Q3k8svZB+r83D3ILBTt5NJ28GLYcSqIvQfL1c5iZpiKqlcqds
aLUS3gwDYBHvSkFa0A3jddAtqSEILwohKX/t4NWQckyJeBYfnZrkfMkLXR4cObbmZ6+tRdaaNVv6
dgmwC5PemcKyhQihUSFLJx+ePjF79vFhFHJGBA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JcVd62StgebmI5ntfCR8q0k7sE+1O39G8APRm0X6RxSADudii/1HoE9x1dMhcRnPhkzIz6MVJCjO
+nVdNqbLhvJg++g7t6y4qcNaG64XJNHqxu42XIT5agA5m4Qg5eODncnGKrM4MGPj3Y78DbEoejqD
0sSZo0EEgetnV0fRP+Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Uv8L6cnBQ0rWS3Kkum3gzbAFJVs8c1f6l3XbEGM5fgZ2LjVBKBR1ZMm2vN/s3xBBLyDinYEiJuRj
cqmtiiBBXTbGTGP6sAjjm3Uy94Q8hbKI+oUMVOwgCiixuW3rfi0EYiHX3/MSKthNNUq24QBmQiZL
JRDVHTt3tDp4oJzBvRP+1gRnqHbxuWwwKGb2HFQpEkFSGpm1Bm3moBgEsL1OqQbse8Ajyj+XbjTA
rvEXHfrP4eFCP82VZHZgieEOboE0C9Q/XL0io/jHyDhVRP6QAP7FoROUZ6IjTavr6zOzBzUWx4tY
WquxcGzItQUuUkaYk5OBPF6i4G2yM1RMu3yUUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16144)
`protect data_block
vH4KCCBRkfZXdv9uoeXiDQQUU/rRBDnX2SIPwtcQipWRNvil/dM0rKUAOEs1UXW3UwqD6x+DUw+U
tVMdtBxsYcOfexAo3+8f+Z8itZFklcp9/qOVSKlRJ61tnWm6gWspk6hSVqblKZZsFY07/kdzuHIt
ENNuAUZLqyHZxbmZ5lSP9CmIVFXs0fWoV3hfINUXP0DVrvJ8SomcNV7f8DXcba2jNzPjrAlacQYu
YYHDCeiwcyPoa9iN3GGpvBITh/nZxa9WOwTUyCxoCW6nsszSw6fMzwZeYNRvwybU2cj01ZlSU3uW
Et8bafPjztRWAga+zuG+fxaZU8PM6Kmt3K1wXYBXhbiJiXkcxyImV44+YAnK/r4+ovncfOTYAmP9
n1v4+FCc1GjyBdffv34f/9jzh5/EFTPVHKEYgE7RxTs2bE0/8ak/wQ2p+LUCFdgiG92uq49vQAsY
XuO8DROp8b8TNagm/1ogB+Rwq85sMZsZFfjvkHRNqRPMGLrh72QWlfJqQBy/lNFfFV6cnGrnex5+
hE4FhoRED8zmhvTynF5wP1P0Ccd+kxeM1yNRMkQd60ZeHMml8AXkcfXMnibL5iDSyQ/1aA+jufJl
LVLJLokrLeZxuu5lcIzOoL8uM8XpyrG6g77sPdPsLZXkn1Du2dHZXVepuBN3GJ7ke2W2QMoswdRO
2+yqcaOM5/Ut98y5Q2yUPdT90m0XeOKLG9BnXRSzufteYjtBCezkeXZttb1v6x+Ld4mnNfJ3DJhh
RSUsgCcCD191uvBjSizmjfg58PH2QxEVJsfAzUtwTWHWzKTBZ+UUVFM210oK+isPx3v6lQXkO2AB
cAHLEmCQmrkYIIihfiXIbh7XqA8no048g5FfxJz8kx70l8qHoWp+N1SUH3IbeF/H24mvoyfTJ23R
s5mNVvV0pUVQsF5N7Zl9vckGnszQOUhGEODqFIUXz/OBUYAUTdqBRdsN22LL5c2bkLQrKnkZ5wZp
oZZj0Pcmhl3fVP13P9Cc+JNjPucnhxfvxfaVNm4SBFZxoG8Wmoiu4OH7w/hDJqOyVoHFxr/hOFMd
yqBgnwpzoZQpMj1lU2zuMYQHek9zs+QVnofv3X35PR4S6Xzsr//XlcdYml3OjcRc0QWEJ+MQgUWe
jhLau4usW+rbQI0e0hk6c2Ou7Ey1nqIWldfnrb+D7PUk3PBUC1qx2FBe7sCuatq+mRE2cyEGPsOl
Qif8GRHEoAuXVHY+1MV35FtQmz4FSSe/ijUifw0YaaZw9S2oaMHIENbzE9pWhq6z8bd52WSY312B
dOf6hNMusTCzBTKottosPwAc3BrAnMlQlVKp7/jdEAiSXwC6Zjb9KoVQtu43DbcyDl/H9fny+dBj
m34RZzs12dyHN2tPWaLmNia0+gOFncVXL1xf8fZljU784feoVZd04GRaRpXBtVGWuZzAz8hqPodm
CKn4hFoAk/HO735kM4KaA4d0e78VBx+BvYg5h+inkTo0ctYBB2v6qjT/BlQm+5y2Mi6+gakmvLBW
v1bThKiWuE189ug3TWbTJPDMB2T5ohttmxNPzDKFxIi0wUzr67Azu7TeCQgt5jezMQzKpyqnwwN1
hnZgvhhononv0IjVxPCODVeT4HZ8M2rcu9eRuSntjqLwsU6BnIw1dCpg6+Ck65yG5fSpXiV4LqlQ
ThzL51a5USEljQBWteDpLy6bWecrQxcCjV5kcrTZKYHimoQO5A/EquifV8iIBIuBBGDKJfGerL+k
eKHbRwlyNeESe36sYMCt47ahDIfapZqy5ZKQ1peWap0IEoxhcu8P8oXMHjdmK0jQs0PLfycfpv+e
R8uMl3w9XeZjSxsx4BQiDGS5vB73TOC50v2KwQ+RYlAG3UzQNn9EmIe6IEHi4386v7F9FbZb/bDP
zQPqngsstuoYyUhTTElsWvzMSjrJpSvPyGTGWpco1jdteRfTx80qGKm1E2lEn6sv7UTFp4Exftcx
bs7v4GoXptiACSvk5OXPpflz49uVoFLOTjUwt9Dz0Cfv1mmlHe3eRliCAXcc4vvzINX/6obziaQb
bVvhMPCw8T1M9Q9wak7ZUm8agABWynQSGJ/0YQRDyO9/KgLGm/WPBpIIOlgc77vjsvlxHaAKT8/5
JXMk2yFrQ5dvUeC3KTnn1sMjA6Krsn0x4ByHWbCB//oZjB8i4NlYgHb5U+4qJ3ifAuo1YpiMwW1f
DmztimWkx/BZflSH8lZMnNRazW+k+uZTWgmodNOAmyKvZyr2zz01Y3ziIZrsMmXIxnIAJqZugVOu
Smg1VjE015G0kw/7Sz05ECbizF1FpPzSYULJA2CRDaguGZk00hGCyJWtr07jfqtYP6HlRq0Wfxcs
JYR5l+uwk9VW7JTQjsQLvuqMUuecDHyI9berZqA4JABdxKQpauqmdez5fiZMJcVs9sHwUZK4YV9W
imxSyw/2w8TGoG6mHUwdOC69833RPdZT2HjjxpVTlB6fHp5KrZd9kfQfpl1VoHs7i00RYnjlq6LD
3YF5keJ24QMJICpSfDMFYINKS66+yRa/EqBdkLhGhKwT7TXE5GNl0BHdhNnC1AywTpt5g2HrF2dp
raPBQc2uX7vOc44x85iT3wdDrGtmERS7RsGn/GidM95+3Xw+e0/GTkEYL6I2KgyZWflnV/ggdGxw
mcfpzTiIXR6or4XjfF+z/m+CJW2mYrzBo4X7d2lD80rDgv8cqiMpXBTW08JoYW39J7f1BU+iPKy9
iAPHwS7F5s3tUMngy6iX7SdYEOAqOPQFwXy1OEbPaG6qu74t6QHycNEH7lMpaff0QSfO+G5dcBxe
Dp5jit/vo1V79oZXLMT7WAISPFK8FoyedrKj7i3pJ6S07Xnou8qYnvWJonoNV3gF+ayZHvq3nthB
gQBhIFYosBuieqdRTv9gT795fJYXnz8QxLkxRDA8KCC0rmBYo9mMWH3wuhHMStkXmccVc1JgX2pd
l/8ro8icqZUirpmDpt4RTJfhipyvcdkgrZOOjbWT7gMsp7tmuWVE01WPddPo8d/B4plZ8jZURA3Y
sVs4V/GilkLls/RJLo7gXUGRNjxcJ74g+f7ywB+wBuahEP53VLz68DZsKlYWAmCPEOjqF4aYy3cr
KZ8gdAjXQYekMbDqf3W79T9OWcV4THIgQp95WFL0hLtjot/BrIXFZta1KAda04+DmGr+F9xhe59T
sPxlOgZqssQqNfVdA1S1YaqAaE/JF05mb1ufoQV943q4DK9arrmLFeUvOOeHkJDXdspnG/hiqfjs
hbpmY7AkWFKl3KO2cVGqGepvTBcM4ymUzluYR8DKsHOrM9LQ+g0PII60Ak4cdHlzd8/I4qiNkFMl
sSM648roOxeeOCbc+gP6rfZ5GCJVqYKwY8eTc729jijM7tqpPe+hjsija0OM3PBKte70jIauWeFx
/U9WKwIjPCLKLTrk7ONF04ahiS8z26deelS3gI5WcIe9lomEk1TC/loEv1NDh5Gjs+JFmVvLoBC+
1ll62zipeXGgqh2+k9I80rKMzqN0FtJ55iQk6OPTL0hnKh7jrhHjV5nbCpbQzrUDULqyORf4Uncu
V/aoZcW9EG0VVG5ckHOv99yFepwq2HZUUvu2PGcoQmsTHQtIY6HZHn0zj+T9Lh7pA2BMrIKfwEqu
A4M3mjjfxgDqRfebQypzbepFYyBJZWQeEetRXdfl5tfenecjiYVSH7qmzdWCE17iG35nCNrgjO4s
sAn9XW7bw9++MqKRM4PosgWE8/ksxsTi+MP4Cf+aDOUeP2sv7cZC4xlk8wrWj7LHaVA67sgylDQo
eM+Ldgg8l9vlngqMfoi/j03t3f9dGVM1ws9a/67KtQe5mECWlHt9WiByHoiXNw+V6zt2k0kFQ5jk
RfFeR73bABeM2Ey9wqEZwjrtRc9JWAyTP3I4m4VGE3VRrCa4HEk5rOgs9rFayFFotyzJeD1dGnvO
g9pflc7z/eZauFIojfrhZUjclfRR+tbnIosXiMvzraSkVtl4DBiHQJpdnHfS+Tx2lmeLZP3JG5Ay
6sduRQPPyAysoM53/eJ+t7FUaqM+XIR73SDyD7Sh2qgkE9MNzi2QYfiXHqyOecQiK7SImZxO6OAi
Rglp0tqSpW/U/PBD1qO5Ag7/AhL9DwmoQUheIMCC+gyd8jPgivTvti47plNy+xTKdKs0iqJwys85
kr45VoiG0prmobPcho+wg1MuTaweuiGoUWwPnDNQDXOeU7LjYtuVw8OlgKuKt7idYWCFJ1UXSZtT
K+QoPOCl2vanWAOljSEw84gg155xmRV/g5y0YYnvUxyESB1RotvxHjVkAZfrWNnL9zeno8XU9VHN
XtYxjMD6f0IIR9zSJSP3J28UtZQEkaiUzJqKgsvlBgFi5XjGDXyHLW7hZodI3/ZikuQrvqttjk2n
ot8nN4Whc7F5v+vy7qILn6+eOl+b5qhiBr6D2lbyPcdFtDGYogbCvBvOlNQr20087+3trfj9Q6Jv
r2b+p5p6ZIzaFxKQOM3H0mWRYa+kJ6CIxP1HjT87EvIwbRBtzKB3iTgjrACOFik3pdO7z0JAYYTo
Z0KczWe1naecdzfvoZPd+/w/poMjJ5ENfkOhizBd+Nh40VcysvZEeiBa/knu3JpjbLhTDT7XUdrN
CHiCUkT2pjUrciX8t2tZ3NUasMBHPcE4xLXHDq6IHOPMSmoSBvc0jg9P+89cBVCgXK/wgeQvYJ58
KdD+VT1aWfprBMXwPR9D8q6X0G4qHcRBoZfTrmfGFcpm3FfCpRkwAoK2SeYFhrLhK5MEa/9uTmtG
N9kWDPjnXYtxDsGYoEiR+BKBLMkvA4wVFgoo52H5dz8T5OTlWVbFy2LSSnDdv75O9qG+PSATphJ0
C4e9hxNVBvgFBYQIZD2x1I1LJujMldDkKoyWwCCzeUeq9QqtmEBEVmHdigtuTySHuhE/r8H03CsK
fxT1sLmaQ2o0HCWACaIhMlvo7+kUd6aKcik9Vvsd4aZGAzWADDRghnsmWZ0EgbXbKt6WcuQP8nEE
MUYjJMrdi40XfWgyodkQb+eAPj9fdRgeUdIOWbMOBG7QGLa8GUgEVbv1c1wFjAuOgIX+fm6Vih1M
b73hjpaVeRxCoQHI6RZyyb2yWaEx6k0KLI4Wvsz5f4XVKHwYH7ldjueTDrrVayp4P9b8f+WQ/k2e
pkUu9dmklFAyBUdvqef9mn7FvNg8i+vvEwgbbta2ogrkVWif5IgiXqXkzfjY31alvGjY6lQgSy2q
8BsA/gaIrEeHQbvjpDM93yikEpdwoa3fRjZrXEESbqAQSNtYUIYPhnwNYpAnpaG5988lAs9RAo+4
NgA4xVMp1CYmwjJ0NCetfL1ejTgoXV2Wsct2eCBOI1VC/Eblo52sODuIEziDet+bgYoET+19vicI
1KKYWk6hALJUJiHRs68UQt3hobpU3035ce1DzoYM6O5FHUtzAsZ+gu5RUuJyQMZVSLn4C8p8bG/0
zkB16qLJS7UOWF4fDdsFbYA60hKXGu0esoWh2YG8k4MMxH0yY828uUoWNV+x4Nr+CYht1ZCy//ck
DdZYraselRwP9rFMVPRdCn3Sgq7xxoL6OQ3SYCX9oRqvk5OguaDS5QGT+DqCCieH1qcR736aqKMn
dXLVnOXIHVcehJZc779sF40pRlZx8jaf8rlmdyZt7fGSNagNOoNXxqXHAxND49+MnzWdjj+U7+fh
nbQY2dtv9CrY/h/MwqHDtKY+fmme3iFj4YbDxI29SCL1/1l7RzXgdu05T6W0h0vREhyv5ZyQcV63
9FutEqAfIbqA/6lu2N2RWsEF3RffW2bcD5sao36iaKrP/XLPyv7JxkawguRLzd+shDsv5J+I7rqw
EkO9q4uPn/fsDkGIPqE8kRSgLpDQ/tRnShEjYPSedCnW942mRy9NfXMDdVbpTtipih4H1dvQQBQg
hrUcI7GplkdSRI7UULhqUjlie//mAWIdT3JASkP1h+wWj+/Wg+s83Z7kNzWX75leA2jGZBqMHbua
0BhPk87fFdjuEAU2yBjCSchmfi3/IeV9Mx71vHWq18lVowJhhCeaFteGJcU8Hz+SKEjpeOSpfif0
APzqGyaaxhbM8uhUlIn5pUYS5eljCY4D5e5Ji8qP6KamAxJ9FMNsclyGLRyYOHMuwhUzT00qieMC
/jzNzwo+mbk6+PirU+/fDEqrbv1ttcTxsAhCv4uCGA5KAsPkMGVuvcEw/fYNxGRQi9Cbap02wRuQ
OM81nCjquzbjzwBtqsNAxF1lcnNZuMAu21neTWlg6r+9bmveqtGAcKlNZr/BEddG95BZ5QGGvDFt
+7/DwwXt7TUIQFe5ydNuK2DF6iD0BjG+PTidhssyYFlaXtOABg6hqLqaEGueuKp6CIwrrwWRV2up
yT/tOzmGqEzcWkqsEckbfeHkmWuCMv3gPFCMCG6e69PdAOQptyDSuHb2FoaPD1fukUi51pSSBBFw
jDi8ZEYTZcGPMyKrXoQLUZVbWV1KQ953rS6uSE5T+G0ZMtFQx4sApMsg1cG2vvNrioi8fiBKmKHx
TXhfKkJA8SeOxj6PDrnArhQjiZOf9BfBqG2yzpDaMff+iDReHhqIjMJkDkx9yMHUAY7rayhQTAZh
A35IbxDpSngGSHb0QnfmoBn4C4x6GxAPuBl2ypQwMiQ0jP6viYEbuZgGzMD2UnhTWtkDP9jNdoGx
+uAkXEIdoboiBi9S0lsUtXYgKqJM1BqM8hy6b/bcD+jmMUR5uJ0zUWGF41CfuzxuDDTeg84reb4T
LZ8LtRN3IlwdZqdm8JMOUOSbDR10rIB0QA3vymRGbBG7QCD3Vvca6cR19d5WntnjQKKcAZGg+lPw
U0hpavnm6V+lA5q62S1c0wyBY4BCX1cirAcnGTmwgF7Uss4xL1jM1KoduRp6IkXpB8LoE9flEn4d
391yUBnM5zu5PnZsp4utLU3kvKfLpsfwf+/RD/ny1Rpqeem7Infg2Gm4NA520JxTrO/rwbls7ean
fOCwjj0vxEPoAfp9lWTHOaR8ME4WZkoYzr8VZhLdTlG19/PaA9OamkN6apzt3t0urnptgP2blLPv
lr0BwIvDQNo8e4Ts9egf4mmN622Djyu5DQRRAmVENh6KEU2IxCTlyX9HJU8OZTTnkAbdkYkLDpf5
p1PuRkbWzSm9XFSKXdUGqMsnUb2t2Ehvc1uJhHS3NJsCPiSL0pExrLonOcXarOLS5JU1hX34fD7y
OKERkXvsLUMYnoQCNKsJ/U7vEl2i23nSoZcvzX1kl4zQwMgqojDsvXN4n2pNcilori7+wGbfHhO+
WthE3pu/AJtdWbJFS/DZdv2AV1cuxqrNLd7ecLkXscEK+paBHh1pZfqGTX2NLNVsndHa/q9+kvBm
Be6B/Vq85gmhFAfIwS2dG1LmFQk+IwzhzNPwzDXKIpqOmCEYNs6bb+LGECGxrj5JFlxqHG6wYxqZ
z+cXZfOZFaUpTOpLm36xOYp3gLiDHhZuM3ixZF4K3iVHrmmPfGT2sAp9RbYORT6AK90VjvGN7lVY
a0fwdwhHFEJe6ECK/nJRWOWcsnD4eDkghgPYVCSft5cnERKJDHEnOQ9HxFdXAqyO3WqZAGSKjxAk
vkCfN31si1XQiItHNT9rLMzCSf0v5tQ5yrgKfgreOyj8jCCuVRDxHBUm5yUKuDFsqtmdizorYoS1
64d9ZlywzG/kIHQk66I1cC+mK/POFOwTf8dRnTFYparZeqsBJ60JZ4vsXqto9L188pLaeWT1cg8W
jIMEF7oTPWEIhniJ5LBV7EJcyywqrIi8aK68qddp0IihdDI8m00cQIDxQIUPu9I12FzQ49KY7S+w
oe0e3uaFguG3DZehsxL2vYLJ0w7DoXfPK4Oy4AVQLuGr7l4RD0QTdXkPR+wQAeNAsW3wSFZd1qXU
n1kzUmJRWhHgUdVlD4MNJUFZZtKCLeoy/fG4yMpPTfK+c+EpvFu+mRwjZvSNMzAjHScS1NgaXqpX
qsvWs8mg+rTxmBnOodTkstJdXyqJnzf56gXG3eTrnDk6Bw+PmPCTgievvEcqDUDgJ+MTMRRVFt0U
IvTJ0W1kg2YhZ/Qb7Pg81nc+zysGsr4CTm39rnhTxzAFjAcj7qcZE44qnYszx3RBvfBA+Kmlgg5p
9G0Sm9TQ9kmzBEoJkEbzFeaTiBRjZAkcQCqqPS8iRZ+OL1p0SnxWev22qSyEFv9E2Co14wRBk800
xHSYBjo3eygQz66Wc9jGT1ld/eDY8ESkXpykXOeRrXxwOYo1kbJ8+m+dcv2hW581MPy5+oJoTTYJ
3k6TyKGveS+DekxE6+RwGTEJgqP6RA6aWmKhYuQBYUTKmWTTfl4m3D4zab0VxY/MntgeXd0Q9EB8
o6igm+W1Uz2CPyHlPJ1Fzw9ZTVGV3mtuKGqj1hyrx7V2dvPBCCyG5cZATxsxFHXbbj+A1syRdSTk
mfIfMvac/SzLTT1qCHwa0/dm+CXi69UCR5bSCFU2ToZoVlB5As3G3CBSm1W5My23AxtYkcm3a8zm
XvMNiwYImGUglzk6bd+B0CDSfna0hcgrAsqmynk9Jroj15FgJWp7ydBssLTOXEj3bGGt9rfYVWOn
e+mm2MrWZlozIVy1biHAoM+CjDSsx7dGA/2XSp3DoVXVG6HwurtWWKOwraBBWXoKvdJTy41KVqSr
IjvwFJzKOk7VdxwXyqUfH2FIvwySAapxSGcuKS61EUGmghdqWWBjMH+ehdT9rXHmEYne6x8EnV5f
7ynJKK6pxXGr+md/Bbs3uLwaGBGK9AwbQj9jUKys69DdxECYo1aKa7vqYZ8oI7PPdVg1y0oSS1N+
f9H4BB081wNo9YbUsEJYJAAE9YxL4wkihk3oDWIl5mbx0HcaCV07Tx+L0J7qfQg4jzot0igVANYn
b2FOguWkOcmavdqcKIeLwGT9B6m5bFZeITY3vXdf1yUfP32zG/fK35ge7Uiqi3Y2BoZOPLFnMaAD
fqK36Xo42nDk7jIjGoN5FO/c4O/dQpHjEjUxTD61O3ntKPpraprkHmJduuunT6ehp+IJDAZT0gsJ
6ie6kuzx+ArIMTlqSx+IVj2udo72AIddlFNDbSsw1DomcHu239QrT7rCX7hvHkwPyD9tqGjrPhBh
4Zlbk48eb9q6IIANWsylBR0XmsoU0Opjyg/59bkhxsuTusp/Qzn5hpjhq3+se2xpSaPSjrlmOi3N
khamAUtPKZsCsKhwm2IOi4Bu5KIfE++Bcxu/fYA7mt/I4JkPzFZMtmNOVtwnC5qSVE3hefg0tNmP
0iIWi0wM1PL7QFwqDkC3yea8TMY/uOmCuBBRuwf4G9vDWSlWB7f7ZU5QGMz8bWUP+ktNDaBiszC9
1cwyEgFN3wHLZnbMxlchcHnhSboMWJ8PQ5X8w50qyVH7Il73UbP8NeVeGkPRVTe5l8D/0CbhwLVz
S9W6bhMj20myhYkKir/tpQQndAhrgSxiI65jSW0Z9lroMs3DyntWqss73Uz568/wtBJL1zdjEObD
/uHYHJ0C+hijZ3OU/HJLi+FAddXSBHUUoLk+6jy5xL8btsC3KpsbJf+Alzgh7741tuU4hvqcRgsM
4AyisDr8smKx08gWf2saUCrxElps5mVWe5EXbiyWvOLl5roXh23f9r/Cv/oKYjH59HRvPuHeCSdl
q4D8ljR6mK2xECB2ZT0oKFtQnd7Z/26CF7E8nSkI1bsK7fmUChIV9F/2D569MPRGBo/gVW1XPyV6
T8PDVRIkwF16hH5oU8UdNUqln5LzIy8RxW+3zYQlAdyR+dxZBrN/LZP9CR/IovsDJQ8Ych3khgXZ
aNPo8eCXAYaH7+DRFwAQN4Gs5ktV4pQRycK2/GYDG8679eQa75MQpE/3oJKE6hhi2oW2MmhoIUTF
rMO89AfoRo3tOOy5QNFiUjRw7USrtETOGiMBcc4RezYvbzI62Km1Azeos5jmD90gU1e4aJSRNVc9
0fmD90mSVlVUJ126E+9vjQy4N1pT6C1n2JeI5VOknyeHrbgI9MREXc18SN5dXY2pGl/2PPpYF6Uf
CiiZ8XVUeL4IVU06bOQ7tg98slG0HaUHMQJm3QjPSUHIk/3J/FH5eReKER1GGp9C1EVHxYucjD3+
AUlZvkqk175J9RkbMiLLW/4a1BBBayOr+hp2lQfXEj9ztwhOmJ1RPeUCuQDKTt03B2Pun5/XD+sG
ewg+H7/ZkEHwDa0cCbqV2LwiDASkCxWnv030XKt7WgFVA4yHr0/jhZ96RMEsCQ6uNRLv086J59Y8
4AqP2PliICyX5LEzbsrkTvaV1pUPmqSPHOfHQhfdM0RvRED1uyBBRiw2slIEc0bZcbvfFoMaRhl/
JBnMh3LVKJuh0ZFvsiBuHnX+LalN/mt3OowQ0+y9abFuoiPK9uNuNfB1OtoIxUZoWETInh8SA0o9
S3z1L+0VZGrTIaseot1JbA/o61duhLz7nyWl8DKz02+DwJ/YBsbSxuFAqFI51zTD+IO5WfAMi9R9
6bZzcPCS0YAkF0SwUAZsYoQOBoPc5VK8A2U9+G2xPR4m1IUfqpZfwv1Sl6IX4/rYw1jau8xxfwSM
EUCquqwddH8ttVX9AFnKCUTjp00yfQsR0PgljgL79sYrYMiU9qu6SLWvKyaCMcI8avFRl2in+Vam
bCer/jNS+BtHvRuGZY3DQQEMqckeso1D/ZCkSrmLTJVt7j6uVH+9S1soy9cuFJuLzR97n8z1vES3
gweUGnmRWb4gg7ohTCaugmfWB5WW+WdsLIR2IlTehnDN+Z/COwfu+QGh1lvUDJePPSxmhAThbLR0
i+D41wdf4z61rgX1yeaRopN+Wif5NCG62qq0e1tSt0ExYRmUtszckiQiNhg3L+f0Mfwi1Z3FCfQf
tfqbKpWS7vcpJn1ZJj20q6KaLC45DAg6P6zGllnyawCYT4XoBKKOKciRygGSHVRs/eHCt+J90JyO
+pznpIF3M5pTb3OZmVXDvVVQR2WkLKsu30dpd0fC7u8cR+XzKECmhYlhAzv0GPdn+V8NKcJ8WSeh
tmqFB1EBRLRI4hmGT+4RpNhVRV/cON0p7x+6Vt5LJrCucIG80d/oA1H399Yl1arHAF2T8vu45xjF
wmDZDHC7z12URRKLhVRS7ZvmLnGd5qjBjkul0uSjLMKYk7QtoouGcWur7rdZ/Om0mdhHhDbY5Twz
TBfaO5w59mhlSEvM3RouPEf5WHINWpHiGczW8C2uBlMo3ibzEh+2ikaS6Hq6WFpbYY9wwh9nc+0D
9EryxLbsRsP1Let6ZOLprOT1ehglDnLJrSDBeVP3Q6dN9GxuKtUDSELOIq2QkeK47MksQbdWISE8
tq57MfgbTIbaHRffAN1PJcrD1NMecUcqXr6zyAOOE8gC1YzSzbCTmrCmM0Q51tJruRp9XNVHzOHI
t2f2eB3CSo4XArp0FuGyRN6RQ9ED6LjkTxYBgV54e55Tw/1qSnGnFyyziGIBq5oPstuy3XbVUyzD
IIu80+ISY/6XJ4cDhw0o+vQCV6Ig9x4lhtvn7Z+4v8ZBfkdAUV7SaotN++YP/XOyC8uDukaVh4or
nUer5DhLdDE7gfJYHxcK2PaQSHinz0IjFtdu9EFcOFpXFI8SIQsIsURGF57MXDWpWOCtKYMWb3+o
wxglYx74cWzqpUUSh5550S/BEv8tSX5+38snTpdsy+CqGmqkpA8fIR6KWxOU8vsG6XLS5QxTT40W
8Dsqd9WUdyIKo1ZgkzQsXZQGgGx/ZvDKik33meEaKIY9ilLFLcxSjUb2T+TbNJgxPf6cbx7HGX9t
bq0i8P4CstfgJEE5/aXOLvfkqRh3e/sai9vTMw6Fiw9Fz9oeHKsWtkAVNwgbRpAdmrzPhAr/20Tp
m7v2bKDA8TxD/FKPobYAuV+1IqLjUVLX2qCa53nW4YIgrKbdAfQCKK84zrhWYV2CZPyzxcyblN8Z
Ih++HjBmKz1WTVO+9i2dd7e9Q0Bxq3m18bSv9TgtSbClpzbwzhSCSEwGvxGnbBwxLDIzVe7TIKmU
tZLSachPUyc1O9278CStfCaBSyeToHT9CnkIyq0KLU64bQT5wRMtIt/yqEqDSzcNz1gvl1AN79oo
2OyCv1uGMHKLyqSh7EpqdG16s5BGedvMz4oLRkzhvuwk8K+eI5TsoM4IxsSi1hDrmEBJ78xg5FFI
dxmugaujAMpcIEYew9c0AUYKl8EmeBlWVLxW0LXcDFzBuoiJ2MfD/+otXtXV1MqH3JR1873jUlLm
96VWFcv2ELChaUnLGj0ijQr7xyqxEAOly5Vt7+dOgAOUwvAFtliBH5j/OqkUC6zN86jsM7Y4FzQt
4b08wyAF0pJQK0peKOkisVVx2sBCvB7x2OR/9zfwWPhebaH/+SL5EEpGguR+OGgmR7UUXY1D1GCe
pR+qVgeZ4XPQepjindMLb05y9f5iEt/8ei8L3CriRKiBBh/LsW1/LUOTH62wx3eQLyP4gF/weT6h
y57aHa9oi1SCV1S+q0TUTNi6lStSIj0H1LlGoZqTPynVxjGUUUXBMSuNuj6t9J65MoQNPZxmoUYH
HIqGP0bAQHqnAJewbS5AmpCu7b+0sJLuq3k/BFAqV7m/wMMvEA7h19VqjfE0uRDms3J4lydrAGGK
nJUvxcq/pEQq9rkCRBAVOTuXvY+7KGxnUPPDjO9YrnYuZa4GjDESNZ/m81DmgYZhONBocxbbe6CH
PiJGM2RrICkF+PnxlUFw57USi5QDQlASMd0YAcwC3cvHjkpN3sCwRi55+IJ8/goXHzojw+AWyatq
xY6W3uIJ9pwVX59THcFBvK1EirhSQJlx+iDruB1t2qHLYsLqnpnoP1HXMuWkA8K5DpKo7jZqRmth
x4XrY7WjqQmdm1boW8ZJKO5rEj0TA5JHYvs8sMmupI6IeicJPesYRmeCSmOyiwn4mpw+tnGKW2FD
+9+ZiLVxV+JB5rOV+fL7978pkRFCdfcW3VsVw99vedG0hJfPnhU5JeOO4iMJEneP0TwLqg2JdOh5
DMHyL2n1u2SOc8tB4hKbB8MGTASez+YilHzdnryu4a3LvigTB/EKdL4kHtzpgeWW846taB4/uekE
ep03Q2qBh52xh+MPB8LHf8M9h7QNmEUpFAiTPHRmh9MA3XESZpyB+G7yZK2DFpFu8vRHDAH1zKA5
hGC8QjBJiSmONEHIMHHFfDuIxH5M2mcOOO4+HjWlgVhLnI1WPQLJM8Z+5QsH2NjlAL0pxGev8M3f
9POhzMrzI+v3dI938o1JDB3bHOHNq4ux6rD27pRzSh/1Tdhg/H/jRkECC8KFK1o0IUUqdYTLt8aJ
pKU0SrceRaNgPBpc7HKDvBWKE1bFYtek0WzTMSjHrw9NMM4aarvkmFWZTZDwI9G3tkzOY1f8bylS
U/sCKNu9wipjN3TUulmP3qkstTueVAboCkWlpa0ntTqNkdL9+2CAIAbB8SHvbtzgYmWTTull5aXR
IC1OXRacDK10mqC1E5Q8S+ysKOTnjaHG42ixEV2wOHQCfS0Q27SPf5lYNk7sLDXt/LaqeK1uqlYP
/5jgr8eEsV2zM4gqYm2jkfNzxXKf+UEwK3Z3mB1iDXLzgwmZXtZ4BxSdVGL9Fbe3mrp2hrJ0GM5H
yqK/X3n/xcwfch+n/abnhgvvzxdvyRQegjpSDospD26D+g3Fq/FMMftoKutZ+hshaOw8HdeJW5y7
Bh2O2sUAWHXn+fNplDcUNdTXhaMkAKzt2hCsoA04Zk2XsgRtTUTrkBdHjoB/SUs+ID+Rep1+H8ht
8whIYqDx4nfbZE5JWfJ5/HfneljNcRDUnbO6s2feRTnE4HEtuXuhjyN1sDlGEUXqRbdVpbFhA1SG
/Lmsb+GrzrNPHXu73NI2AF+J+hxKWZJ8PPQKNW0CEAndjGFA3p+OmAGeBvJS8IvX/9xIjbgqvT3B
y/cQ3r+sjlTX09vT1dKvfau08fFxbD+ob7OeOjCrejr5d1ycWah397vqrp1SzFO6NQqwjDSIkYPX
ytEI+GLDzb6ijcn5m9SxKv93R2AvtvRcuPK/v2edXblCUmDRNq4VUkXfMr1+sHQO2/AyNkRDr+Ku
JYLtIwh6TCv/dMNpiX7881yCfis6f7656iMbSD7n6AWj1E3W+Ihh8CI2Wce7P+BlP5Vyb979dz9C
2xLcJD5lIg8aM9gZho6DfOrBmeI8oXjt1UqAg+b1cbSADaCWmEFQbST2uh1RnSh9nZ62saD6IeHV
x20CbtGupWVzEmK9oV1jts3A4hXN6qxzCBJE7dDeD40RVX+co6aFzP5L7ydDGO1RWHvnqw3Zpb+V
eTQWuN7KkzOrZgwIxzrvRfbWSsHSD6ZJ2L5/bsAoH6WiG09G83AsibimBZi+xJ4z89882npixRuv
rgXzjNzs/ku6LBORnh3VlvwUYtlJs7nvR7MbyC7DCxh8tkhNvz3ul1Ikm+K+7r2qyO03ZSFmxeZM
IPsGg9GkKLmEtXS70iUUefRMnmT/lfDzadsuEi2t4XawHD/G6zasbG5uB/maIc4wX2SVvo/EnvSX
RWVN/R97c+lf/30KdVKlg3lxJsOgnebYy9W5Sep9cbIKuh/V/u6i7HxzlTTnnTqMeDC2ZphSjQ4g
3qqFMqrznEkGyltpCHE5NDbTguEoN+e58Nw0HtELkGn+2ju5HAAGg2nUY8cikCTf/XKC5zoaCnQs
Eh2mY4H9/Y8TBMrX35JPxAIS1XqkezvZRlSYhdEKMAUengHOeddppdelfTcoo4deBHG3NX0PvSob
FtfgScQLrvGGhOxan7uJc0vAiPSocYME83bun0qCcmlVrmQXnO8Mf165WrA51ALC4dIj0IwzF08i
hDq+rqqC3r/fxp3DxIyK4BDaz1nJLPhjhAx80zs4NHicYRXfeZfNKUH+2n/Omc84+0GZnVVdk5fl
0aXGtSXf6TOfhrJQsSH0CgkrACNHql1zHGa+xecssk877+L7uLBOzcOUr868RWAl0uF02YRW3fZT
uCe5XJW3ar8N5DGsBwluPQUiU0C9yQuJSSo68uJhkgx1NNVYVlTU1D5ar1PNgP5dzMv3Tf2skgSX
BQyP+p/vFjtmoK+KFwH465Y/4VJQb8YwHixGaGBIDj1tAsR6ZL/rCijISrObekZ4lQYmMCNYCFUe
EQCoziCLveOh4WCy7EkI0LFx0RFVFt7LOGLqbpu9ssXcmFbGQZtTWKFu4tpQNuhAiW126ZYYpAdX
todL1/8u3FbynpWzrvalQ5JFk2QBApoTuTMlky+vMMkQ49sdFE3VCf8XryRtQHEcVh8PkcJyr0QW
rEUf5xYfSsuHcBoqyNBhIhR6C8g4NLgZZp2ggaOeMD0PrntD5jTqft3WRea8o3gPFiSv0m+BPadB
mQ23YF6Xe0VJRxeSk3qNv0BEBgUWIFDdv0DM4vBKZrrbQpL2rxDKxQVjMqgM/spArsvBow5w7Bih
ifzn1zOotxAt42Wkcx3Dud4blsBHKMaHF2jDyNpgZkfuqlBLOvq2F05vT7lGmFm0nWGPq17HL1qt
uM+XMnslAnXVp7F72ABT3Y4lBRz9ZbIVisSMjFib9moar/ZhL9+Br5bVd7gINPbbvxktSfBlPR5l
+4jb3ou/uAfOOGrn32ATCY2++IFvUzCGaWnCj9urgVraPqjSbAT9qFQN7Bx1rib0FSeM/PfY4iJW
15HuFondnx9C+dsHtIpxOQKCToS98zQxfWkhCWnpLQw+sVmajA8mvGopNSFIE6Xp3ljwej9PuzqU
2iB+0qfJAm2Cpu2tWeSqeELfMuWay4cnG/uff/Wvm7vzvkwe9bLULoNb/YL+l8yoSLy0nNBV4Bqw
ZD57eR0TgyuIJtALJtA7YDEdmq/hls2JEf3Tm0h4Vu9mecgYr1iYNcVh91qIw2Wd9vnnNdNr3frJ
MkRScLy1H7WLe5xc0Yihm63psfxxhJVPhhld4stg6BHI0Sv/LnLaqn5bm8tg9oLiFK16CZQhoCvs
hZzHGu8Qf5gG9FVJ9pnzqURgsLI7kX3meoBWs7Z8UB7DFB0nEKL5BB+bAzg3leAH4A9fOLEz3C48
HZYOjKaICc3S37FJLVxW/0XbJmuHXSQbv2fAqGwY9vd282XVp6KMzwqNd4E/aQKNheJGWrcEU3zr
zxhLvqXC3nU7HNoMZb9z45NUeqdWgwoW4D+6TX6EcP6ETeC9QdrnkV2xeRSkCD0TXZ7SBewK/0ac
9/IKnGdGf8FlyCKMRwVjZw8z4pKGc9LTbE84pqLP0CCpJZ9Den1actUMBle+tpqoieSJXYNvWbYP
lvtnP02hEBSYTXL7oYHZFP2sq1E7CV3V/poPFprCmjY2jsRMVogsfkGRIZuWR+9ca7XLgOqYp606
pUv+HlgxtIQ49Hdp2zi6T5UPqpGP/NP0ZLULjocnYeGFi53YOqFfRi5Gi1T+bp//nlpETCW2jsrZ
VM8D3xb+lA+9T2/HmT24VGBmlWEFtIvHqim0pGbtPY6E7VwGi2OqavgQ0yRhwtd37vNBBqOoLXsp
AK1qx0nEWRbu12vV4AjjyZRTYxUm0y9OLnSRKoNBu+ZPANfc0UVmAvh3OcNq13yCgyDLzPH803fQ
wbjgPXK+B2KJ7XnIMrSloBhyU6R0aSQgLcYe0Wh38oKgu+s5ocTx9RJYNVc9DC43NEd42feSc3vR
Gj135IiOcDDFcJWCN6z6/QSwhXi90DOG23V7LJqHkvJz0hh643fjc94KiQrbmRFmLtFFlAu5Mhm/
OY1e5OeF1wroVGNbGcDb4oWYDaMhiaW51vRMNJbZL49IptAoqP7pEP4e+XHhg1HxmlVJ0VyfOcLp
LwGcdb5J2Jbjx4Hh1ElRmfkXTS56qcv9Uq+P+EiuqHwyE4kSDvY6vepJepImmBDPJAwoWb5bEF9E
xxO5HX8qEVEDZU+NrCPQWW+naLBcCgKIydfKH5bHtqRdMA22lU1O6LUkQCsJ0Rp2JLbz1vmfAI7P
wjR5Sx4DMv2VTd2daWZPIjSDVAXClQoZNBiAJ3Cz1qbNTgJvyZ1O4z0a09VJ1sZzRQInX2W+yoA2
h+PIjFmaqQCRLiyEuFyU3UvilqhgE0B/QW5nQGmH9WYr71AMu2wBz6KDMFYNhQ6qQjitYYCtOZgn
KGuLPOd0pNlz5wUJMYE+H+GE7hCp4enk+5ys6QzhhfkurZob7ycCTxQeaU6tZ7HEqc6D+7ZZcIul
2dpAoR37okH786/qRLoOfJnUyoaoTi+I7xkLt3aJncwpHBQYycpJQGkpNzH5nTNRmrV1e5lqKqNb
rfxXG/hbCt3fIN6rQnay+C2VFvpJiwC3q1h62odOYe3aEUNrtQWLWTrfZYEvWYcWcdMm0D7Z7Q4w
Fe52Li95eW9iigOu+aJiNBz0N7kLMjOwAGEHxlL1/hOQG9dyo0+0AK4Smd3yuWNXlkxihcz4w+7U
CJE93gZHfEfp09h7yCyoq8qzAI2Jshb3F+pqRXM5WpaVGszLKGQXxLtIHXiwpX8jp1hkEEqgrxkq
TqAH3v+B/ImDhi+skA6+RzrQKLV+xA7qmlrgu1kCbUeMBPCJg70wQhwrVIaGIrii7WI+WyKoTHd5
F1tWK3s0M8ibCZc78h8SEk48TwYqHVqA5y8IREMNMsYGF/ZXJI4zRwEdBVvorSawTTS+bSKt72Mf
UPKsVFOZz8ATPfyOTNAlLI/d4uiDgdFFhsQSguR4JE45FQG10x/L0Z78ob4lGtAFC1fNLTGRzkke
6S7vSKg+j4ovv7/vijVtGtSZ4HK6mUsGIXrgN24LBMr/Khyr1tMbXNsMC/AcpMlaV84/XWtVTLZ1
wDqgY7BzB4bwP5gFG7QS0GDPyrRypWvQwTCnuoyjPx5dvVfgmdzc92SacVLQfKDBPldDzYGqsJFL
ckSk2utCJ8IpL04kLbnxejJ1PFg6F1QRk+uoLCVypO378VXvVkz6pLCqbDn0B9KVTtdXk4ZFEpm0
Ng5EArXYf1R2KYmN7Li4yFzoRKRyrhaTJKba1nqcNtvwJRkbqb3vRfaKcwfPWNzOUPs03qTqQg98
t2XWQ2LVJ0+00SNQAvfG+4Gv2jeQcQiOU23kvXVjq6w5r4Rd3bQ7HupH2cx8g16iTP5JrsW6yAsw
38Ya3rMMV5/Kxqs5BnGk7XatNZfFkZ7nv61yzViWbRPWXUukL3tnI4WfmrwwcZ6662JxT4ULS+zq
sx3/CMMa4Tl6w32GzPC0ke7sbu4Gh7W3q0HMSNDu0jt01dme1jg1eCVWfZazsoxJThvV4TnkZZMH
Zw64dlbIlzXhUd+tv45EGAtn3paAXVy0R438OuyZ1X1EWcnVVMaObNbp/W+6LMedMIgH7ZkVRfwg
u2R9K8gfOUZ83DJ71GlJsKkYQayrXPdFYGRH08rhtgXE2nEaKIjMv3gb7DQmub4RnfBaviuBdDXx
CfQasYJSooCdcUQhHQSMwkhFg3T9sFouAVl+pxqVrHDIwKWtiZTXbR5nasq/fQtkXOK2ZVBph1e2
EZ+seC0vjcuUJUPp7Lrg3dL3NE3sQEQ8w8s2/cUp/hfXMe79JPtdF/744a0Zde+pFDi1INBZkUjR
oKVaYay82i+HkES21IA/hmWOgHB7U3LvIpJYld4ibxYPRZOrSINDNixa2fDeigD+IB2kO9N6FVQs
a+3kSRmEfHyk4U4G002shgLh5OpKRN6UzF3wc26S6d9FPHvScP0mbu/ShR2PL+nQV7ZOhd7hy69H
SVGZqaKDEBgazemNqgAEenZ0MexH4Nmb4zXI7IvTC7Uo754dE1W5Sk4o4oFu5JATrERqCrddYqn+
VmK9jUyHHDLpXrpjgHMqCFAfW3+uuLguIBh1l3nD8GZEPY5uRknM5oMPyEHOX4m6CCWHaKjLp6yN
ggXgFYQit3yxxI6aQpJEiRPb2es6AAJYntFIWi2LoXrY0bp3jbQVl9N2tyeguNUXBEKe37iuh+F7
tHa0XfcQSDA9MBtstyNqCpeMmBBoTB00RQVd/PRx6pUt22mWyv2VLdZCA9bTdzOkxEUHFlrMFMzY
1TNdNOsOW2sYlYPYGCUt2TBVLtzpm10nXa3RNTIRxzf3QKy/zg9eEJKJeTp23//d1UOh5dczUMRU
UD7d45Tyepj0003W5KGDhjZOQk8hkkJABf4Jztz9aDjS2G+3aAfLV2wtZx1Ife5YWDj1uYKQY3uC
F+9ZBvfvGPB2qL8POoEntyFoXE+SkI4xB4dTavegi+rqt1Oj6ZSh+IqairT6SHDl+Sc7cfViV9O8
8EgotIirzgL/nciiHi+g7D6yl/SE9ZB0V+JroGnbNKF140sGYoUj5J0SJj4J+xzCGrGCRrapc6FF
fRUrGw0J6jbOscmFR7ZMLOubizB49XozbAy0N84np/yNhof6cVrHApAJhmI8ga/KP8fQvyZWk1Fj
mCUGxLjjDQpkPJR8VebBronM4y7tNfBpeSrJCYucPgV96zSJmWZBKhzEj7qeVKG0OodqX2OgfKs7
KOBqonEdCcqNGgYMktbcNxycA0GtiBb263GvPemFF86GjeMulkz1JTKv1wDzw2NY9MtAeFYuq4zr
IjIz8kHf4T4mkXeMBZTOLas9Qndr8036Ev+i5eqIUAI3lmD2EKjPiF9vU5sDl3Xwzj7RzaZuW1jg
75/w13VmAg6b/W3/9M3krDSLr0OhHZJZpI8ha2sMcZ0HcByiPgwqa+aYJ/WUjTAPYsRLGaEC9uRf
GcBitAuSR4rUgiKstvxzTuvv2DGnTeFxP12Hd6tgV7AtcJrDVvER+ugChJRxdbqKzyURq8RbxUPO
9/twYtzoj2UU/YoqG/nV79UI9RAHdAlRYAia9jUhVsuRTpOl03XKVX7thQha64s3jpY1sxUli7wv
q+VHvAglIWpQqhMD1tQxm+Da9lstODrFH7H4TmaxcxmIoDkNVygp/+0Xl85hqhY9+tI7edwRh3bs
QtI0g22Mu+ql5PtGu48Ib6diy1WAA/+tmMmXjrPFQxFqUpi25bTdwWxuCcevg0NxuKI5ryhuWzaY
zp9XNFVzm5QESa+BzX6DRn4EPs15sdDxpmL4C3X5QunAUWlIF/6vpfCcAW6M+rm2u3Pkp86Xn+OV
XmDbAaFlsOV4Yk4O0RYzf6WszACurTNXmGUopaJi7U5A1zSil+/DIVBOh+9c9JF7Txl/u2WsQxl0
KY93G9ZWRCdH3+6+Zce94PKgXFNOZci0jjuqaWN3GXhw5ZSWFVTrPYKtdyIVXQlUqK2Pssr68SCk
KjelPtqKfl7HPpDY8XIuLPDs5VAeFyVtJd5B3uiEvfYZv/MzBwD4tgqQPCmvBZOpEt00rmgjsLMt
mfX8SVCf0dYzU1kEHFDiEgVUA5ZX9GImQuikKpYrJ0/oMpYrODkiEZFGImVmruhCLltvPcdc80Qy
HlfjiHO+vIut6lPx8AqX29met5JtakH5fJq7Xa6uCFLt12GawWjZejiE6eig49zVQgaK7MQMIs++
qiNXH6JXKv6oxOZg1dEmWCdNnGQhf9m06K9HT01okT1MFbvdz5/ukkIqi5WIsU7TvR2hzqZhw6Gw
FARFb6+fYdCmJIopZVXvzjve7j6FVPaa83Beq/Mbh72BuG87bkZistknoMZ73iBMb0KPC7vpOAZD
vwqKgMdpZIYTvAGSG7rco8QUZmGgarcNs7n1X8R4vom+Yo4cRIXvMrs9mB3aVcucnyhMG/fT3XeL
sl2i6DKKYmxFkUQVNLSWC6k6kpX13Sd448OcRn/RvPKwPsf8+tOF3/5ghU41nH01NBcnydelwfJd
hT0C4G+yD6OT79TU794RopCQYpdQFmwVTEOClwulb81mTS/5RAmzMpDYzo3kI8j4s1Iq0LmYV+nx
pAy9/RqHnTzuWGQzK5xyKTGWBzV/lOvUKtZIRMDRgr5ek30qheYIoRtoouDzC7Dk7KLawx3NCO8G
o7+QOuN631JbW8WIe6tssFITaXPUL6I4JYFWb+ldkQlVRGL7q7XJQBgD/YrGJq8KlBqutN1K/rsK
bcHXNhnS9FIrBOttsuX4/TXTGf6D3TZYWQk/8pzJQtHnXOS2HQ33wvnbBpJmmZ9nbMCMqih2RL8Y
lawtRjo+k6nFOk09rsNuem3fy0XcYN3mz87edYXpXeiJmkirAC8wXX714HcjX0FDqSgCmCasYNj8
p4A6cvgQ8D042wDWyAdJpw8d64MGjMRHr0V5PxOSkG6nqJiW9czkAgPrgK7BvuUfaEm71llorf/Q
v99VMK7Qx+P0GtkK636mGzrNtKDhmw5NNCcMhngdV7ukNyqlsH7vQB9xIWpOgLuVV29yo7AQYrX/
Zhxw7B6PFvdPBLNGeTeb7WotmNyyUECwPcwa5x9i7c43SsqSHWtD2TU6IlpgI+8kNvfG04+njo6I
owvWFQ8lcpJr5cgsVNAfHRW+Fzg6JvshV6hBOaRpRzvOKXh4nXt88naKfNDnBc6/Yeek6KF4z95G
ipwlOLjcVkl1jnk+0L/RvRe1JL740rrSx5Benn9y/Nkw1BSuUIYZe9jhq9G7qgUvmKUyDhkMln9g
Pi16zoncXtSbUm1nsQ==
`protect end_protected
