`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Tjf29iORrKVIHRvtvrk6aRDqmKeJWaLqE1aCHIa7FYxGytOGulU9GnP+DRN4Ow5dJ6Jp1iyZrjQe
ymvaTXXJjw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgpyy3TPo/idL0RHeTQR/rQJdwyhIO43/HQrJDFJpWqO8q7ttJuy2ZlTHW9q9LrmnqRRiWbW2Irg
QsFxHg/47mjvd89BDzQBpdvWkTwG3IGn6k/sbFF2v6BUfI6WdylkjhKIJXbedVukWBl68vW/I4Rj
bk+yAuO7cmWdc3a3Fuk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zl+eTIIpOqO4rV11m9bG45TodRndMR97jnZCKF2wNgWgUqthyc0QOqR8l5fesrSfQFmldkdI4Aof
Jf4DME2EaDxN9G2zq+VgK0o711fQ7DkW2J15l+qhDYa0cITKyqrvJWd/Li+FqLz0tefkpN72tBOm
sjbQypImXMtkGCRSM01mz0vvzRseJo4OXyjBk9KP69bDSB8Iiz/KmpgbH1TiekFd5o9bci6/SxGA
WOOdpTTlPk9Qz00l3OigR8SoIfCUUQTkIyhdjqHmMEW9Ug80lKUNz+xIidgrKiNFezYMx0KUHMKP
Unri2OeUgvaFgsZL9EnMNbIyPKaloqHHuC64Wg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sVFqhKafThpN3kYCJZc3USKnwjYfeMNcG9MlLTuMpwNgdcpouFKfXxycRcYhL6K19lHY5TOol4z5
sYHEZ0JPgNjzZY+6q3g+kc9yVP+rLv97IDFczDE4lyAjLpuj7AdTpQDl4DS14M2VmZ0vp/bp4vdH
g4KvtccX/Au7XWYNjjc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rqUTz6rDUDK4KRpsno9a+KOnh37IXTSclFTnVTGDj5ZZGO/4vKjZsLvOVQVi0jrv2scezLOZMHAF
kA2z8eT58BkjPHwGLyPXbfKGaiHxE/Kd/dGXltHrhDGc3mlJPK7oE+EWVwV+i9aSYzHuMPs1hNuY
GJbWOTMjVIHYjrlCfoJeBYQ67yqE8LV0IJYav9EIOo9n7hqx/OEJEW6sAUxsOIznQJ4NcmLky8hu
KX9SOkCSjltdPQhqeFEr1YoVz0z9RfCgr3a+6gZMEGL8lOwvvMyOJ8ALuZPPfC3m8xX+zv0OX89U
45DdRmgwSZgkjxY0Qjah8z+eFyW8r5ZVZ1+rnA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47984)
`protect data_block
e1EimmuGN5zoP9EctaLn55wgAuub1xIRRe8zZErDfd4zxJAdFaFsOxakPPCngjv5LZVSNW48Sz4B
yFTWF2nYHdQJD+3v9bRQM1UM6LntSx5vlxNzoTVpSEBNUZMrKE0iAmP4vreEswWQTbGl4b1jb/c3
tNLBVbXBpHNEiWOZ1LHIKKSsQdt30SQHQqT4GTPbVepw1X8Haw+Fq+nLUmawaFCGz+iw45aPz/Tm
keojMyS+tRUnRJMwrva8rtVQY5D2qzTRbGl/Ku1Ur21l3q4yy8+RJYXlwjPLpoh6oBL9kCeUep33
47uQUwc9lumVSCvQlMncpQtUyc2MLZvYYRULmw7i8GKBXP+75R2NCJpRyrjeKvH7rQ4bRfjuVQOM
JCHL2R8gh48EryldcF8nwxDtzscdK84Egtg/ShxGxOQJBBXyECL7PcCKxEnytLEpfOJcyVCk0CW+
vlByFDM0HflB8cscwb0vTlMHwRiq+6jNOlgzUf99OEz9W08wIzw8BMljpaBivszN0n7pJe2WuL3H
OkxdGFCsLuux5jGZ+VMkx+koFm2aSFxDwKb5nLK6xUwphSuk9LcZQdjA0fjt/7DcFbv/np36EV0G
WOii+gQhArQATNWjR0rTycrfWru4BeVR7rwGn5QCiOZES0nBgUsFd6FpJ/sbOxB1l/ez7038lwx7
Epc1nTb+zj5p5A/Y7G9VrcEvDleofD5114HbR2zYulxGlhqsj3YAtNX77nIgJ82G25f6PIPbDyxb
epzn2aqYYAQELpZIPlmleNeOwChqhen1dfI6mXkgenPjgYlkZCwAVsPiJZvEZIJzaa/7IJT2ag0q
0VTkh4nqgVEj5Q4tEGmjUX0ZfqOZMNE9kdEGSlmS40dQedUkHLjUagXYf95gPcKc2Mr5qWL5OorZ
YEJ1ofVeIqNxnyCjni5KNlTGtOPSK+8QyXbuUC0ftEVaywYc9nF/tPGt+tUMPQ3skavUS1uiQlT9
5Q38rR7oMhBvL/vbjlqBNs6yfxYE6eWAdUFsjLJSI5twIoIyn4jdCMlcMLopKk1v1p9+uSbYToD/
asYthZ84e1dex7Ujipq5XhNSamkKOcIz0IEyU7YpqqRpyVSZ5S7mJ8WKyzEw6FUpUrvo4jxGSGG9
C2rgSRY8sQnNVFspUDPl9PbuS+UKlx0iQS8KI75NgeuGnAs1esxkhuU5jLyx9m5xHXeLXaQZCAXJ
wdx2MjTqELGbxSyoN5JvK5jlWzmlreGmSIzWT1CqwXbSJLudf5MKwfwPc9ws54y24yUpOnRjuaEF
KJdicYnKgkn5JMRaRP5X4BXTXFVtC7vtRzvNDxaCI6jCOTNAC6QRbWSbGttJ+uqBLbf3f2uAOHqI
3VGVweUijLp3xH+Bj50b6G0or3g4LHvb4n99mLz+i+5DytSOcuHb7q5YQzpexDZHEpDVfSmaPv5G
jjIuKDM1mgSX4jjy3e+ij4+0ATcupPRZOa5ROLVkdun9Ni2DT362XE1NZeEeMCYKJVM3SVLKb05D
vhUJlGfCmy7w6N08G3B6LGq9Vq5c2X9de4NOxS0mcvs22VEaFaeLBXNse5qwYG57GVCy2k/Z92vh
qfcY+yVdqV4IJTYdUwQYfEhMfhIusgsQ/C2U7rrACOK3mT1gCREUSWuhO7T3dD3Mr5kbIAdph+uZ
6VJk+coMJdhcbcX1kyEnS+OySv7GG3lXyvSxDfXS1m5Nz12/GeMNl1O6N3NgBNHmT9qxX33roBrw
9pVWNU3AhbMYITBVZFCZzWnD8DfG367kcp2hLKxCp1P5xCoyo/AyTHrhZ4r705bRPSdk/2QtpROU
2kXUjqP3i/213JX7VwssqKtXMn75PF/RpH9/SmQ5re48Mk5OYBAT0ADJPY2y5SohHIE8O+eKThGf
isPUfFmPDKL3YTiDcYQGIhmtdZhpUFr7sxPLFDgD1LTfBnmIsvH9Sjo9YQLfsqmk+dRAtLc4XPsW
KMaR+Sn+VsnH2+cz0cv77DX2aql6JrFo85mqE6Yb0xmde9GltPPs/56hnt6p8C+5Zc5GZFrUXXSl
kQafQz/H3d0dacZNFjyL4QXJhY6n9ZGERt8+9Bg6pF7kleNSFd+THVorzS5AxbnSm1AdtzAQVK0l
7gb9z7BU4uvI4fSbP1x+ty/xR55wj6HnkhXSfIE63HHL1FqoFnv/ij9CFfAX+N6x3HVcqiSCPXdR
qmEe272k7sggj+4FXVYWziK2mbt5F/MB7Yiqy10XyzAuioqbkdDsvL3aMFmbjmqK3mQ7zHMLQf3W
QOBy4yDnXvOrdkUSmkGaS4NkPKGJUkJlQ2Dmno6hckPTCZtZIJZ/nQNe/nTIxsJjiZYKm7zIwn9F
/j9n95QsR3wYH4gAZEN+iYREYtlh4QrcXLBmj9kJyNFTEaXnljN3ByYEsjHvbN4GTt6CQCOx1Lgg
n34qqykHDV3M8a4nkT/iZM1tCJWCMOHrrNWsSn385kcjHGIlDStQ7BC/W1O+gg3BGbQ+yc22+efC
nJlUAuMKD5Ufs2egT0BbeV/gGkUhZvNnd/oz/gfAqgv5eIHu4cyLKQKI7Q3APSSA7PygaMU44GGl
DdFMjZaPLLLzXXfjYOHvixMAULFTQ1ZVHGpw1QAwM/WiOT9S/120PkHEgB/EXHZ5Y3C06EseRBeE
xnyntztNDTFcnD5uGmpTqeDN8vXkLIODBxiF+zOVSCyjjVslUm8KRoE2Idv2MH7AcJl+AUJ/fOiw
EYRM0ZEt+9vK6cc+193HDpb7t/NSx/JTWlTdzRI8FGwX6jZdnOZd53rbK06VIfHTsopWk0imQhWr
eHfy14NJ/eH44KMxW7XLVqFScVU/GngVMFBSe68IoROFvJrXNw+xRbA0EKcvYRjnlbzaKtkWZ3p8
JW/gH1ZifsNGeD2s/Hj2AA+BstZBuQueLa91zCUpIhxmfVyvEG4u/CswLfngDKNBguahG+R6KTTt
iXi/vN0GqwP9/HIh8K+sMfweGa7Bne6l8nP+6vxpSxw/5CqcJAj4GPbPdEpgPL56nnkUBpLhm7nD
yZ135fSqMbAlA1ul9nTHDl5jcNPJnRfzr0QWQ3GDYT4KMPm7lWFjgXJllpGPAtY2W3GMiQQ7Spub
jMiB270jzkRbqg7NL/nnjzfLRRWnVRitzYCJkZgtmDMXu3J0SJwy96YEmrQg+mUW0X0zbuXoJvt5
0VpYgUaMHx1tNX8elapS3FfoiL+mINClyBnUBlbHnC7/jxwuMYRuOnP8oW+aExHrJXNyqZz9yvH6
zvu0/2Y/L8g+SBFhomJMfj6AA1TZupc/Bit+hVkwaaS97yGbtTOJmdVsMNPMn6OF37V0c4lzxPHl
fCeyelIq/tHq+rO3KP25O4OGNhKiDVLlTMuOZyRo3KISCu9qn3o0g6q1XGY+9AedL3OdV8Q+ZbRi
QhlToGQUel0Q6GcXBeCAXRUIAP3lLSwnXeEQHc0F8ZSSTszLqMYaTqSUudwewuqvL4Lj4byxNYE/
LAgkP+3IkZyDTatshD70Ny+x6KwKaAiCI5YwjROLH6/SyPPZ8MW3EXG7fi6hzsJ4/Yfy5IOLiU0w
7oJSCqM1XfkEX6WCIRVpIz5TZN4qhjN1IuTchXWXdjlvB651JLfMtUkCT+2V1hW6OZLF1WoJzr9/
1DnPaJLP47RtiI1Cb7/OqltWQH47cGwj733gZ6NHuC8/WMHqUHjtKAeThwx9cRkwMtmLB5y3tqeO
ZyQ+hG3O/ysJEeb4nopk9aE/tkaXsEO4u06bujX93cfNgMZkMTdK7VYdvvg0UoI/Zx7Zk8IsCAua
FwZ0u69KdyuudNydpl16a9a4bRM+jp2Jl9GPJKA1Kal2Sucshd80oWTMSHb1AZBtlVYDGL007+d3
D/bnDg5RklP95J+UgnFM2TUHi3uW2k6Iaj2ZC+fstmRvEIW6e/POkGpTbehQFisLyA/xKoSsk9OH
pQpSE9A0xtySirpiExm/a+XCs6zkTl+KQBssCYlUoz5iIpW6Y7j2fsv6Xh6rwvJnvsWveerqHUaO
r5WY9q4LtM5/ITIKK7vD9EPf7HVZA5bX58qY+8TKOlOZMkJP58wmTQj3F9o2bgvyjK45i2yOjJhT
+MreA0DkbAQKACyn4pQ8rsnEw58norq7RDL7AfGDsS05aDgh0QcKxzRZCXUMhJ6+BunT5b5T3B+l
//02HX7GGvfe5qYbT6L1aDxgVaM+q8NQrWl9gOGyhiN4DcMLr5fiAEgRFbSiQoIn1ZpoFyEUDKo0
4oj1FGE1TN/LaKbLGuNmzA7SM1SkcBA088MFIYgRyQKkdNVbjCV1xqYySMeD/sLxOfnYhwiGufOx
fm5Jjxk9LZohA15KF6qnrH0fgr/e1p955w+YYkbNoMyhP0+gdt9p1eGilMIHMmL4rRFF59yE30MY
cPyCv0dyaDGMr21IbG77ANcOth/+mwbmsv0ktaMEu3tBDG4+/jeAFazwaho9Bcn+/y3wKuwQoJhc
KJnaZ1nqlJdpceWnB2JnOtfrGujdFLwAW2CkPGfP4mK1MLPRl70OegVBtfTOHSuyaqSWhbIq3nUX
4wAv6pGHyGmhMe6WayeIrEpvcA242ERtLQpZrB0DvamCn+GF/6dEZNTw78KK5wCNQpRui3T9tuR8
qIHKramNke9VvgLvUvSkDcyo/RmdNK0IpQL/w4qFmixsxZeH4jhpPMyTRo7lNrJu1y7UZWBa/Tx/
M6p9Oopuqoy1MwwJfgM2hNKBBMdTlybPXJLM/4sNlPc96Kv/SFi8aQZX+vYqZItkS8j8VvsGFECC
rjBu+oQzes1+DqHdOl4uVh9QcsHTAL6hJ/FSAecdOjBTvfnuS18h8kYBpcinDdgTuLB8u8cQhFkO
WhM2dScu6rO82Ok2nucAwyqzRlHDOlQJUjFe2NthbphOveJA5ERh1Jv4LcXmDA/h6UMSjjrCjCmU
qfh1/2mTCcQrtnlMY6T/72F6vTBkB/6C7ccYSUTeWOzIDFJi7ihUz0ZzfW2spduIwPpixYQ5QC9h
GWu2tgBZNkp+8hKFkgWfHgCrH1EfiOsvG6p2o5gIxruitNHO4yJqDScMRcRd/fYcyEih+gMH1Y2s
cPn89qiJvd+o4WNLIuI+o/7T5KxjJToMe5ubhUgJ6/+GTJx1ErQrtVzGonPbvWT6fQ2ssfwthOvv
H3UjLPwWJn+4QmGQ0LAX2MxB2b7xNphPEIOudoEQFVpKcKg5mPlxpIKWOKWv7nG2BJIlNdfZvUe8
qdY5i+cboNzBXiaFISJhtmkLfBK3R6EaqaATmbTOI0Dy43p2+qmTM0yPR1MjHh2XRUea3Y0j8xVR
/RFo+vJwE0J6paBP6wcmBhWlgVbZ8yaGCtl9ZZp4gSo2SBrkka1mALakkRwy82ArOmYfV09GG+c4
cxvoaHNLwP4jrzJFSWNJgYNBdAiwNNsNVIzT6FePMtC148vEpUrzdZTyPigvgEmUWJYijk2+1mSV
rOpBPndbosP7eSP5coXJbVey7BAmRpsURrD32GF7G/YQyKXQRaI+UE6diC2aultqZxy22J8FvDMS
bdCSWlk6VwsSQni9YmE7VpycxbYkqEElmp3Z3izANimZvCXjlIHpZXld0sdauu+Hnuvn1bGvWzKU
0IM0zBel8IXHwI05oz7GJoG2/0tjW3O1rBK6Sk4U0FliOE9iGYUfVpH2kK6HV5QG0tYo0agYkHnh
G6H5aqFw2RCbNiBFraBjXRbtkBbCbWwcz50zHnvFepurSKOBwr0PLe5jZTQH4u7ZeRfR3JujVd/C
YXbqpANL3Q98xkyKF86NRckY+mJGDBR8hmM+pcQQKn1ZtxM5IMkAnmWjX1YMy2ZtPB2A1nIBrxSr
jqXMT4MI5XpzDDLt12706EzqLvzB42wiK7ZdF7SFFmItUMKVWdK5BNw9Szql8qWsC7hiv0kB2pp7
rgAPgqAQnOHua8GF5mICvlRBEH9j1KkYvz0dKl54B9FC/Vp9ePllR5Qubp7DApEay7lAv4qwyCp4
g+PI77fPM0H9Y65BrHzwLRo8+SvPkI9V8fZHwijXXqhZvqItMl+ZOd0ITTadWJeNH5su1Rkf1pED
Q/ORgzkkW0i2+0aPzyep6PBfGuxH27r2DSy0UVZc52ar3WezV+jDj8A64j+k+t0wm9KzpcvZi+fP
9Jd3rXUkzhkKsrHEgtdNjYE1lKCWC6iDsfcQQmp68gBAYoifAWTkMKRxRV0KGBCLgQGvzeZjtfK/
z5ZQdQ+yy5N6mfE0ssu+Zu71Iwz4RbK/vRByFe5XuPopDYRPiQRy2IYpdpOxA0bNE+5qGBCscJdm
BMhecbmTKf3ZYSbWG9XvJ6HRhNuGnvyi+Xpt6mNy7QDJZyfJc5s8axdgb87JSfEftEXJSPEgtlMz
HKFwyfE+kC/0LPJYTjoSgQRll7nN/fqCV05blG9WZ5Gh3T76GXKppqau9TfTGCJMWR7XM6UUsDlz
42+PdQ5rK7Ec+lGc2WiidiiFf1sLXrECxDTIwvFKSDCHPkH8BrClqwOK98Pu7gyWhi2TrcTpuVuO
pE3Ee5/lB3/lQOwDEbP47+jrZVmN+jqz/UEu72Sh9V6+EsA/k8JktVoElQffNAbzZUL+7NBFlfSs
P6ZPbZCDWAyg2qJF3nnHA6ilZqKwdl1qDK//Ig/qFtgRE3BwbTN4UfGEVNFBUQmgf48hAa2ZRIrA
qAoita4asLsttU2+MNLjPyGFHCSyF63u9mWwGYeLbIAtW7y9HoyG/tcJ+c83VuNXCqMVsFtqy8VF
dGL+FvxbUPYnlLY9kQRbWpFM2hsKbUMmHrFLysmdWvSerz67jOt3vC/eqlW7YI71GHQOjzJKZmEp
QvNhJk77n+ue2g1IV0JduCefZTSMnWSX4J8gQEASGEgqPDlkwcZgAAbzrvTEnGjvwitM2xohBtfe
jL+d6gQbqsZZ2mtX0wDLYq3Zd2DRvmGUgdALSzKLykzTIQ4l7RMBH3vlcbaTMek6n72zo0LQcSvH
J8bghRmyxccE+nD6XEmC9CKuwvvVlbq6xyPc03/MVJWNGhZ9q2iVC1RTnjncR4CrsbgmsmAqrJ5w
hYtKksC/Rh16CTpYCYWmEhRpCsQ4ttH1aQ+NRRsJGXeXOkl9klLqq0BJdmCk0XEAlEhpFELPJNGf
W5wLIQVdWsJMTTq9gBDXNQvgbKmVZawSzLvKIYyLVuqwCBy5H6xWRivb6nRhSKvto9fmguOUbjli
sxYVtLlsw4P0MdhPhRK/gGX4Jle9gt5TPjhLHhSdkZeqbW3kR5wKY9beDsp0xfqYqpMFgLnUTvAE
V2vkxU5Xi8kwqRnc/Zga7qIu7HDOCGuDEajseZag3p0zOX0kGi+fyor22wqFIR3xOBrCO+VJyKHr
CmybVWTNJyCijcH1Y30WagbZGGwkBGJyd/fBw27cIgZ3drW18tWWOa3yVEvZhnoik2JT8RftRhXq
k0ogMdB7d4Vq5tohErwaV7wQWn3YkOG0JMxllA6caZc6nPmJXegu1df7Et+VpQ63dGeDHGgPBDkh
ZgdF1bCKabLj3HPE1+Qu4X8FWiNUmQAQH3fuduihE88SD2y5n2a0cjIh8bHj67cB3/cw++rI5nAG
jG83YhWWnrpphZeh9VerNMZ9BuPwRWXlBiBinP79KrwF2Q3FDN5gfdiRb0Kiryww/Q+/iXksJ2Eu
B0x8+MViUuiS41SLhCo+Q3dbueUQ8sDQ8YTN00x1IAFC7FmyX1u4VoVjdZL4PMIz1dtkG9fea+bN
UrgzbHRFNpbORWMhwcNdz2LDwukWY0V+svvdQMYpPUysMpxdUupZVG27p4VFKvzSpkMkMkWx1wjY
t98I2DEfGH42Ta1GsIgIO0ljk7E6hPvWDC1q9Cwbiv2eabGE4Fnm98sIeONeKJfg7eOOjNCL2wPC
mO/2FsD1/YTAbVnjEhp1YnsXSeddoLu3Er56LpO7c3jite2gQpXWPEqtWb3srxAhvxUt7RQ4C5iR
pEn60uOPcr4MtaycM5O5f0jfJxgflfwILiRNZ0DXQ5dINTlf7HAgsX4jCGjIiaWxhigP1Y4Zj9Du
1jr1yXK2MdLckaiuHuQKzQAikDHG8pYZ6Px8Du/JVQ2ClL4bSwVGoov4E1F/9e+Jzwcbe4J3EtEH
dLoVf0pbgP8l6eOjsmkbcG0RnijH/k8dRYjbMe6S+YIkqSjEb5CDjEwvbu4BIljZ1CWU5VFcrBNr
ToxFyDyXz6zhJmpR53pyTkixMgZky+pWupEBXiajGQOg11kFejVLZPkWZnq2C/zDL56pxFPHl/zG
ehIS4KMCgAa1eXp/b9M3aM/6nsbuVoquZVPX96MholR5Jn2sFhG+C4KZ/K0ElMEr+WQ08t6+uz2w
YFtcJMNJfYgov/auDFP/TBmzPjucfid8SgyNIKv+58jgwx9o4uJWy9keeoDS01XmYxxHfYxv9zjw
h3A//jBnB11KtHPP3BpPlHiBsqItcqOkqGxSgdeNo0CBX4T3wmzRCwdk7iitQlMk6arcLVgwyujz
MW6aagYXMZa+HwETNBNFE36g+XKcD4NmX+ixSy3Cn5YkSStQNh17yZ4+ob27BbfsYBe1k4j8tMgf
RGxN0umJw+maetyv4w2e7wr1DbAwMmcTFE5lFMdLSyeGfVFxeLLAOBy3j8t3kG/7LftgyHiIr/Jm
y93aBfZbThOC1p6huJ0MXF0G38HgmCr73d3frUjbwABvVk39ojYX0itxx94w3Si9kSgw4IRdKCWd
mkBwGBU0p4hu4AdaqDeXodRRg+ZbAw0ivnbbH+EPtBv0512CLT9pVLspqs7ny3Lz6xCMctzJmh3x
FR3KtZ2sGUo5dG6sIEeA5xSY/cUb41yND89vxZtaxceL9PIcTys79Rw2wR2EJfxu7TsA4M0GPKUe
5h45zMH4thjzVHP5IFYfAv+0OJkjq/u6AUJG5KaYaMBF5p58Of3rJA2fpLoME+wE22yXQ/CqxJsO
iciCQYYwRt5ut0tnlGljj74CwU/dYoAtax9TXmNvnR5n6AknMV66RwPjtz/2slYBFxneVt0igE6r
l9iTBgRU/klkbxWrWg6DPvhRxbBt6VU5qR0a/tHoCObMbd0CGn9/EpDH3gerXAXfOi9YU5sFWBPc
mWLPO7ej2KIcI6ypLAU5s9Yus7ZoqyjqOP4KdlXaHldQe6N7PI4JRDpiwR5YHc551llLL5frX7ZJ
VEH3L1QfO1s3Yl8/90WgAYiokpTYgHKsMkpYLGUdB8EjuN+UBpKpKpylAWDNGbZrbxt0nLFz7qVb
q1m4R1uFtIJhperwCMXqJCdANK1TJg7PHkplCVnzjlMndfNcTOe/l9pllI7peuAVplLMThKGjx/e
+ye1nIy7Edfp1ajCJ4KKIgRSUQg5qwZ1J0/V3vRGiqiri0f5VBTDXa40580uKWhREKoQqWwnLi26
Kr5q7vxm/bWLLf5BNvDiiYhMP+L1uHv2ELkO2jv8xXc2IhIYDWoSpKgVmakeDlMZGoRBDTjoYXLf
sGtQ7SvKKVzGb2VFjKqBlFS6DqKT5sPY8a12n/sZE+2RD6U2LLQx3xse/3U7sf0+omcFitC6aGMb
c6N7o6SncFDI3GLTyB1bDuyBPwyOSkSrIPzwsWXXhcru59vKeosoM6BIFhzQP9toEEM+BMJfFJbO
DTQ1xCOD3YVTyVBGDwk2/Lgpopjd8MPCVdLQ+BpsA5x0eCyDmozAwmc3cC/+8PGe0ZhkGPJRHWAA
XoZ9WgOJyt4Xe7zPHczKDumO0WPpf+mUDqyJVGR5B4l/W0eDISQA3Xs/kczH/isiGQsBgLp6fy9I
RS+go+ldOeDY+rPUeFCkq6jx0e2F41v6YWUBfci29ESjeqXQCibupowL6JZPqTWPh+ggnolmDmTz
cLS7Qj9ZyC3E+iosdPaQynstRXZHFIQDWvM67meclxdPXvxesMHl2jcfAw3kyM6JBElzzbqXKnvo
JPyn+RJt3ppbpZD6ZY8MlIytLy9/SbxjX1jZgqpkQZsrXCP4v2Ls82rY9iOz+/dWqkuHn6J/bhdu
db2MeRr11/QJDMtM+Pw9u1Z7nJhksgwJV/9AKLnOcAcsrvwl92LZHBkMJ7xa93EwS2874HkIjSC+
+8XtbWtIduL6zrxiqseUC0Eose7TrvoTt+pCFADw+kCQ7EbcGW4j8bmLNhkHVthaNnM0riMc7vo4
rrcrpgV+OaeJ5VIT5dX371SCgz96XbQPxhcuitxZljJ+iPhIST2eQqNyF0kRXCrRJF72xaLzIcrp
CfJyFbrLftleV/XKp1sq8/CCGjEUxerCiBiGYc5lxv8IF0n7Aw3ST3wlIoLi2Nbw8b40shlPlJbh
mN/keDZKotZG3h9XsQ0ozMXJUFS/a8SUKZruQfXnTRkxgwmQsBfoPcMaOYIfh018rJZqk6+aqK6l
I8L8AFBVRUcw9W/joVWNxS92WIzISjaJVWqzSmmIAXsOv2vrylGH3hSSm3pDaBzhV1/7ibq8UkDR
ckgzP65hhMUALk9Y9QgxTJnGzHTxMhzdahO39YN1JIZI4NCpM7ohLc83QavYJ8M4bnC3dvQITu90
vfV985JMtPG6crIjg+C0E1sXF41P/IZwpgOUb6TxesRI2pl2VGUavsm4ZThD5OBy5zMFdiL9JYrs
3iYKpySiAnigbFkgu4UJBwhEaLLrwZm1bzkKGTdvChoSvhMCHrsKDibbLOAHN+ACWq34puNa8RTg
bLbpBKv8Z7OEfECcqZwcfbSEWcDh5aKoBo8FKfTxYyiuwxNi/cZ6bUFbN9RZapf8ixvjnhUcfIed
7xzzk4W6sV+G8iZvtP1zYUAEu+gf1xMh8ycmA7/K9NzeTd3KN8kb1I+ynMpVVlfPTvOer3eNPTAn
qYspGr/ECtkTxDa2CC9LHGtUIQxjYMdV9wEDyuyLixnoSpGXWqpwQt7J3HiaCn9JwxuQfOc86DN+
xhfT7zYXOuqtZgfWwHLP3CvNmue4s1iLUfulUzZ/YlQA+RV6NGuCsIb8T+BwsZW6onMz1j0qAXGA
HNZBSasMZjbktnbyW+NtFwRwnq0HOyTQRR1tNF1MfboYjiUMs0sfk3HKIKq+/9f3GsT5cHDc+uuc
0jPYie3+2Ap3iM0oiutAuWW4SOyVELz4y0F+b5N2pUzDzCP8OllIOmgmc/n6qyzH73i+AtqyYPOS
+uRaK+Qf6wjkOFYovtzB2dEmena3xjgYDbeUKxswL6yE0n+nlEoL/tVYs9DfbIqk9yBEmdTrNWOa
AHdBFqCz7QAIbKDoFL3W5Lwy8Aa0vXnFy07hXX46R1qiac/H7yRVE0qKnRKB4hfk+RPO0kHQbvm8
wYOvT99ohHswSLR18qHsFnsKEiaS/o3onyqLwoVIdG2990+LeDpOkvZn+JzbcD/W4E83m1bEeCWW
ONYIeOquMIXHOMxNZNTTLYMlWCj2C3c4HeydUQFWCABooPThYj8noiOptjFvA/iRRQlBjwoTmH+K
P7iOiAHTI793eOq1YAzBCblQP7sEcj6orJ4k77hE0szucVqhAhOJ3wNI0YtWVd6lnOQg3bJRWXPo
CknSwh+NejPIhbtKFtzhLDDXUhIw8LDXTRYpENEg/cydkyhYEYfNpyiGmWvMkVrgUqyacxSU9yWZ
YE+/huxljYsJ2cWWuLm3deXUPs1SLtiaEFehDpRSbk7Vka8qZk8r7p7XJDwWvWQAYtVXLAYBskYq
1J6SRV+Cxn+AhArg/MXyDKN3z5XxGyj+53dwL6YjNDkmO3o6brUr+6QQ8a4vz6InOyKKiq5X34h7
qnIoY5tBNnpBMYuBfOA8gyuLAL5wWPmMMOektSDcUBqt9U2CRMRfDHk3GA/X49aJyi/Ia55B5yZE
lN8yAXXCpf3U8iOmngmrDFHvTBnbmRGdshLM2rfoIkrKD0ZxPgpM0tomvUiKjfjRATIHFNVoNbFK
wuAGmaIz5taYvD7QEVeT3ntFyhohpYSUC4MD+orX5ToOu+9BpTHVyelJWNiIXxHpCB7WGe36Krzg
7DPzgWEeiznTBbTZkc/MnL9GvC3TKt0c2QehGAJj3c3fH5ok0qu7NtiXTQERdYzvTcmfy60NcpL+
Hka8OC1tNeuBIjnXjUWCVrEU3M0trBR0Ked6SqjfshcurgDibXR2FQKgY2x/OrJECtOOEGAzxFU7
Y0aK1JZh0YnoEuWWEbiq7bDHdfkkSPfSjDLBc10h4WzLumtv5ZeyRTf2QF6AGVFf09rMKNxOCFCd
rPQH6DL+vfB4M4RvMJUgQLMRqYIJXxyIZpX9giTvLA1yWLh7pJlX10XBOcbD38mFAFrBX9ot5kS4
FNQ2NCJ9A/N1gW9XTP0pFXR1OD0z9EP+NT8BjOuOlu44RlP+Rwc6+6WaH2Zt8/wFkel1s+b4XU+8
MMx/GaW1lhbZEwhdw3MsCMksVb4M8/CbvP1ZIqfeGD5B1P1oeDwmcCJL0x2UutRxhvC3bT3H94L1
FDHpQgCRc4PtWW54PuGUaey0FNnUtRR1N6i35B/sM7IxPRMR9JIFMQc4+a2IqdqvzIUluuQXMtr/
lV0poo8YsrYpA0Mnzm1PLkCZAsbMlm7rPNcCIWCoGkwAZlNb8RRyT/wt3pRuGyXa4l+B9AyUUs9s
JABkSbiX8ol6KZ7bXZjzviczNOb1uS+y1pj9iQQuXPJxKdJWHC2ACycdg13D8dvOQDkrEiQh0HqF
6TEbp2qht0nTjd363ZBrf867PcIej/+eLMT6KUu+Og5xPa/RnTnuq0ayg1tv9TYNCvbikvip+rJg
k1fMfHX66FW0fUDTTQN5hNvAxgZ9K8egyugcw6GrmaAD8Enp1fCsNgQMGl5X7E9qGgoPPkZg1ZXF
9XvGwhxJfrZj0977rcfW9m2GwunRM4/wu0zYU+0GIZb0DWCIqz8StEKUEgREpgK9LsjLaFPGTnXZ
v50uDUVt5fURjF4RrBTTTnNIsfmi0lu+P5K/lKp2nXxwuSxrO5LtJ/Es4NLRtwjJrYtJmcyIgrTK
/nfmmS73nxz2uYLuvb2n2rDCPwHy2G/SI4dYEPXYxCDhwLT62C0YOyRbRhApaNG0uH9QTJ26/fHF
N+mjaNZlKVDsUa13oaDUEEydpKBxX1k5tU/H16+InSOdfH6hqeGp/TRSQT3WfL/J4JgTmFZI1Usr
t489E/dHPDWo4NW4Mt1Z8O0Tp4yfveD/w85OROadbf9O1ork8I7X8kSzIox4ER/s4pknDHLCHtSY
q/Lig6Igl6mGz+VbO89GdAAzIE2ngGNOUjyQ6rfOfCVPH5Fa1wgbU4tgfIUV5VG4zq6SaOv5QxAo
fFYUslo0vaEbfRTCavQEdG5BoEQ04Q5F+6qo30pjOqerTYbo7+gVhaUUQvdw3cEhFD6ZqPJYwQqe
7JNaQzzAKf7hltlHJ/XWiLhqC03lkk/lgf7PMHK0vVHftQCVoa8XKpYkw7nILroN6OkD7+1hP3w0
B/HtJacPyW3kL1UTOro0vpkvbFHzzCI4McwhetGhXfs/rJpxf+VHpEReM8OK1+4G3JJFPTlLggj1
k/Q79UNvpAN3fXMe4kUjAGnWzEdy8esfK4i50epYYF/I3ZvXKHBza/aNtlUbarDNWNlXbLXG7OIt
mR4OWx3o189k4r//WUTnpJtnf2SPcZImaDCzXkhq7kkAdEI1N4iIgCanJjCaXwy5mtOEbT+cD8UE
iPd9OlyuOTBwC7BsJe2KTZFIGTpsqSF15HSJn5grSvL5k+hvtHoxzzspOoDBxsLHQAfKEXfD+efI
kZVRRFuvBUsqaakr4HYTJk2/WOBQNHN8K9K5u/i6dYkgYxwYLN2OY7XrPoeKZzKS2I2PV52T6YOA
BZP/Ex7FfVunf910ezUBpFAJNs0Omy6FO34K9w5LmFixtZ4lsC64CD67LL9yzPDg/2jo+D3vofTg
tP3TgtDtzHbcEJpYqcNk4+smo0HNyVQlEJuaQYflDReftFIkbEOBpvKJaV1gKZtKus1/ifq0bOCx
ikXI+JdEUzy+3P41AwIsGEElV1QfOK8x8aQnoZgLUklgoCjD2TG+QPI8QCxB0l6X2e2sVKDJt5FS
xTRUt8Xetf4LGNGGyWUztZmlmHjEHn9wp2FzQnd7B94SvTKxpHiQ6bihvpWTMplvSik+ObYs/ozu
OC1Jg4YdVUPnFWug6i/l6hVootjOMrWRTQhOQ9JTtO3pSLDn09VHyJNqIg/RJBAysWFMtHUgk4gO
3ksDZKw3TC2wpD70fSnyKthMycBiALFVlGDyGPbjqSxKQG2mrhY77Rx3E5AHqgdIVHCJblkkkGJz
GKn0z+d8LXgEpyQ904rQpadUkfykTTGExykg8FUoDtr/E6NAvj2sLCMl20xLdiNV8Nb7odjkxhlW
snqqMSMSI9PX7PBSc4m3BvtLKgQK7QmrvmEBL4KaX7/sO77XbMeXxrbW1FOW8IaXisV5wO5Zvp6k
rq9y3N43K6OUuvXF8mTdBKlajNBVLy2CIyhSHVqNQxQv9izzExjgrWVGbzbFKOgAuqyoQ6FOoNxT
di0BT0Qo7t2MlHtf0H8AOCqmBo2q4R/Bqi/p9wGnjPBEVQotEeUm5HiuRZZyyILnxy2ULqMIP9xB
cgsdP+GIjxVlr9YN7T4no9PXutqnaO1iJ7KFY7poJJvLfbdlFVflAS4CXhZUxFxH7Bj4x5GZd9qF
AS0tmdnmqZaVRTiuIX+CakFtsFs/POUxFuzLYratxlFUlAB3TKrrueJiaSbh/zmiVeO/8+8r6EUE
mQgEWKet0hidOHCkUP9igwsB3ZcOEyXCZEHCF+p7vSEnvsqhQ2lhDVIf9BQU56enn5O7+M4R1Sue
kBEAv4QOaMEcNFd3T+/9u957YKnfrsTUouqGE+vnmczynubME2c2dVBONydgJ6uNZewj/vZdb6X3
4kXtSDfhPOlPs/4ULdpM5ynwoS38e+Rk2U6eKVscq9YX/rPb6kWdwTq01Hdje257lEy9g0PlUdDM
rTIeEHV/CVoWhWc3rTgkYxGwHKyBDuaFTir4QKdVltqUTl/zvZgYKFcUVg01OpFQzICwSxeXZxd8
BgFnIWBu7lBj7xNb1nOSONvNOJBaaBwb+YhgAX3JvGMFa0F1x/4YsSAeRAC9ZAUJc95f1X9tV1sB
2wEX0roQPhNZCg0PpNXDk7rezhCiJGU5j25zXwG9qyvAb6e/EwfNSLwJVXZx2ykipJ+4mG3wvQsF
S3Rj7cBXhsf3/93d2C9dH1Z9dFUK7olD/yyrxwfCQG9AhjB8a/Td2rSbW7vB5ShKLaeoYewbvWYp
EwCZx0aaurj6i8TbnT5gY60rbe+NKVLygHywZp9GwjF/O2noL2XlanTv90B8gZGdAmExgmr4rkMy
uu0+v4+vjGTt0+Ht4PPvKJW7F8nYWV48iuSszVZNOR4OW6L4NVQ2Ab+6sm40egWYqcmtBmNIq0ev
L/xLJXo89QfInGSTbGSMqxRux1/2tfjG05Cin3acLiNbaGjt7LPyvd2hdBzF+s/1+o2x/JKKakM+
w3igzUxvO42cWz0O2bnI94RA3LetuDlH51PejpyaXCo6+czze5NuX7HVtVNvrtxFGoDpFt5rZXL3
XhKdQ2dc2JTaqMAe9gxoH0J27Iiqr6QHSa/VDx016gyHQsuWWMAzC4hNPosL/AR9/PSwUu3uFFsG
/1XYVpYX0rIq7wThh3aSEj4hEjyzC6mmFSAwpP/QMPmefYQsnSWPKvxRg2vkPpsCFRt1Vo2g9FON
htcliCVAtH7dI1SRI41SGZN9IV9ypCmN6rtDdSWorocDfNBQ3HIScAFb/MbuI7idt1qEmAlN6xoS
vZFaHq56LTqU4dkdHku5bsQDHPV6CMLhYeVf0p4o2ua3TPSt9BBvz42K4R8GQYnevjVadF43SrEn
LuJn3Ha6lITEj3xqqesU6N7RmQu7U1xW51ETYQ6Ya9KGg+ksjWsVmnMMyZZwjAZhyUJwf5mv9bTc
vQMzZvu/ketEH8RARBtsWMylFFLge0IcA7dYl4QfjZSuFHK0u4vnycxOOZoXt8k/ERQzd2pEtGv/
QEZkdOgfVuYYYm2vgHra5Y7LuFs64ePKFmvBKOSVVsVh+qiXcvBWmzhDSt+EpT79V0C66mkIYyas
f5Z10+jQ/Q7GnTcZajdFgzoUcbAXA3qPJKt47ncToeUjV9/eh2OGvNxEBw4qGVHZo7XA7N5QX78N
0c6HGJKDcL6UzzhLQTPHljXTqGaUsLUeFbubqYnwuv+ges/H43G1repRLHD9p8ncEextEvdRBXpq
dFqydM1YyNrZum5uUimmsHrghoOvxs+JpaFCXS9+YWeNOgeLGRbYnjerBXP5HS38+aHknrSfgquU
w2cFDYSoHBkDAlVvOwWIDoB7xmhwK7yXk73pTfkw3OR3/sfwxBrJ+TBkzMZ37XK1ElK/uVfMfm+v
MnCZBOeJAEB9n791viu494nDmt6V/Y51GpiHRWiWilbBNpDyjtgjCZudHOXSqNQweYeuz85De54M
qGbY4sJD9Gz3Zg/wE8U/w6zzaRRVuG1vSyA2QQGXb2bx1+ZUIErgDjGUhEb+IqOj/00KJfeyD1He
zs2jonTJibc+0yWe6ri2kTRH97Ro2QSkuK+nLWxhfJ/Phnk4KzcXE0aebLJ61V9GYuxxyaUkhWGQ
5bBvp6xY45PA7CRayDpP9fzP8M1lb9121yhsq8s7jvTAHsSATUJTQ6r68IfxlVsn9XL1fckgmvIZ
MPx/tKMEGRUoM/L7/7O28FpzyfwNMqeGd/1XUgtTRSrluMi6sILIXOrPvfPpK3Zw3IkgAyOw3lYP
yvBd7SyBmPAVFjOgcCX213aHFT0HCSlMPGESlJ+F2amcW5wT64tqEwZr/OOfpVX3Pa+g3zaTZVuR
VUeq2491bXggfGDM6Qzhd3ZAjB0dsTZKp+sVERiEgCW3WLPsL9Vygq6XC+pXEVWDp3TBwKhhEAQ8
YyWdO15O3RU7zI69ngqOlMjFEmMQZZhJK02lfFiMqgZLIK9NsugdLKtp4qiq/j9C2srxeU3HcHfo
7yUPgDm6xLuUhFT4hSbfvVQFG1rgzARJeS+ZTNyt7ZofbPhmz4SqlVTRcLHxCUqud/JPC8KEu+hm
GrDWt5cLDFWEXKeZ8voY9s633cuIPRTkJ/ZITXiqBJ9IcfwdJbBABoy61wX2DQ6jp1bepNoCsJ8i
yKhclu9Fg3/sZQHsfJvKEaZZXaP0pl1/ElvVLWaHzhFS4f8Plui5QkN9QPKCIldz1hK2ZV/982hW
Ogtk8DHpn9d81BtDu1ocvCpyYTwaoIjbaq3ZO/+o2KiVKoo6AeTyFlrgkdTCYY+fhe8oXgasXlkT
za5ajtdt6Pp/dYH8gkH/t9zTWFQK3yoVzz+avDycYWdNOOFP/vmfYw7W0p5GWEx4cWLxE8OiiHUS
ViHbaUWF7xq/5H/B91JtzLBbmjJhy3IwFnM90m/ikLSn9T8tQmmmHqVHoWDPWLsnFpstSalEX5HH
xl8QcLTtf99epfEgpOoPrN9r/4u+3RbuBbJketiBi/LPxCFezZ1l/ulb0V+8kChMSUJoDya5pf3O
vHBSrZ+SFp0OFs7pZXqlLhu0tIbdIk7+m+TJAOEjbc+Y5sHXmW1jsxqJXzOA99+231y1EQTZaQPe
iPv5BT4bduq7mrSezcLfysbxMexTJXftIZPp+ZSOla5oSiScxNF8t2Jg5++BrHp7hUJorrVj0QoI
ODlNp+fdIb+B/hLJfUpMP/3lF1+s3sPYuz5D3b750YQnrMBLpuBbNEK7fhyLc6lGFGeVQDn2Eii+
p1itPEgq02CmGosUWWcSxflCHEhS4y5J7eFB3ILrH82QIaENSYQwYDq+YzW+mS7kA1MiKJvFt0U9
ok/jJmAMP+0tFTM+MmxVTrnVvPXXkjH95aiNLnfhj+iYej0ZazeI8hJDrwygUxgeF5hii4IkOM51
xtETgsvVLxHS1Wz4/vvlJ2s0SH6bHRhBZ1KcRRTRW1GVRKJK826NR+giEKSJd6m5MiZ86Hogphs5
VuEmDLx7+Jspo/07sG/1pkMn+1WYHTRugtP1XNG27pcg1GuyA4C+5j/Xog3dD8sJNAQkZwvEpe1r
ZYmo35GBNGVrfu5Sv7yieGcPnMImp3tz4inhc9iqd9gV+uXToXILxr1pbUHOEi2bZ06Us2w8YGu1
qtceaphK4k2r/p+R+1HjLYp/BIzK4WnUImdJouTDWCgTSWJKSLrFg15V3Uhj5FDsm3eDppnOgS1U
jN7ctb2Yi1jM8PCs4UwypXrlM2ChU4t6vwqY1zb1kE+AhZDoA5qkh/CIcbeivxsPDfiw/0SkmcsC
3DpuVljuBbZu0gGLEgUp5Cw2B+lg9slH9L2VyVW8NCanMjqN8Jnl0kfodE8nbj1IrRvnfkZajzvt
Abks+9jk2GHmz7OExRYgjPcT5VHCbMJxVYaeDjU4BfnIN/7c6bIga8VoczaRxspEWp746IkOPH10
fH3ibwTm5HtCPK4eP64Zc9pKAdK+aP85/obQk+I3GuAzhG3YSqVZb47X3LnFfmOzBnynuqhdexH7
pW2xHoOqAYcZnkhxxRahrwyQadUtUyErFONoh1Jd3P9ayKeeM3mZOQjxwCwhacCd00cVHmuWfo8p
T7wsr939XauSxn7t3UuHRCMr+FPsfxRCTjNjQAgei09BmOwQslfMkHfiL/mCmUWPy4VtZjj0vTeD
YiCc8sYFMNhmq2zGoQAPUyaAuo/VaIT/S/65BugNwEV59lKvvlaUV5mUdBS1lJhI4Gm0I6KgebwV
DkWx9Mq/CO5rwFYl+Ee5/X1Pc8zrf0GJ1plc3y2yMT+Xw5Ydn6Dnj4LZdU4uO4oB0mFa+3yH017K
OjvJdyPH/fNT5jurU/DwuotLSqtNFGjT4RWc2d1NHkZLTQnNgN1riFkSHYE7Y0ReCGWa2w3jSnYZ
nXV2YgID6Ob47k6aocHCeGFQizlktQ4dJ18ut8QWLDJrZ52oD2yusrqaCkFzfBsrPnHUAdfzzLU4
7miLGG+ExmSRieaCmjL2MWfewgrrS3xct1Eyk93jIEKGgJ7ytl+9//SMEl6JJNUjNyj7qZb80X4G
3fmsdsg4s6iwO7FXGJZfX9dmemuoEKk/IFG4qqYTixBacDMqeIz3sMFwAjfaN3rAaF6j8ikCUrYA
iLgZ4X+1z6c5GD2hjZSKFfsbASrj9SpoJdq8U3oPLjwFt/vctdvAz0mEtIaG51gq8GQZoOtDFL4i
4CvjJjUlkfokbRFPHrGIQLqzuCrCO/wNB9bAfeeCrtzT1kNbeFI/ISa78Fden5wq2j3AEoUQHzxg
PYYRMgajTeIE/QD5SjKg6rGovqGxVsM/WLgMFDa45GDHACDRUNDCbGPgbg69n6w8Ewh0aD1OEKx4
DWNJLWIoXRQgbpjTm/VBKuzvXBn5DXNTWYBQ3Y9aWQf6u+5sl/HUaJ3Kp17bNIphb9aX29CISzpk
BDDwD9qAApc47PBN2i2elhYPOcLq13WEmV8PeeZJ6RBb8as0SZFxHmpK68Tn+zZJcohKXkLKeUOx
c0G1Usr4VjNtKo8b488YUqF/FephPxNEWBNDnQX6svJaMzrOzd1BKAWXaQgwdTHa6Avymo6J6knB
IIGPE3vnVrQW+8qSPXVcu9tnhFJI/+D2yVxeXGY0J7qCwjRUshHPxW+FFUHbWed+j4eatWRK7yH3
NqnBRseLuRwklQSyO6KNwvEz7wZbIYjt5mGcYq9yOm6u0GJa8rt2AlnPa/Yo+3S5pT1ruODrYktF
+kCuQj5Ve2AlXoUsNiqT/HPqY1cFrGic4E4q81amPuARmrvgKUCT7MEhD0uE2ZqsxVL23R1d0IOM
6ub1ek8aZBKtQiWyfPM+7N3KLXdhIj3l1ik5vpYgB4+9COK1+k8LlqhT3sotCF7AWXeU0/jlrSmj
pPuaX39wUIJLv3UqvNVY6xJV++QERBLai5zXKTjQmQt9CHP1MPkbCVXPWfO3NalM8O0kgDfp6S0s
tqSIWo6d6EaVAb5PLcmgLKApdTjMmDYitL0AvaY6JMf58SG1zUPukG50clqBV235rjFb3ENr7hWF
h0ctZGGZztsNeOTlAnBppVM5tcSnree9k3F0ZDdN3FhXoZNorYrVXOiw2brkrpA9G9cf/H6ob5q7
V2IQnGhLzBz39OstajHYlWMSJY0myKQMgHkOZhrt0MRjWGQnzKvirPrzTYuQznllyYEwQtDJ0HnK
96K3oS74AJ3ds6PUP4yN0OAN6HFPGJbjWZoyQ/VyLx76kMTDtFf9AynXC/CXd0Q+KQtJjJZaKx5n
P0+8oW3uILwekq1e+E2+y28cQQf1stzAzh2Oxeb+AbwkJE7s2ebRqBiwaNkVRhZ00iR4E2B4gp5r
8IIJpD39yiuVPFMk8OtJiZ59ngdEk6TMsry6yYZYH5HTND1qQ351RpjSNXmW2N6zns3JxXxurXPc
uUjzCHSslSCxMrK8FPod3W90vhKWwXVsygIH1zRooESrV7L+XS519dnc9X2TQX6wriHiHsyZglno
thA43iXPtBHbVE7E01TdqAAU5qfxhIXWIr3DBQsuB/TDyNfUCNH8eRSx4yzACqP1fkGUxBiwHHOO
Ou9AMQ9/Q/672wqsPRKxjm2/ZqGzGmpxcmTU/zk+f92j5z3vet6W8YHMFvJCdq0lwMSGZaIDdDK/
RsABxACgXvcCw9HOtW2iOrckJCd8zSIRNRA4mPT7JhM60sQIxfL4qV52v4Vm//SjM/VdoTH/uowM
NFtuRFUC3e8ajdmxeVMiQkjqtYMSmPyLR0rJLsY3XmYFymMRqRAlDMWrYBfhGrVQ8ABu/LMthEaE
zYaBHBzcn+f4GPNYas9me6tsvViNJHIeRaf7WA1BxFqJkULnSuLug2nwgMN1U7M0G7x1pbZZ6Qug
duyLFxxRCqGV07+NrDHT7Hu29HvYH2LtAAoa8FLRo2HjqkgLmRUZK9FGmRMx3foZGHopDHncSpUx
zBOTxGPBIEJZguz0J3bUD5DJA+8X/mew0LD70eQFcoXpLN+rqHsXXLFfkC5l+zynDwBomBdenb6S
jU+eI6xxNqEfvuaYuOXcs5OWPGg1vVlPmzZSrahvY33r6n+3i6YaWkiJmvhIIwOM8w3Yok3a5Rxt
lY5Di2mS42GgEw0ekbVIFmWHulCKcPzQwpolz3K1gFBVyiO7yL9bqcioUPcrwI3SxMVBffFCWnwK
9jB/maygXqngc2DT7e/s0INCaSx9b7OlPp1QqxY2WwEXt0G+aeQEv/H+Y9n6KFN0MKDRW2JYlyk2
eQjrKOvSv0jqX/5/YSPJ20LBdENxfJm1uo6G2/YVCm4TVT2tytYBp6arEn5ODUWqlhCT1dOFAgfc
ZQNJa8GXIU88vLDeJW9CJwPlBoiFkeGNQq7QXWqxUrsmzLz7CG8D1WqU6L+WM4TcpmQf+cEqZfKI
SFkZLtNx7rLEP/+wN0n5FuBl1m1zlMeqYOEMam7sanPrYJuHJuXa6CVBgcPf3rXsjf6RXJTPB4VT
tkNQTRSlzH4A1lf07Cf1ajk1aOky8SeEjyRsEDCsygFcc6LjuvLnIDMUriCW5qsVs3w5vUxCcGKL
xfiQq22FBb851En2UGVLaaby4jH/lDPynBeEmvBbO4nkb6yJJAajCJ0yybTh6/ue3JKDv24wtZnv
FDVTDg5/0bRzpnGJK04wWTSPMIh6EU4BIMpJtQXnRPeBaVq70dB1qGZH2FVgPkjeo3tyRAL5ylmq
e7G2P0sNuhuysWga3n2s68HeMFXHtKhURcLR50L3m4x9w894QwHSUlKyNbqm0xxHjVuJnEC+/b/m
8SDUA7WfWmaPiAnwBwhZet5nx+4RchNBeEEGX2DhMToyqe9HrRUMf9kA/YC6zRKd9Gg2D648pnFj
r5Gy+8BJAvuwIlEBx6UVyqOZFXXFEhbXu3JgKF6esbp0/ZWvv6bKodeYPgYW1dL0LgRLL/9RX5Jd
eX3ooraH2/r1S0oMkBpHzKrEhb5DayEhtCCmdzhjkli5OzcBJNXIm92QLcXh8VBrr6M/2rVx8vM1
prU7vtUUZHV+ohj/B1xBz6AEm2F/hujd+Z2JVaDPflrrI40e1snUi94tjgryEo4BTuU1iL4H+f58
IntTh39pUyNcUlK8A4HeFE1GxL3tA50/MQHb3mU3400AFF/eOVUicx7JamJkaLxVbR6ZHq5DfBQ9
98diFUpXLB/4HGYp2QpREp2Z5sYXB3p7M76ZWBEKmoEQcPQPunj4DO0+l7BP7uftvS8zP8PzOJbV
4oIVf786eIw1pXhA7E1EHMVEUJPYKQNvVZPZ9nfBIZxa/02r9v+Xy2DurE4yGJh96nkNNtOCdkvN
h7rqJf+Igx6oBJ8Fb40pVS5TClsUZcNIF9xzzkBAi50QVxLogiG2nco/eob2RuC/CoABOxaoFiFr
3MT91IsjzZn2l0F8Bxx8dZq69Vy3k9vBmFlbo+fbexeHoofKrjwvydfhFkLiM3eJr/hs80ZbURCk
B2EuwAwupWkl7Xqo23DsZC6WCfMCq+0bredoCbItU4FpM02JyPgL3zxuamxOe1YY6KHLy9Qm3mD1
m3SkGkQDStpiAVRGRsXkUBXiFoaCobZc4jaibdKNxFuYXkh07e9XGx6b2MmhksZhdC4BmS0sCgmK
rzIuQaoCFrGo9SdlcPnH0dlNQekrn05KgkMW4ZdeTcWgg/bjUKDep49sVK73WPuuwStp+fBy04p0
pobV52boOvn7ETEm+OQRiLE8eZxiDkm/pnebA5RS278jhOTf9ZnROGaLN/lqHsJ1Us5bSj19PYyo
eJWYLhvEfGycxToucrq8uXon9SDVd1X6d40ep1gQG+s2RuFkMDyBLGK3pSm/sLsHug5SAMyz/nYD
evqMGZRPCMFKinwdr9pmJVU4yfT22jTaK39yOL8ljOeCHMZnFbKz7KFL9n4w2lUO6r3xt0cDq7/q
KRW7hCmlPK21OeNdzzVy6G0Pv+zPTVjXFANxscAx9rSKJ3wg3dMdfBOL97EhbNJhtm4pZ/HQS7By
jgMq1EwT+MmOTcdRlU4l6oRfjjdQtSBA2IPupcT05baPOjL7KrHyiiTuDYVhnV4ERE4pwyFdkjE3
i6qLvyWTKz/fZ9YQmUG7+ggVDVstHxTeT0WokZ62o2DDtzsMpCeRk79mNcT5vIvjO9PxhmB8mmMn
1X4OMdlZ/SnflWdrEpXbLXmt+PwP5FkEkZIs1b4bdD4/oNCxlJgabDt0zBqar9IS8K6cFhNVfYGD
vy8+lbQgrs+kgypd4KyGvDK6TLOiC5MN1TRZc7F1YVxYmbWW/8Bn82+ttruuVEQwWuFI/p8QKT0v
butPSP8ethDY93DrZEwhJRo4OGyrI5rZW0CzAwC2tbr1D/ae/ovHc82w/1MqDCxd4XalRSib+La5
6nZidhiZz0gQWO1Er3Uv4JHvphNh+PUxMUfwyLWnKMgaYVZTZJ5qoi1U6Q6OwcU6ha65tyNvLFaa
hC4KCVKZEGLiBAevvbUsLpcHzojE7/Zi3ZQyv8L17+DQo0K82pu7aIY87RTPpVmUN6eB4Vq2ZO3Z
9PMtgd02O8Rc5VbkM/gfXj6pWykWZe79osUppgli4aSiUKN36IGWgHbsvj1Vb2pLYrkslpefl3NG
9kAP7biUY8WiAAMJltpwbOOYoKva2+x6GaGwyeR0km9WQliGX34R5M44e73Pf1kzC1U/brPiXLOt
W22XFqnygQnrRLkT/U0yTx3Tidw/DW73Q7xfKanI11bqnIplxr+ZVJAMn+S4S4ZxFE3ibJjds3tI
m4kJ84iHdsSUgH4nSOavz7HqYrY69MXj/yaMXYzuVRyBGHpzZWSSJh23dcl0VyqvTCqTiZJDa4Fx
+Cqs73OPp+kzQ2eqWJSZqk2knG0jostS8ylQOVl25o/9MNDtSzh8RZDMP1DIzSji3IsQmrOiPQqJ
Vx7/Na9ViBzyLHB3r1BSydbXhvuR3cMEPfb/k1Kt5D5ci+0ysan7hnGR0bwX6XG8BBHsowaE/3p8
y+eWgPuFImikkHQ+Kmlsu2DyenJkWggdQo9RK4KvbAhBff8U8pYeuGm+XuEG1XWmbqdxxAvMlnSw
EM/j0+bCKa2k/jK7UGTXW5ngW0izj43IVcVQecPdrY/6u+AI+ZeiT0GNV9hI8DP0EGh7WzSLMv6Q
k+LnsEjj4SD6NSeFHOynACQPUpCTt6J12AlYAG4LZjQEkanNkEBvDG9wnR8zONOkD2NXZawvikk/
Q+80eIjmMNpSkdxZoAcQV6ZTT9D4mH1O6/ZFWEURokTwNJzzx5ZWaI0QdoOKtycL2wNG3zarX492
h+UbU7vhKSkLpVHZzwiSHgEcRfE+uoQmslAfpb0tyurK8B07swsbKsl74kWz6AETaK7Xpn50pOGv
Mv047anUGCLoidKBVHXvCnUNAjQq9N2Sz4HuhT9OwlOPboQXxb322SA4KpdIF4NMj0BqB6s3zmo3
Iq18PXra4NYSU+Xzft0CQ1yslsHfXNnGmNf7AB3HF1L3Bq3t1rXuYz8Lcrt/86/qn+O9SI7LScgC
Qj/rJRoj/CCjrU6fnf/pHgHHlPT/7YzM53tNPoD2trszzKaNoRf1rPYwbuhI5w+UmletJfO/klXq
pkJ1+zUsloJUa8tJ5j3SN33++UpEctYadYN92fpuuqrJv1S4cuM5nUohctkJVdfEbt8djyI5MidD
waZK8w9luPKS5qncFaOPQZOR3i9b1TqybRKrQ/xRzECwW67gMy3q6L+81VskGVpVULO7YTi+MUEJ
b8CIkmJAqL1ayiIf8WXJw87dFPP7eENS+cqjllNU3T4sHPTy1Uw8z/nldxazwC5HsJOVsgcmCp+K
27uH9DItDNlrlMFM027iSyOwf249RTf8sS91LIdgqBbPTqswajkQg4PSGs0VuMjkksEK/+/kj/gF
Kp/WoJEKqkIun4iRNwaNPrrEr48Y5mFEF6hz7/uSMaZ2atILPIM5eDLkxJOZxyd8k7xoVviZgsLE
jNis2jQo7XSGUr0L0U46WERoSJqEHoZPzT9a9cAOiTx6HZPaAAE6ey56sMVtcgiUx19h4TTTAzdu
/e6Ih6qlOok2BnMTh7dDZFzWUgltEYGa/5rha8YawXawbn3FoVbeBk8EFqjtEm+pd8z/vMTzDxLM
776s38bmpIwaXyYGbI37G+psdu39OHHm/miLo4z44odsz7iVj+6b4MrAuGe9LxapC8cRXnxJD51L
Fx5+Qp2UKo/Y7P5OYajUTkTzcIGoLumspVtwwkf72BFy7MozXD4N/mTTu8aif6c2Rv3BHrwOk7wg
yWr6nujD6Vsm/pLnmEJt2c8vO35XKLdrCsF2xcwWYqxjdnwFqTa5XzKBwBO9PHB9IJiFpz+LO1oC
LSmJgXTPbgsuHy/F5Ibk6uV4ziBzwIr+ilOqA9jMxLjiBIMgNZwlqPadfjzdduTZ1gX2z05sPvwA
dT/HBeU+vrrZeoTC6Zpiz36mgpTZjKl03xDdHaTGBiQhdeeP8UQ+8jP5yj9M4dckYd347eEd4y/h
jKTCYjB05dYUYfv98ZtaQC4gnuSnQ5vXCjMqMyH6EHnSKWQqkwzlSaErooLqV/aqUBfdzeR01cNy
jLi4u+Ok+c4Glq8kXIUpJ/rC/q7FHQT4Lo7eKb3+7JXrE8+Uy6/CXS4140OXgUtkGqhtiwqEKXFb
PLWXXWcUKYa+FnLMXBZTr/bbufGrRyi8stZNhwQBgMTHfNYyFVGAJIeT8cXntLakQL9TEK7lYTp/
8MMhkpKbTDA05SZZW/Z3Fc6mt6GxkUGn/AHRAALiEjyqSBqrokeUs1hGep48NWCjcYnJ0dUqLqZd
2wAk5HTcrJoHr5lTX9r2XTEtywFLw8uR6axObU1k4GjzTmfSYEllBw9MhhurJ6PK34ph5sOPX98B
CzMKLf8axjFeizmgJn6IojDBSEPwBBMgZkGsH8Ep4oXxXJkFAawvCoJpwAkIO/UzjJQ2DA3sZ+w7
kFh5dcKBBTZhpPz1DjvnWQHvWx32UX2cknB6eh6jxg1JiEUFLgT0U20xDZF/lt+KrocYG9I2cBQO
hPKxoglWFAySGYCLf5PRHxE/I1el1IisozSkrr9Ow3nVrNWM4mLDCbodbBisy9MJGI62mVNI3XsY
WDQrnk+HJZ25ZupKmkc1YiAHZllOtl+d/0mtrp4i0xtUo4fi3cbKtQk/AuBRY6jcePhXQDl5NAfZ
4zTXnxZY09MiriMH7RN5UqTG5BESom8UbLDTvVrl+vM/tTbGc9zm89gcrr5DVtg2GQ/J16p4OUI3
ZlMlThGwqrtZah9Rygf7imtLxQDGRkofGCEGqoNb1qIJTWSnc/6jzT59L5C3txiPTNSR2Ws8TwbR
SSUyjNoHQ2unHT92SSZe4OapSuCwba++mOt7uiZmEiiqdv21wUt5a3RItA0B7TO6Mm4Hp5d4Kgm9
ELMSuLT4Ebydsuyv8YA2roqwyFQ73XM6mtAbzJohUiTgXlEzRikFX1i5T4hnfDVZ0YfA6f1UVGjB
/ZtFe3KibUIyfZXGTH3Oqzf+2sXINrlnsQgkNNpvUcZrdXyx1Zc4dkUmroefucvN1IoEiAP5NO/W
3rNkmnpA3FKvXkJgIqauD6RSgrtMuq/7zyxwySXYP9SaqwdhlLQLckFHFiLxHs8NifpzEHFkYF/j
xkbWI7pksjz8Ga9xL8B/P7a3AAcZeSyehoNuPNe9iqhzqZcgvj8w/D9zs/3Us0UBJszhiV4ITx/P
9kZTZpuX9QgGEOwL1+qhg23V9qcu8z8nOhknUrDc+bJy4wftPjQE/lxrIWaV9DoDHvgEsycA2uG6
QVDF1QHHCLfunDmxp1vNaKxD7NXKyl35jedWqN098/BCckmKzDWigr/rRnrHTkbY3JpQvQcEr8Ik
7B06JmZXIEquNnOnlBmgpmswn0BKIqpXDW1TFrn+FKUprRZATqvdvDb5gAGo+7yyjrgTnfYx1oyR
wopazo8JVReGK/s+54MHhn3MvTuL28A4iwkFngIp3tRhog9c/jYQYglFPT0mJxhklUFekKjOmK3m
8hn0kSl5dhgLOKNMsA5KHq88NI/m0OTArE3Smvr7Ht3Wninx08qdpOqssMqrRRSm41URoqSciwRC
ENKbeaacjoP9kb7MV0lBe9ggWVJmLYJyN7tsWjNm5b0RKnyvIhfiJWL3GFVJYQ/a8Ai6lLZ54AVR
MO6yDPhIT2cByO/iY+Z4rjP5wIYUTwbcXXbgEkq3zaupmLAP32NpqwLevcN9heVjmOAygR2B5X4M
+DEtwb3rTJIAgNv7NGj8Jfcbj7TgBmfI0orkZEySjrsTOSlObjNuXyLA7s+T1WqbbBGyjdxWWjsC
HHd41f3KkJjd9X5wCSuiVEuudKI4/BFGsGO4ZG5VfG7GaG1j7rVf9eOOevq0JUjAUrkgqBB/fWbY
eKQlhibruzowqOE/7gVxMa3lnLXQQI8tSzdsQhKJJ10DTwdbDmz6ibP7F3YHFJ0Mq079uHQZ9iWb
NRRgtyG+VtmYC4cBdXq+VGL1Lq7ihLeEf8sNgZMMBZWQk6EyQzGZXGbp+UFXwVF3uyh8Sf7bZOiR
4iEmDQU8yfV0WNYg6Iojh2XXSCp+SSyzurZwXJzijUGU8XYEKu/y6f76KO1GWi1hdhxgzJvR4sl/
6Q8zaBJvow1rdT4cdN9uqfFzrfSnSAEaf5UAePtaii6xQyDsgZMiDmlXHqBzaTjcNbuWxv7OBHim
FpEzoUoWIbXO6xLPZaLv2g9wKcVXU3a/k9KRkvUrqFo9Mxa2S7xtIcNVYNnWm9X/icWliNna0203
R+9Z9saaesNyvVACYOdg/mSLTJKSeVyDGbywT+VT2IPBxOuZUkmj3mDd9doa/UblFqET1GzV+VRp
M19ln3kef1IOsDTMRpwxMHttUhQq12Jhs9Ta4ysukKMK7w0Kf2DzbQF3R7fql7xInhmJZVRn80z+
saRAKcn2EnYhTOqFAJAnvR3VE2wtSxA22cj/ZT7JscIi5ibH+/2Fnt7RZINAJCR9FxAsQaYDIe+6
BeriHq6JfjNRm9pbq5VhNndWpxODoBb+bToUcs7KtRAT/o98xjkvXGAE5f5rf4ak+aWYDyt0YDa0
g7jR6ZMCIsYMfP9zDBzlz48KePKWxwvuH5bmVVauv3VbfbUOdcrbuE86L2oD5RIbDrbskGXmIEvx
xHFDLBxNoGiYMO8ajnqqacV/sXKoepdkfbniXel+YjVVDbyYq+zLPgzA1thQPYd8VlvMDpP6wTso
WQSC7bMBf7VMPliVkWKx4iFU9sbksIIXk8OhSBruME2Vj8urjEVXA/2T0R06E9HTZR2PYYnccoEv
d6d+el2jBZZHOe8R8xbb6z1wQyMon555zEUpKGHsNGhY1PQ0UxClHHNWlxuXpUTDdKj/K+jcFHBf
bb7PNomXGC+qY17eE4xsItGzOXYQdHLyd8MF8TIpzoUdzhwLjIR8OnFedGLcSlK3tU5+5OgAcX7S
l1Wq6sRScIM8PqnBu4CjABKxd7oLwraHvSn+xnsRlPUn3GOQFWfqYmTsUam8Z73V5kJq9cgPAhkF
8xM8lDg30DZ9CyKZ0AIYKMxct7fl2/YqiLjm51eShsdEAFQIgAd/CQ3R2M4xXGjxeZ/QioD1tLm9
VaO6LpiM9Mq/ezWt/INw88UVsMOoMnYimp08tXhrmTFqLYxZO+b72en+bNYSo9jgngzAo9lEyKBF
8fSfmRB8jlcjzDsKe/mL9ZPcH55ebhCxF9q1z8FebHbeiupmvAn1rnVhiFJlp5oCkwiZzUBTYQ5+
+mCwnnh80EIpVVP/+YCMkYvCZ4wddUHwB6hFswK2HhWwu+wf1AXA1c3Ln6uMVoJXnSPm45DFc46R
B8unzi+dJC33bWv+a9Gbf43V/binf7bdDMRTGoh65EsSA1YTRi6sQ7UFufsTa5ec+/HSjCCJw1NC
BOo+yMdGXveqlJfwIsnt5aVkmeae9qjh+wUpBJZMoWG72ODZPfNNgIc8o54rYqX/6SyJi4EyuO6c
R5gNuHsb7oVunz4KqLU6ycZHBJU807DrdHY6U5pN42Y5gZjXcQDVa0nHh+XmSy0QWQOYcgIQwWu6
8JObsdym1hajCih5wRDV2aFJuggFfDQqSoxuOVT8c2Bcv9cRVDnpEq0rwGKedoriWHIZbaYFV06d
fUEbsB4dsrVKLj1ZDusNWHN80ttYnPTD0FhFab4kdFPc+8RjZGD//O0M1IPrBG0fzai/CPBC8iIF
J55TTU67+JpXQiNvhsawIjadBAPysOUyktwDICggRaw0s2EIzEdUBqWATgru0UTXzbyWaqXzg1iu
4I+SFkyNLoeLXkQ4XMC32t/5vTVXNM9NRfaN1SVxjF4n7Kxij7zWdAPDyM9MahhneYHCJ+wlOqxW
G6o6By9oEHP5z8wfKHegWoevSytQkcuD1E5jVFGkeXWDzRQqpXHpqC9zthz08OviLJXdO+3eBYPI
ltPC27n9BdYVuktVcb812SQawjEe8HlBdapRCRRIMu1n82kAVyuSBNdr16V2vx7xoajbiXPjfq0g
VTSmaeuJOKAkriNpK3Sdw85c+O3LoFwmq4m27mO0d7tYg6qvgN2sIX2O6CvpaH9zFSSLGaAtebMd
m1rcA4dBIP3TZFbLbomJwByVU0mqXVdIgiMb3A4x/mhtbZ/Frqs1V4Or0xuUrh6DFs3XHm8Xa6QL
8a1sLbo6C84KmkiLlRol3ILPARPnUVIyDpBPQB7JMB1M77fDVuHow7tj0e2sXMDXlbqYc1MZ9pu5
OaPQRw2/Fu7BqMDbmK1vBxqcwU5LX4Yp2cg4vnhr9YXJUqJLAdrMKHcZi3fQfnIW++aD7I6zCC/9
kBugmrWF71KMdiI01XhI9egZBTgR3oHT1CqFZ1pPXGfgfaKlKO0bLd0/7BVeDslzVxAV6wpdd964
8775nwefFkQA6hdWmhQT4E0DTwPgg95irQCYFlJppfCHk5heAOby9arILRMlTCx3769i2KalglIe
3haF/tumXfdL6Du9ZGIxM5clctmdXZwhwWzcPm7kDCDkHWugy7I4jhR3VAZME1vbMxo3xC76YKFu
9sOox6LbL9DlZSvi2BuWD9v+cl/9pEQLN8lfF0y3rFG8qmvhANInPH3+urZfv1AMwbGt0cdn4tUJ
fveRqb8MR63ENuaUrqEPxctQaqSfib56fXDrzTkBZComKrVSz+deITJriE146nFwRmfdeksO8K4g
SJW0Tvz91q+Awk8HF8BhiC7f1YAud7ZaQdzGdGDUQf6D6eI00uILxN8Af7e1qSpTT5TOX3jUSqHd
xoQvhrqCF2BhUh4u5/Xq9l8ax2aN195p8KF3O5PWrf3wm6pE4oN5JB3aRZ89g1BMshZTn9TSwZpo
TmWjK3nkms1SQgMbYQUBm7EvAIYbuqFlpFAsP9+X3iFeUIDCZbZgj6dKw9yZn1FU8NYxHNGvQoDc
3tmZ6NavYDhoJiEGbPwMq7FA1g1n+cIlLMl/uzL1oW5ky2C9fAUvEAOJ+I6VY9VBT7Q0+xSaalFC
hiNt6KztP6VDqcqbm+NBD/rGpo+fZR9c87ZQx2jLQsq/6P/rzRog6FQ8WqV6UlYwLF3jckFrinI3
9nb8ZUGfmB3zI0r5rQYAQVCBAIJfTL0tCRXSILMHRdv7gf81Mdge51wZnl92UgAsxEgq7XDKyHi6
Qbn14KekH1ozHR+b7JZ/4dCpULNDCrmUhHrm9EBeSAE4fA5gtUhMFrCGslzF88d7OKx8YLUb989v
ARGok8gk483o+XIaMSm4gt4M2vLDSkabhLY0nzBGQm7PcseYU0PsdqyoxfZkPzxL8GklkkbdRd7i
kkveXTMMWDVzmJCGgI0ImXWqtewj8sSwOudizbW5boJL8g5C/CONKQVXcoI92LVw6tmRiLQwcxf1
qv2UXRNJqeZ/pfbCRCnXj6m3KsGwxpg/Nqn5CnqqRC51wq6z6y2MxCzYuQtWiA769whB4PAEA3nR
4HtL+fPrg8B8z7/6y9CeDqfsunuX5no+nFTzmczKtuzERueU9KmBXsEF1beui5+ebvAaj5B9/ZwQ
G7tN7vMH3faFVng4p5jBvGPjQBUTXzJrDbRun8+G4/Fp0FMEyjB+LMYDXxkVNEC98w3hfNqImAzg
bWRrnadKMcYYrTd/hEcS7FfNsP/vCA5ZD/n3+sLv7K4bay6D96VnSW+AjHCMymWMCLoXPvYZDbvY
Umnr2wzROK839tZPHZfmfGfrUbnY65Aof9KzDK/eskdKc3/hr+84oDUkSZE2JDlGCeASDf2ZS8oE
SDqC+uLIkGSUuNWj3n2E8titjyRemrweDIbMAG+6E8H0HoBR6VjnDhMMPJ4nemHUcCosJ/3Igxvw
6v9nBY1/WOhPcB6ownSfxUY9CHTDwuJlUfvlrey+N97u3ltdEQ2cLvAnOMSIqpEC1h1BuiqMa3HA
JiO7NjFXuokl+ZhpWzh6Rr8KPAxyUIY2lObk1IAuX77Bv4y49a56BKZtKeqJeCQNebNSKo+yWj6g
t5C192s/RNaQiyF6TTUmDKspeJFA0Hpl3EinEqF6NaWW630G0jVaGZWNtJOQua8OGmScuSFnlIZT
XSnyPYliJTuPR3xgVJ4c/EInj/3QFc/QvQjKyIVj4c/ykbVO7DgUneaQqhJfwkIfNQZUSmrHbblT
0NDNPdfdJbVs9xzWMM5QGA6GiGs/NWCAv/p6IH5tNiUNozplAcLWemHo1wTnFjNy84Z3b+TXg3a9
ZjLYeDbtNF0OZdNt8K4YftDrAFvACRGJkjrzYfvD2PBRyHpSykF+rh6OW8qzrqzw/V6YP0caorzP
Td0QKcVuYpyEE6FyJvIQ2B/cg2KonoYHX95XGX1cw7MLiNnXqTiZg5li3lq8e67XP0q2i6aSj96C
UgeuuRK8/kf1Iaaz6BroTs8bCRcKjMtzaFzHmi0Y2Si3rLoQOt85hAUHdmx6/seXmEzCVY/2IM0P
QWgJip1ydom3dIs0umQRo/62p/AbdzGP3HJopDdIXTxDK1N0ripiNbLezWSELMUK/TYtGcLhCgnO
8nH5lACMqmFv+xIzc+mzHiFsdur8ScBKVGEnDLkJPN/9Dh2n5uLxc0ifYZBfkdyhdz6HkaezqWZx
nGZR2XSzw0GkspuGtXdjE0u7NMn3crr+PAiC+oNG50EW0tCF4tbuT86+dqathFQU2HTG+I+UAt5V
pxq9PBeUOz69JzAW3VoL5j8O0aAg0V+7HxW0XpC7zGIXSjNO73ajtIT5gc61ZUoXF5YewaXo7IRb
x14aSlZYQE40eWcNE33+MhrGhva6m13H6icRonRZijtDVTt5ERYX1YujU95LKE/vpfIVFE+n8GD4
IE/K/eVuSkYm57OckSkfMn8yvkp7LuADlx16BB1QsoJi1anMtcE7BVCFdFkEVera50SlzOIDv1S5
/07lKXxHzr0oCHIgH4ywEGKOr/USqxZp5unoBex+t5HqC5h7V51vUNCY/LNoaBCp8catriVi2+mK
C9R8zwhmnhWjsQKUD0TOE2EqzkjD/Opshdj7qZN2FIfpToOsnmx/6R6JhKayCQnbS1fhUcwyQKwP
Ywl8/kFuft+ZO3oVVgquMsmM8w5qkwAPd4SvW+F4lSCGzHpjDDLlQLvoci22sSmWaboLVnHv3SLb
c3JmpqJ2l6Iehz16RuLvUGWMXu2FgTsRhnt4ZngQruAX7EbFT18CyjRZhYDKvKeEo28bk8KPaz0x
gP77iemyUSCg8W/1BVlFpVsqu6akBT/uP/3TymktNrg+kxwUGiSanw7SSzg3cuRQwTDu6t1F5go7
ZsvCObsWTMPCRUXl/ADyf/+MOAmcE8zzJvpNvnqd7ITtvemEDmnyVbR5FOAKNR/j1YJ1JuqH9Lpw
Read7xP8Vh+A3DSwCB2iN99kcOBuiA+7dSlskqXY2NmrJyholR/Df9chi2yM0nYmisGEW1RK29by
+6oyi4sdh88l9zge37zJgiU73tSDR9u2b7Qp/qdEPdKMJXrD0YrazK9WnJU/lANoWdUtoVxIzGqH
6c2w1WmUZl1atQDfzPohGKaOTGR4sO9xu6vdh10TP9yS8XsX3OtbURm3Y78dpr0xksL/h2YA1rgN
PaL3CZ/AsXp2buKC6RJ1DyPlaTK3xw5IMiAKzCiQaG4LVX6UsGedBfYZc+nGrJCxZTqLDtz97VU/
kNvn8cKgusVmkxfjzwVPbcUdNNsuCJOFFx7SUKWP7jHOhUA5ceml5aZuOkPGsAdBQtosK1JsLsHf
d7fJpqEgZ0XJgq3cBic11FUYwctwa6lc+0a5MJWf+bi6cRDVR7JqaWaAOZS0xylL/gUkz/mBWFRi
uGspzgr0icVfM4nG9yZZ+Mxz6HOhivopZ8vYZfI5CaiEAs/IEoPBUpfrs52XhSJtpnIshO+yucnh
fuf20xTMP+nHaU5JxE6gtYk9UF3OYKrQoZYHnk0Nw4nowuudkR1FnxWqvl4hE9HiPtriG4dACaUN
rBUt61zrO4h8oPgSAUwocKctIcN1gK2ZxRxVMXYFpCDfaEVmvTHeiRcRWxFogZhQ4tmnd35nJbZY
GogYV4wpAJfZ7VrG84F/KoHgQ7eA+ONNHhkwAq7QRF5wwuuUw+WqABVwiFz0yzahhSiJuW5yRurN
b4iq2PZevb177RBAhz+YvKO2VBIYzenmIE12v4qsX2VTpHd6ilUN1ZgH7XDQKQOdg46UI2QyHoht
rxXj3Pj4ZLR4HaxOb80Btzeal4tPa0YTUzIKcSKsAvtLWP7n6rT6mg+67F0PCnrkN8Mz0CeI8Gw4
NWRwHYa061q7fVZfQh5s38sWGqRf3XLew1r0k1dMEbmGJEukpkPBZVNB5gOQRsEAiekH6j6lzp/0
hrZqJAaOHxL89+kGGn/IwQDiTT76z8XIVe4bpPJ6RFStOtI6berokt1ZlIKJoMujLF8dXbyjjTtx
xns1Zx8MQiB/fXJI2NHnLQ3BAMm+uuedB/tGYFPB7uYRmDJKDesHDWuS7MNjkGIKrdAvJ+sO3Wwf
GtyBvtd1pyMrUPQrnztm8hJBwB4X7fo1mRuvcaDQ9uTP7E6YAzMgrsdqAbvOkiBnv4OXjgFvtSs+
BWh11vampe3lJXrtd7lfkhZBNl9YidqVCUj7GnIGbYoy125A+3GWXTRr9KtNQsE71rLZVi5AKcxh
UGx9no1GqypgzWL1LOh0epqcXv/U0CD5CRRUSI+jMFSPLRacI4DzULCwWjcbmB+O2FwgGLDdSc6r
fF4oyS8BDOD3lb/fA06c4IbL8tyBSrxFmcofAOSZDo1rgjef2Li06oVAfLUSEpRg5GYBYa55wcas
TzKbCa71UFDa5dQ+BGPt50aVYwdVkfwD51nI7FnCQuTFWIMfOO7WwN54jMLj8T1xxkO2JFiX1jM0
JV6m8uT7T1ku3WlY2/j54q3lbdWmajkDSYVGM4VPA5KWk1ZS4ZlPmmTohnixqY9f709HCLh3w3rM
R5CsHDlxvUGRbatckuYABs0FsBpqHe0lLFGCzUySIdh7h9nstCRdmoSDQKG2mV0sFrLfPLBReTVD
G7PMwsK/b57M+Snh4AsxRKAZYI+QyN7Y7ur15GpQR3yyDuFp+nkmF3hIJ2Ugrb8ZYJx3sT/ogu0O
i7eqcpiZwxO/B+rUSSdgUXj55Qs3wPKlqJfE95t7qqYQcb2awaS3cP/IA7lTgf9eLb40JIJhcC9v
IpNAD4P4+Ht5pVj0hriLiMGpdVEToAiTDu0lJnpi0FoJIWgTK8KRClEOxLUdfMrbfImNQe+u6al9
pBh3jZA4H9r3O5lGEak8r+U3oi+KpFRZxyTi+SENPoGWnW2bZYU56rw6QJmZay+PIdfZXW+I2Qi5
H3Dt2HAHtj018Ozp/6GARRAGQtdBXXzYqp2m1FwoH49PK6LnRDwd+hYCI17OGiHPfrGv4VyLAigN
nDx3+sD60P9OQ5EUmcWhbKE6FdE6k7hZJD0oKJ7Z5TWscrUr4ISdQCJAVrWEnwS4Vih/xKEGPb9t
98mmAQZCHHsqG/0bIMIeEwiVraJsf7Nw8XeixZjvhk0GK2i4lbGVH1kp4iIoxi3ZfJIu34ZNhEO8
2tg2uXhOW+EPPRseRC3bAp9LkywXqVcbuu2KkTl5Y+epYec9L1Mx6SzUi0JYMtX1QRoSyRUdpVVR
t0HwGaXlVyu4bawCq/W0P1ayP30+n969+GtNIPCE/FZjeOGDX5N7ZPiElxP3wYY9RwU6TM4e7afz
c1lc/Pjw9tJXgVLNRD3BM9OZPaAbYQs3OK71bCRQEIAFQOEmiuNm7TUehfEiHpi1zfO295kCjau1
kNdqqfXcL16MM61/JMCY+5FsDQlexN4V95UBP++yK9QRGZ3BiJPjn0vHsxa97LNmSUxY6kixG81m
X2Kqyt23LDVaoDGlf3rHKqB3WWwA0oX6dVwEACTP+h0b37XDERgFkvKLLLaAUo6CWiaMuCMKIuqi
bS6n2/lVosmsBpd5EYGLBvRUTG48QqfBvQh4SpEDWrYl/JEZogniaiRxurKlZy6lGsIJxPBCwm1h
/Ucqp2iqnqNmGRJvb21H48yVfqOGoTwo4qjRMlznlx4RpxT8Kj/5+AhCd+nThARXKl6PwHbg3TOt
6GXnWS8TG3aa6A+KxGHmw2dtPuocHSw+nwV1wZ+29Cu2BKVhpeW3YXk0ktf8KxTTNQVQHpRScn0Q
xlYJEaNW+k0OsAn/mcoNpWuw4kphAk/0uSZc91rwYz0xekZX2aSBY/qYWk3G1BgMdb3eT9IsNUxS
ZmCp1RKT7mwHsT17Aa7QAYD27P8t+BxJFjuAyAYhdax/DcAruDv/mEMGyDU3tHWb5mMWcF8EO53v
llvvZNpMMzT0CxktrcVFVNCqhamOxS4/4uRfoRe/BZ3b09E6Gw/7IfO05XcenZHJ4txbbswZEcwh
i/y6tPejKkG45+WVvQ3UkEr61uEb36hkX+wEMwA8MuH9mZtdgVgS7CysqlLSRMipLUghCamlf3AZ
rcQU3JPO/HMC8wGla0tOvfAHwEmPKii5cMPfBpRmeqI1OLfiMmE3dCGjd7OIcgviCMzLwuJ54jo1
PUbUFg2sXCVzVkFUmuCgn5vE6rs/DCyJ34FjqbPhT7nxp8f3axATK5jgLey3gaXss3i8GvoC65tk
CgoIITcFgP1l4IV/+VSZggDyrEKFX/pkBCBs505eAKhzi6iojJOyMxURXDHgL6pZSKfMHKljoYi9
7wGL8zJvKkUPdrqdSOBFqzjRrFkIlNRTJAhfeoiBepHT9yYBVq59sXmPjjue+cUZ0gFItDC2AAQ+
KU+rJruCEpkWMDxJsc3cMQiIDTjWWUQXOMH03yw+0oaj4BAH4NeOFTI6j7PxnDucDj7mK1JIdX06
ZksikA+D+PhCPtIy0Pjdy0xrDidBl0P8UQ8QkFAzM29DsLMHmdz1XGKWGV9SzWE0gEJMIRF5U4Tm
To9kec+0E3bACDw/O68AW61IFUIDTHHnSoESChmutBMzSs6v/BFUkEElONST6BAkgS7/bEZ53wJt
gBmD0aomAotNQHtd3nT+rjCtrf819uf5sY+IVaxgUMwXG8L11UbAkr63wHuFoIfpJmnGMlncqSFz
r0z+jTiMz21q+9MvEFLe7kSHGF2BQ/M9nLQeiIPkGD7o4nTlCwn7WqQ4jcA/CvYfv/cBgiBdHHJu
mEsObB9lPDV/gJL1fpcZn6N/+A8/FxudiFetRRIXYd18zeiVQ3aHHGXD8rv5CTrjwKHlrTT2fH2O
ABCwXjafGLi79lKf+zR3qhBsFyZvofQMGJHMBZbA1+C2jTRj4VGapcloB5ed1qWNBMO6tJa8ncfh
X5A0U475M2Bq0/wmpgt5/jRo3o0nWCWJ0y0PmMhlkylZ7wl68Q52jJ6JNwSKDxUgNKH6tu0Qjp6D
+6YmsFJH4Qq8a8uGrktdfO0oyAf13v2hNoNnymGVoBkFbv/nGLv/QCZ3S+WvY0z3LhhPYt+KupRb
bf0b48LAmXKny3mGXwGGf6TdPYBoBLIg6mSETA67zXy+VLbKoi+ZUBonD9zFTKUMOebNoxUixZ67
Isicu0oGl1ZZktG37N45xHkiK9m6n89K0FpJUno2LdewjCeVAo6NF5ofsQsJ3exd6+QSAKjQhAw/
4IW4wOI2telx146yfdmaZ+mZ0/m9HHg31bgY6iKFwQB6CobHvz9Jn56/aOCZZi1VAct3EC2on1uq
+5sXSiAF2zCu9HzvGFMka11V4ubXcPG/tKUuG4kgF9C5yvBN3b3YeaXMwyA/hTjvx4ZSGY02VlPf
QAIta+E4MY6l+HWRwAsExkZdA57n1KK9MpV4YolZfTwUbvQdrUkQAwkYJLPr8AZSi5MDzPjFfZk2
nOVAI/1uiAK3V0yE3RcwZJlni0DtVaxd8AFkGHOwvlw54JTONlXnzqJb0zevlmcRrzfrGm1jHkNK
oqhr1VBhw/SPapO8jrklgqDgu7NMp7TjKOOMhP/deYqXO9FokMQsKUR+iPzR+vMAhBt4CW/G8A/+
4jlHu1PvZkoaqEbIpTUnB4U5Df8N6o5bHH0U9XqXdfazxxYJFck34SKVnOfiwpvlLnp6Nd5NZywW
FmLWcLxmufjMxkeTK4JGIcp8CYyFWGQ9zi293Nta+49ZvwmLywQiRmCgU6UQBaiu4iliflj7sCkW
c5tk26+o1+TBc2ozp+eVnR6E+PZRCsGHMGl97A/CzTvewTkjmBiVcfeOyC5G0Izph19eJQgJKYau
z88wmklgKVY8ruRbmb4aw8RPbkculYHhUpU9Ii9MBJLCZttnoX+6Rigb1AMaczh1KpdAHqXX/9xJ
nNZTVj0BN6EzU0pQXwYDC/NYcOustLbzxWZXavUApAGSaMPpEIGigg1YofN5uTiKrQslI885seCI
niVo25nlmFqbFNbylHKBs8BqqXaA8LcJ2s/UzfT1I2E4+IP/Y4PcVKyuYl2NXtiOWiL3jaq2Vwku
QgjSdelNA5cFNSTkkZWbhAZ+QqDwvbEEPXtvTLELJhbyD2fiV7WgxXGmY8Fq/mWjJVHX5hyc6jrP
US77YxfuoQ1XWSWYwycb9guKS8ZO6GLepSqtsiJXJUD818gcaEHSdaJHGY6xwSYs0ScQNez02dvi
P+91xvV9Mb1aE/+F4ousRdnL4Tt/r5FGCcHYk98Z4Jb/Ldzh3xVt2rh9s0hoPqytOa2DeNZJbMBh
DHWpEfoyT6ewhryJ7MUG9bZefMGDXep4wnzvVXZgeJBkVFYQ+T+vYXj+fD/nqP0dNuZh7OxIpRbT
CRiZ5Y7nW/8dk394/42TFJ+qNcSN8/ix0oEGl31TAIJR9j0sZ08EE08Dnj8NMwPERVQvW3ciBri1
sBnxLXUdQGUgDqzoF0fN5UMmTPlc8/CTN2rKhOErTBLEc6bc8bbU5hmnZ33s6JDQ55Fa0oJoiChy
jK8YXCq7zdVy1YCK9kM0kPmF3SYmmtLwEs2TCz2NENE6ErNK3k9P3cNOr9BjDPghwi0WqftfAzG8
1Ft7wu1vjSnAswtvf5f7IvDHFR8Vm75SJQq/SUslClPz3fqqM7rI6mXpDsUW3pVKh0FIZDvNxmUd
T5GaevWoMRu69b2I6CCHEtsEEpY9wmTWQ26t9XjL5en5r03O2e/jNTz4guUXHeQ5HdaLz6aUwQN0
JsoWcdzAJ28HUuuX8bajXNq4xBvG51dR6a7V8yo94Cjd8+HqgwqnRkLDR6RovXRpHRQIjbp0sTFL
SX7VATDTX/v/wwtioSAtLdDRSJXKlt7VWTNEiShSP8AOdS0Hl1K2TbIso/lwxoUKehCi67ZZ3rsE
h09vKmfaj2jiRD/pez9GP04EF0vD4lyaqrjtfivx7G/Y9HmmEH3YS2WfxYIB2RXEHPullE4KPSVB
BJ9u8ZYv72/f9wP7BIE3BZDB1O+avjSvKFkbw43FByNFjuC5SNpTVZhu8dYVkclk9R71ea2hutjQ
ZS6H69d2gyFlnfM2qwXNuNkE9ACBlulIo3IOs3p2hlBR3VqFNwGZgHs4lgrC941lUjmv7vrptHRL
cX7abVGNsXNRXaLTraf/RE3UUst5+4mn1MNKTI7/WQP/fO11U5NAXazkhbf2CdsbJhHz2wEbvsLy
TJxFbiky5gmM/NR7UWPl1U+711q7MGThng0oxTxTC0rKNBLzS3FDza3LXNlI3+UVTs4TnvhpkvQq
L/A9ZkwGZe+HDWWQdY5echJmBn/v2NkvYgxvJQZnOeApha+M34de+qZcdZOVG9smaRKP+v/Durpu
5QcrS/P87SelDh4NOfSFuzXPisH4sY9URukZddqWHtMEQKuqqtSzWa2uYOYCl3MQ/Gvrlla1jwA5
Za5o/lQtoDdeio8/1eqEiFTVSXIfwQHs5nQrSbU6gtUAf49ynGgiXnC1WJr8xRF+Mx2/H20HJxRv
b2nDk6Tl4NAAbtpoOmBnUD3BcirJ/XLaBPas6GJAxytzjpZpA8BRxssR8AegdHs1Kp4bndjBFCon
80Pq95uMfdNSDK+9thuEqVVIJvieLflBi3W+DEViToOgObzjAPtvwDUCcYS8b7h+p/WnxoROq2zE
oEIecAXV0jkFsjmnSqUKNaI+/TuLNYs9eRN/4iiAIrgJO18Z2fHQW25Q1Q3VIc9G7E9YaPqmJl6P
Xs46U93lAjICeyLl32RtMPSWcvq3YvvF3D+ZVsG3F7G1OVhVNBDdYQiKFZTZ2rE7StS4ufj5yyBW
la2KyIIJmZllgVrtZPQDsYJ5rZFaimc5qs3wjJRxrhvzCfkst6fwY5fM7wNMEyI/UW3cfSEcsns8
SWg7pXAoXze20mBPPpGHM/o+KvQld7LTvlQ8DFS9Y4oqqGlk48jhvSYW8AEfRk0b+FpB7giR+RPd
YlN2C5lBzzTtjYOdxG88Ia540jbSuUkNv9y83GKhFe1zfL/eqMGpLDrahn56HudRSecqLsZJEy0C
OhNCvMJJBy35BJsjcdi11TkZ4XiQPW9P1j23806L4N7wOE4U26hg0c8EFeILshCxemWEVN9e/QO5
zlctBVRLxTaUhe0TvKGqcHyULTmRIldu2WyWh+swb3qiy9OcA9EIF3a0VJt7Qan/31pJNRhIO8QC
B4wUZLqzuqsJ/wuwAiTqipaZB7hjLE/ZBNQZlPIXId0uIYFOFJEDVOLOPpCHks0Lc+wCaNlU4ytn
8qkRCVYTbBTex6PwGyIX6b5jCkac3fbK+9dx+QmkcJdIJOsZ1irnjh1b/iikgOyPNsYLkid23BPu
Fb6lbjum+ZUhDMtIp2u5mMKoyZQPTZcrvr3L77yl0WxNsp2Hhl5WVfgSHI/afhkTWSioqZtevop8
oN06psJkVV+oBLExLTD+XSXWL6kJFuKYmeqC3eXhuqIzzQTA5B5CX2di6hX9qExcjP9mnKoj73SY
MaChDeipeDvMx8XTB7XJoOe/q7WSXps0zsXU22aeEn32yr5bR5FN5s8W44v35mQf+6QQtwgsaQB7
pBni5X1mk05WUEJuIIHqBoyXeM+gk4KKwiuLxEGrXakXvDnE3YMcpoYJuhJ3C7M1HG3mtzXl2I5R
L65L5okNuYnZ8qrNfiyqaqvwje8TYSZa/EZRZi5XakbXdNIRiVvyb8X93IeM2L2Sd3Y2F+WoeUNY
7aaUJnlmbTs9TGYzzkmyjCP/LMRGFOW7p6VdKskzeB3kp6KNcXmwc4vCsFeFAIEMIrxREgFfbZjS
/kRdqXFCYnNlK6cZadxor0LIMTL8u4w8I6ToC8znH4HksFdNOrAwoGpHx4wfLTM83P1BNndwqpAQ
zeXDJTl9edCAzw3SiaGpalOwxuoNBfE8vQ6rrD9vogsRVDayKQLPELZh9ekrvs2J882vqLY+ZNix
qvWlcxFKtHSO92qZqovTEW1z9Evh0j78lgNiR5UTmrcWZqEhlQ7JMtYnVjfUXvNOn6rMFPqfviIb
QYjzGdrkcCjQoQuLdR/j4GaOdxvExN0dnfK4ZykukyAXry8Nv/A6xodCEJx9HzkuvMtVc4BCAg1c
OMKPGSHnTGuF7rlBvvUW+v+arhTme8SlzjA7kW3QBekVl/Gag1qmn96dNtxQ49ebPszt5DLsx6v9
Dp3hQO38yFfOzMRrrSzAjGsObHKiCA4dahAryNCGRxlMcjMGO9/NlM0+H9XNuZjylLZCz7KexW9a
7buybghH7bsBx6wWgv10/uI3DW6wEfKzXGRhqUgC1DX7NusOtSQt9w7wtreaLFhp50rmWnRLgFEX
1XGHi2lbghSy6zgBK9RYzxWKCvAA6cX5jjwtbFtOuKL9xGL1bGeg15o2pMVRfGxGR2EnXLun4qaK
uWgYaTybfr1ttSIVink/AFc4r7sVX1NzdS7fFGiQ/ptjIkZ0pxwPlS12d6JFtafLvXfhb1oM2hfB
IUpD9UNh9JH3YOfJyZ9gzAW+OmUh3bhq54Tq9ISo9RHASb23+I1YMhZ1ueJWJpQ2ISIUs1FTCgpg
Qzsr2BUZiwgpiWcbC1xah4Co0GED/O0sBpzUpSDJpiN9bzDDB0QhMyPi2iuRbTrn0ZX42dC0vqRM
Cwsn4zEMn+vNE4aXvZWoZ6Hm2I/cOjBt2iM9IIFYa4puclNpBsBAIReL2OhnzsET0D9Kwn9Oq+A+
j6hvEmPazakdY5pgTniHkdeMORjDUWxvHWeR7+cxeo6gnE5vsbZxoqTr5Ycs5W7H7UbdyGHiqxt3
zdDx23F3NnQ5lhxVLMwveFTjgUM5xB8dZYfQRU8pYOXJfyrWAjvbq5oaj7XfX8iYvC1qm254NGtl
SCVlrcLFfMC6fB14cHCUO9lt7qK2gis8P91G2/07lyNIEnvWQC8E9luqCJOf/BGCwGGfjQHsHK25
OI7I40tFpBLLnE8AqpTa+VZYV9kzx9kW8L4uFFZK7bjioNiKrw38sg9v73+tcRmRGPfmZxLSPm/V
abqDAijVDWZqBkNmpoCguecshjcRO7/4+fRKzr0e/y1NJfkxNcxTfOE5Li8+JsQsPIi4BEXEHxBd
Sx6Wu1go/8ExEa3AnKfFtT4aQxrUpqwSBrQGPGy2N5W4pOfXX5AHolFKib79iaIwUjjISwosWVVU
19qYi6dNB/Z6HLlQDlT/97b+svdtmA3rMAbFh6dmTZP+xj8LpB/d45QgDntOQgvqK05LD7CMwJhG
K1VgWUZ6eD+HMLeOsqgSW5FR2DFcjcKRy5cdUKrvj60/z/PLPr6Wkt0UmvBXzV1U+luJBMZ2gB55
9RgC5kJP+Ns906Tk3ymaocQ0vGsmCyQA+GhRNCP0oAM/CQ1PgZw31oBiMyPrx6fIKHWHGZOCHf7F
1OkTEA7I9V9btWGggw98SMpUg0j4hERiy3j9Xe9ESNRXaildvmLmWW/1BXth2eJ/kBre1PVr+QSv
iJhC5vk5OP9XUNe9cpBFVl7lMwQY8Q5YA6dE7ppTonmSs11fw1SCR8u9YA93ZLIBsz2PKPbbQkD7
gzyt6IaUyvS9QoSGLcK+4DQ5aJIfzkoYZ77yh0MnCUzJsomHxUpdtMmt/5qNmteqJgkVu3ZvxtaQ
qjquQVJePttCBRR86Q0cTaXHA1E4s8EGXm45IkpNg6bsENAjBv4JTvIYUlVGsxWLJQGkZK8MSx+D
6D39kX6O50U5Nkjw2MteaRd1SDo6imIu5H46yeJC+CFugJ9I86Q0tJPkMa6ZFyxI07DIDOKSQtM2
6onOflo6q1EZ8B6EIDgqG78hrYLzDkSgmFNUQvqXeYaORUrPvrY7ffix+7GQmmCgy0Y194wv/DTV
lUKTysR4rrpQK4pMGeiPO//NsCouYE66iYiI4UpGQbmeuoo54KocJDiCG2j3kIqlRurq1x5uIZxb
0y/n1EdTUuOnMwJf09nAWT0qUdUoa14R+khzhB0R5MOXVZl3S9LoYvPpRDymhVTfNX3/iCPPC/ch
PXlG92GfS9Gi/rNo//ssibpntOtksoiBFxHmTtYM+gGknwnozoBt86kDcnnNoBWjOtmM8gf/vAQA
Xw7YisxbViKnyB+Sdncot4vbeGp2c4mMn2QLS+mSmDww64Wqk/uJ72SqwOPK8yvCoYdXMyKFvX0a
u0YZgrVPQDGU+aX8yqm7nNVvO+ZrJ/uiwvycxT0AQMaKUOHuCk6hP6Fc2rcgPmVlnsGVgQocQxTc
ctK1+hzbHNtuhtiE4QVS4Vkv8AqPSn5IVQfiQOPUokY0/f/MJivKCKAFuKS6++HR0bFvQ8C+bzIM
xqYqrYfPPeMvtDBDS//f95DS3Umb4tVuFfKT/hC2j7+Ckmj14RLB5oZ3YBx8KV3OKEIw8MmFd1S0
WKA18lg0+Mh8yaWTSuI20Ix9Mq7y65u2G5Lp05oH8lknxroVT8fGse9haQ3kyH8D5KRX27w0rggr
JLilJL1vzsaGcYK311VOXkk/9r7YpZDA9UIzoZffmBjUs3UPWSTJX3wtufyg5FfCmqZ+gNr9GRgp
ZV1RFrwh4lpF/vL01HD+moMbURIOHFwJPEstpeU9x3PT0uDUwTxLJ6+YnR8OMlyD5+RYW8wK/Hk/
DHLyKJIMJHBqoUyIyRBnt+cO+nch8rcpiOGVHMBzDSjfI+S35TS2Wt5YXkJJlen4O41EV6IAHVkU
XVmxZCgwsFQn3v0JYkvsNoTkVuT07XYdbGVAKoaWbcFLcTnRs4xGaqEGAMLS+B+18+fBIe2+gUzv
m5/EO5BTeF/RK0tQgwtWZh8mNhFhjigNOa2KUgnarQdqfEyxQC6hBN/R8eC326DGCNwzIfXXmVlf
R8FuJ80H9+KrZHpLU7WZmAXn2HBznWROsxQ7hpXWBEqfi8G1imj/JGS5Yt5y3HOeVt3LSaNIAbnz
qmV1GRqqRo6MG+mW5tmHrKCyb88XOvcxx9HgWN5Fos93u7zDF/eAhL4lhGM25qujFUWS5mpw7rxc
FOpbMfLKeTneB0Dp9IehyVN5kuIab5IUc1oaMsy6dYfaths7d8ZtWXwFyUm7HlTYKq861q7AaOIn
vtwwqQ/y+3iQN7fcXvYCRohOEJQusMioNN8LbypdxR5fSxM6RTcMhYDS01BaixGPTWNNrsxb+aLO
wRmrj9pgwu4FtkslnsHp7Al0SiSJc/bE0Ja3p+YLxf9wm74MUtUnNwsWCzIHZguOlKvtcgFwGf2v
/DPEssCARb8ggFi54fL1E0XJE6zWpZufBb7pOLLkf+xisvndzI6bwb09Uynu5m/PCCikCFr6HHZX
8DoYCSbyWAaAAde1lE5WfvYdQVg5owN4ycKqLLq9NUlGVSErGVZBwh+TJOje2vaW4wx56S8T9dr2
qW0LUR82UeYm7P4kppGzGeJp+29OT1JDTBpfDaaWPSsRnBG3asSbCgbnEQg2rskf/Af5UtsrWJ/A
OBz7EfgoslBBwg90lTie1HzROsh9udjDqjCSavpzpk9SzVErTHE+YF7Tt9C4sbYb3tCTlr+4EEEE
QhllB3yqJ4ZhWcAZWFkK720U1ojQz7o2mW2wHRgHzPJ/RMPlOqIjI5JKI8+o9XMtqLtXfED6+REQ
zcGpYhX1QYRkMPr76os8WOMEcEGlgvlaToC1iXLNNo30nemy2VMuwlklBHWLmxh9WulzADBOTQzQ
zZ9GWyOvVNaEZf3xY8cSjfJdoneoj0AYA0EWeCknoMbpzk9sYF4UhhdvdKx5l8ToznhR/BTdwhnU
8A/QLOcMhAqwlUcA7any5Nz9kV+jRk0H6Ude16Ki507lE9YD049lnfXlwiuVFQa+fLUTgPoG8yyM
OHkJ8b4VF7z8iQGoiOKncHiQaHBbvnJ+xbu52sonwJkcO8SomTUgQph2DZtJAbXuObG+ZBLCY5HC
k0n8kBMDVSNR3bzBL77ctA6Vdf48xOvTXuOWzlvuR9HATHb0X5WmxdKEt9Fx+V95oElF2jjq5XJC
ykZ38mxD93tS83mXk/dXp3dAvRGNea4v2EpV1l4iHAQGuXh0u4gt8GdI+fxnp7qSokoncYe5NYMq
6Vf7l/FyINaF3A23BxbfiowHLOzgdgilILI7UoTyDJxtsgkH2wo8y5tjp6n6qyrXAkmVdOAbWWv/
mj87B+A/c6gw5fBByNhVw4uc0qdoAuQnIzpENyWSObByAeg2NWEJDmz2APzFqnWYppFB0sYz2pUK
LduZbFvVVC0cS8bp0cCAwnynlHegCYz163QMpSWEB8SyH0mHae+o3ehj9Fu243Rx8DFPuuJsLeMY
2NWEtreYAkETZpOVec7VJ4NOucVpFDeqwvqUC8dJ1qCiUom4A7z94UKai9nq5H+hleYOimxF1jl+
b56HzeTgM12yDzheoriN+RQ9DIQORcofbaGDS6U8wjHd4Qb5sWk6xCAUnkD49qSFHJgVyVRfp/q2
sOAztcG/CQyXATRV/xGgcTW7OkrVkYSUCvvuRQ6tZ2ctj+QBcL0OGhLyOwgh2r/2tYewtoP2/val
MIEa6ostFiPutPPlIOr1IevQ78eg1MRiGwrwVrXhZLviwnVPkR6BipPs+dxMkMr1k32Qbk4R0ded
UNJc6Icq9Xn2o69pMoCz5COuevlxl6T2Opk6L1BAowu0paPoGlj+ZJ4uDQP4nfVLMh4kBpygSuCV
XEEQKqaes0DSdx1jfkYCf5js8LeHWlqM+g18FgskIvpljuYFp+u1GLiv9wGLrxU60bzh/A3k9V5B
KXFCq20KN2R9ghAYI+GcYuqU33pK4a8Y439EwzRiJryytb2lyDY1AnECTBqFlzUkSxYB2T91jn/8
M2ABXqfZo9vDBSfDHBXJOIlJLxkg7SEpZ2jb+LO8SPUbAZTjmGxwGa/nRwDwuDjOf4ol5rEOlcpk
cXXFwR6lBccstzpwV6wDk9zOtyMoc7HN5SB3Y1uUsNa/lJn+ruwPLPglDs3+Oaz0SuLe8yOgreho
3LDwxRNemxwX6rzGiHrhnEqsUW/EWd61C7Y99bWLiZCYnF1+vyzYu2FyXrJG1oCtt/rqOxNNmYcG
zvprECKfJdcP4Dch1hO7Vr2yMdD9bFEBy60gLasKtD3Ta0y0hBy6gCu50B9UnCaxM4VuWB8Iqvxe
FABXhMPEOYhzRRWdjRjH127KZGzdFJM+sU/pm2Tp27Etx20MP50jFNVp7AK6CDTSvMxsk3+2TCCp
PfjI6zR5Eghgdf+UH1HCpD7qOS28txvTp/hot9cackLQVaX2YeunJRvUZvT3H7TajMrqnW4vg1Tw
dpQAkMcE6NaVcY41DBd30aY6OXuGGeFk+SjfJRTkpsqvy3SX4VksRPwZuiV3HrdozJP/HDUFd053
wgu+Gw8BCzgNjyESk6wbya3pFbYzJbIqB7EUtoRLW3euZdJ3/Rhxtjypzf8uTppc+cdXQYI1sCTs
6QoSXpUFhjLufujPxZQp6ApynSiRWxsvdV8tfv1l7KqZVmj4/JgILH3f7sFPk+aE7UB/pmKbDSel
46rn+r/Nea8UzgEyTyA021b5rQXtmtc9esm3x2uWWhnzlK7GhJa5PRmhyc60u76J2gNs+lWnN7Sm
BRuzv/TtAv0NHjIwoXpM77FDfpakKZC5ffFGUZuWQK3z3TBMdacrFbxdgZSjFHqLkiRPJ59l6XcZ
UGEabhvh0IDfuZDvt64oUl2ca8mkpJ1YP9mlmipQYc2qa7Q4FiD4i1K8rFbUba9XRV8R3N54M/i5
ZICOyuHt6ciR8kieKGjz7DbFP5R+P9hly8GyxkuAIxXFKeUFoPe0SOq9AUtNr28eFltAko9UQUWQ
/Fbi8Hu/p3TneAXDlrTW+SnrTYPmKMz/qPadCbJLYRZtSjrQpvFRbQwmXB8D1rpL+zqTYlCYVz2/
7zrmejRgExSOkq8M6iRfxSKyghps9HNbjIzWGRHvHGhtUaICNc+qlOuZzyZoOqwe73b0mrc6TPa/
57wpXxo8yBTNOKBGkuMsdIKPRvQu2d67imHQt7XDNQB2kkpGBasMaJe9nQr0WFA+bIG17tA1AEv0
udlhkxIybaaCqcOawMV4AH9WB7A/rxTwQsxDK6flLnerOX5QCu766IWu91ceXYRtaT1eYjMLrVKl
hYYXP4t6AzpxOfExbiBrkW2jO5GUSMUsP5X/AqtDqv4U3SHWgx4xrSyXByxJdlm98xHp4Fsp02nw
hFdxGbIzjKsYzPgBi738QOp4AuJreet2FQG0n/ipdsK7y0zcHeh5BylZ6uTvnzJZt2GiRZSxfvQn
QOGnT9rngBT+l98XDSTKe7wqR/9RRBpg4Q/YVL10fUvJ4k+7CzU9ZWw2XCZmS4OT/xbIULM9bddY
ZoLxIcWeXYoc3FstAI0rQ4W3aBt/KfNK20IjwvZNPUGX5zhlXuNI2EM8mxDk0mM51XH3g/+ROQLo
M3RwrPQYH0cudWZ0UPGD/ZDysdEov7Q7eiSocOoXfxKv7TrYQCGANpZMxAb6Fji4zV5e32utqTaH
W0j4zXlM23hJBeN+x3Nbaw8Q1KyMyKn0Nl1/B8/x4ynUXg3zsjkEK/IcGAPIL2ygelNKCPsgkECn
uf4Yruye842rwNm4caQfxVKUxI38ABSPry7b3raCARsDNPkycIpFH4w3eV9tiYKfDVyii1DjZ04r
h/mhz/RJGOCAOT2H5OghuX0bFdQwpnXFOI2v6maXVPLgeK8uZKi8PKEVPrRl4PNAMBAK2R1qXg9A
C+YFcFFI0VHHNIFDXYYkER7jOAHuf3b5A7UToJ1CoOfLpNaoZreVN++AgUMZOw8Yimlqf7o5pcXN
utj8X5iSrjB2CD5SLOJofiuUM5irQ26acjzL2HlsV+3U9hv1YVJ2zogVfOChR/YApCCv7NKTrZcE
b3hGeIHNTqBd4rG9mVXgFRul2Cca8aqfIBRtNNI7S8rLPK1xa6mhNRSO9ubXdefuHOwpT+S9tOJX
rNn1DtNO73gK3MFw82Yq0HuOqV4dMpcdcXDlTrLEDG/y3ftuFO8thO/ikgEtw5HuYUeGvWEGTf5n
FppAESYprIc58FgDL61Z/QrvzgPuKYeri2invOStytHrROK7SUh0bfZHAK+064anOsTZE+TDSw4e
k2LYIV/rZz9gVdWSmfYSIxNFM58ZukYjq0OL0BAqrhoYoA4atp8AcG5S8RNL3X9+okdStnFHpzty
6aS46CSQEFQJcx2JH/pGqVBv6VMQsZr6ccEI7WOHYqY+1p982q5zMLzipha/Aj3Us5ULPUt6lzzg
hn0CHLW4n/lLMC1DK6g4i8jlpTsIuJMurUKW16E0gAd8jiXc0OF5cd0mTlhLceoObWKlAKRH9Vu0
hMoLkXpKIsjIvXARUVbEE7V5l2peiHsvOawwpBm5cmF+/VG12ihYj/u0NFwTvJLpN1Wj+AtzZKDm
prJ6/me0WnqiRz02ilKnaci91KuQHQWLUNWcMY00yOJBZe7kar+QRs/Jfqpg+cIBNhii1gAPBN6M
NXDtYDxzf/3L4oFejT4Oq7fafcBzrUlDwGqsk6Zli9ABR3Nzmm7siWTdwSwE26jfg12upkyTu1BS
LvrQ/8xcXFlywmN/vxCZ8pPSBJvzFZ8J06lTtaGJJ3dGd7jVrc1D9/KelNXpPm4Zj26wlGsICWDH
EiwyX/7xv1QbXp5aJIAEpRFsZaVy9kqW9gSnjxO8cESfUL0Da0moLWGSr6PPQ1SMN8OuBQ8DNw30
E/sz1ehSMAaAnnNVJdz9h1iovaQO8GMRXm/blFOydYUwPuwsCJpHewsObEetOQ5shxCG8v5pdRRm
+msjNLldE2qAcKq3cMYo1JApkIVcFD3r6emVxnBrhGvTLDcojLnPukdC+r+NAbEGCLCeVmnwDEES
FUw/brCBZUsJ9OUkTbGKFi/fhKmJO8dfX12CCwabgIHRXLTmHXPlrml7lOSvAUr0l2Wkoq5hae/0
1D2Em5ZP7nK36JI+bA5RjxxWhsGoV6pmFuXTecQIv9vaRUABhAhx85kTlCYKNy6aATbjSWfVV5aN
UjgjdcPuazgMlurMrChXonLXNI/Ww4gxmS328dA2kKPyp9s5qY3oT82p4f8CopY5jt13CzfZ3sLF
f5oacAdztT+vr8ygPelx4Gqr/0Ld4XeeaGgJojW6dIEqRd5qEXhoR1yNLSj9qF59FgVOOwMETucy
n0cF9y+P+pS6Qfc70CU52WhZB70ONk0gu6zy1qQKXNTBgW0osE360w1Mp373XlYkYi0fe4pmpaAq
0R69GFI40LM4xOYptkz/WRZHJOpb7eAFyQpwJy03kHRh0Sed5Q88SL7ZtfWxxTMbqKkNVXDPYRb+
Hls1/vy4Gq2PFiXAd8bqPg/G6TaXFX/HvD053Z8Rij60QE+lskOxgVZrPmw4RWj6TXj0H8Z/b7c2
LDp7kl/kDUGinZhS3Uo64TgeBQWjZBKC6P9MpRl/JxL47K19zpQpSuMdGCf0jzNmTC+COIWKBDNC
/Pjc+dP/F7loczp2lufl+uyzKhG019TF1VqLEYVUXQY1qiofjqcGNTB4OS8ZnvxpJSSpGeaem38K
B6qcvOQgosp66XkG2m2fcxqyhdt4zsAcwRFsttrQLpVzuoLW0ad7w5WlyJp9UCrqQr6dXi8z0fW6
ehvp6v48T8bG/xaeQaly/1GGgyBnXg4E+W4KcsRobtuOnlIEYxBkr+j8tR5Zwfpgy46snDzV/o8C
DJEXgK/G9JdpqYQVbr+/Ha8hueVcYE4fWNBmnvE2ohI3XkXo9z8XgJBjQSiqag6TJJ2zSAEGHpFi
yfN3VOZjGM4mwwG0i/4EpLI2U10CrtSTflOlNy1GaRP4mAuyc15VWAizUk3hKRrpNkjNXxZwW1uf
UH7LwHziXrgiH/6xqfs0XCb8gRojY0nJjqW7yu4DV8d3br3x8miGPRXG9AddtWWchdwKEOL00egM
4xKVV1iv18N/OoPvDROxGJXhPtXiNKGeuyYd0JzDEq4114XEclaNI/jxnCiJ/v3wdnULSNBaTzKs
1OSLyM119C1YGee513gBQpYHHKqeQpOlglYssg7tFjcFbF7iYHSgZFa2uDpUZKJmcuA4AU5L664M
yObbWF/kjqot3JpOzK2jqClkZHrkZE8hy3Bce0tuREZruuyt8PpjolYxg5kXBbvZZAPyKBqzTVNX
S1F9FgvzFj3krV0MLNcqxB/bTAJd6yirl62xGDQta+nWK/DAHGvRyr5pIhoigCVN4MLHZSMaTY2R
DNKJiJlZiinyIELC1AvBSPqGf2Q1lsBiiRPPvTnXKbdsLvMB7s135U69gEV1ms98W1Z7f+L+YGiD
WBmK+OI9EG6eU1c8mRo4of/4Zh+af+51vFiQEt+x+l1zcjhwkiUY4rEu9cprirPu+ZijsJdivS6P
YuLgV4hnhBBGP8LlshEsnz//6vZHkFfmjt0jS6sMzJ3BIiUbI8YQ1s1GSWOXXaXY50tJ83GftH1C
Rljtm1/+ziRQlbpomFo/083soX4WazTiTPEuYBOUo1kBuIZq1ape9da7OqKiUs1Gz/qPLypbXBW7
w3AExcm3jFpWNYF4VhhhGDC23qPekAWOKzWU7rTNyJWyt8K30kIrZ94GcB/CCCv6Sf6Gh2tmXNTm
e3LEUtQTIhdeveVc/NZUq8/d73cMrVFbuxrBmAp2JcUIFsB5exs2RyowciHEMq9/OzPyBOrNE9YO
cRVeZ3m6vxyp39kaw4LPzzRX3Lni5nbwXukl3Wz/G2Wm/vHeAZ22QaVDY0WyplN2I7V+hxCX8eDH
a2TdEOirvFMtog1CO5FIFu5Q4NfPjilIGDLoDfLAbjtse50T0Se2J3tAFWdShuv5q6IQ9gXkusTx
CmOmWGtom8VLc8mHZpmqNiZKbkbE14Zet2lrEzRfFVtjWluZHloE+8IKAhhR18u7p8JGobay9H5T
5HY/lEmPIkUXvt58IfmUAY9TjOZubnkqd8wHiiEgPb6axqc7GjIgFdkreWk3Ffdp0t4/eaQCly/U
Yter0IQwV6SRUbfJTgz9Gu5Lbm7d+4fCtPnoc+d3cM29dVIeTVvHYDEHLFisaHncLxKb08gANtWS
siQLqfIOMh1Q2NrKTcXz1MvaL0IpdK0pry8zTqD2tbCoKWMgb3qGz+9HWNQdNqsx10r4NAPEPvWk
M8qgi1WfvQb2av4gEQozZzt6+VnyHwz9nvzGO9WY7Z6Y/f4PKtn6oETVMC+n0tQZlUMCWMvfP9Nc
ZR4vmB1yIwzTcBUArFBHMsnhBy5AVnEIthOsZiWRCiUyHejsLk2RB918pbW+3Cfg+B0HoWOk8Hs1
z4S+/s08+6GOjFblNYb4P+1iAYHRG41+koAsu10LlVj/Klf3vj1rNmfL9sbioVoxnGVXtgbDy1Rm
AxvSnO8GruMAeY7082Q9mW2L4PN+3cp21dYjyiveXIS7rV2B7i3tNB5+u3US2KBxGD1lWe6gZSkk
OCttpEodTG8Z7aHbD5poC2CqEVXpBg3X5USFT42ZhPmWoEfCE4jOVmkNo+Ei5Fi3A1lY+mYg7cAV
yE2Xz469N+Xvp7CouuB8LPaMxLz35RhRuHOZo4MsIA3IDeZJTAiG/hKLKmw7gzXngZUeN0Ffx7+9
99422gbiCbNzTwdqspLegAHeBNKH8LRKq8BmarFnLP4MVDPuC+vqsw+snk5bvR5DaEk8iSEtXVpL
ON34hdO39bwF22sXvNeTmdO4HPhiCCpkfzxFYP+AFfX/6n1iKiTm6bAXTsx5otpuctCGDld7m48U
eYxUVn1HULDqEAzrDA1hnWBLderkiXyD725sSnlaKyNign8ZD+kYVA1syETtrs1HiPHgP8cu36qj
25qNgkHNuD76HM6GJMd8LgEAm+PYMgpEdCbml7hG7G8DMyU0cL3L5MiD15+HWaI+1TPViitzWVsR
SkDEshcIR0JcrtIWC/nk4EjjCDTgZ6BzAYc0R/9J2PIKL3YeNnUdjsyT4aPfLVORx9rr1BOpTx45
tEYQXYu2oM0qEjM3CbdU1p+4W0R1fekk/nuCIUvELpWLoiWScD1suyAtmsKJlAjzDOYLSWIsiR1P
oqLodVjiT1I+ksTvkufxuUCbqxozbSWdKQZ+wqBj3iNupVgrUcDI2M9nNNfT3xX+vrrVtEyX0dvm
ue75zslzbXe3cdjbtIY38y8LmHyMdizbsSSa9r4Fpd3xLYxPnVXt9I/w1F/LLt4EW6ALjS9FFVCR
4cUxZdPFN0s85DrRQl2S/JdO2WIVLrH5hBRcl+CfBF7sdrokQEbZEa5mv10mR3atvJisdrbuApGl
JFYOaVD8gv/skHwO35XWde2RLKHiUj1rTSOVQG7HCiTglmFDWf4kABGYuVqm8jD4VFJY97OoaDjX
mT0gak7nVqHBBP7QtGi9w5iGTcq67k7Hkgdqs4KHnMnpSSRIyAi3vuOz9tTawygtBikcfNNXSgVO
O+nXNwHd2PEkpoghgWOWGOqwaizOPxkKxNZYRoeZ/v3ELUjM7mnFEH4lKhufVBenvdFT2CTaMuJu
LF/xnaVMOXqOvhPtEwxPnInHAp6yAyhUU/HTEtglGv9qmCVsoGtKjdClghahOdaD5H8dbLzGUxMJ
iFmKc6i0x65duUzpavozJesALZBCAN/tgbZGbXNXv/4jgShE1OY7zpJFZziJ7207IfX8VUkyYhOH
W3v7ZhIE3U8gWlokxlHKsgO/MpzSKBidFfg9kPT6+Z/ndymAWTpRct/zNloVWnP1gNUR6RmxMOam
zg+0Lm3zkQ2h0ZWktFLjFuGpuRFEInJm5Ty7OLWLqx4+jlRBKitC2pCVYYbCARgOetk2O0LDmxv6
Ucn09/zGLo2f9Cz8Nu3AbM6LB5CeFPpINoIzzR1cElUMWjaLCrLMH4ve7wmwC9ALex2DhNX/T2s9
WtI//0GIACTkFcIG9+gT9S/LBAt/DK7dVpsTdQMaLQiwB8oF23RXjh0U0965vDpPxwtcghRSYFhr
tAf7mSp8mD06RtjZ/wKf15u6olND2pSasZ2j5ytfaRsw+zTfvJ+gHsyZf3AnVmdLXYL4SM0xm7+s
Wfcb1GvTqN8vaMtAiX7J5M7PbTIT8qqFaCy82hatp8mtBXC4LGaFcuUdh74W2jPDqgbDNhlE1zMc
vYSZkSiL72pmJK5Lyi0BWxRvvP5KUgepz4BbJMfV3DcWRPjeN3eQQBy+1W6YrTgDjCO8OStXZTx+
ebDhTk2kCZpRzJyrxfzWVElfNVTsEvXO7u0ApeIZ+jQ9HgRyTvJEuXWkaQMGCOlQbBPKs9DqCvtl
ZZh6EhAvAon8QxsxbQwMB7QULXKfWL7ApfVHdtubssc6h5F4b0sWTSLbwxDHwKz2/P3pQgZpfIzS
RYbzb3xiGRcaGRLw+3tq6BldSgoA1GxxpKiCJrfZs+xexC7jaBDDw+Gs1jFOqat2m1/szALtafsZ
KgoTrAWQJcroxhdtRnAT0qHtMCM6G8JgZmbYyByBYbrqR6/g7MDjcBjck189fpywwRytHW8S+qXL
1RyYN3vp65MHUW3K46egm8gjy3cZ0ELEAtrTvSxiG+STtlLdbVGVkmxvEAsVCPKg28j0ZnShk1/t
ZbMuvsLZrAZV6cPqWhkynRDOtz7XdXMZDzUZsh0X7dXoPVQgBBEhdo7Gn5CybMSmpa8naVd4JcD1
X3boOmp0HsWf064y6rCXbxKqAAgOtycCr5gAXlOagbRtv2F7icxxqEGr1XwqDcxTiR7P80hmgN8u
AmTVqhVSkX49EHst2+hKtOvZC6E5a7xvODh4OXyp+6U3Bwk28FFGzrL4xO9efMujYkFsrc1ZecO5
q06RWvTOi2dEReK7fjCINL8+Wl2VX7x+dKuaSaPAqgi7pJ0il/IgmQNAZPpM6u8TRvMCOjvMmzhx
QRDY/LGvm8F/8TtdAFNSAdDGI8fReUJnr1p4mFGsF2QSw8BoDRzD93VEkjPZ0saYosbPhykPik+q
Rm+k6+Kc/n8DpkO/yBBip6jdrgyHycimT/YY086n3uHZqvUxmX3lP9jM4JJjkN0Cxp7BFGuAaItR
Uf6fwbLPLr7SaezuVHquB/uAySsn6HZ4ON69RXiroibgGt2uBrMbKa5E47f3x73FNdeIRqlWX74X
TasBNTviMTgpz+ZBQNgy2C2GesVmjroMj0E+k74NdZk2xvQ1dWhlxHFT1VqVE3Mme0R1v9xxKKYY
1Are9MYEQOejKfY1PORt70lOj3bt3kxoQ+oU//htVfrLRo/ruUHLwa3To+cqbkSuOVqUcIpm5XtM
ipA/kYHX5SSWHNHAl+kjFyzNuB/D7xbnbhyp15jnObA1sJq95Pch85Iwy5mCTxZjpkVetktgYMHy
c52z4jGLuzg92QfcuBIGlGLHAUhkkgPzi20gbnYitCgoN5S6q5UQ1/vvyN9aVKyjGgOm8m1iKOB+
4iHN/kJk6qlIMttnhbdF4EJCmHVqa3fxvNq27/EK1v4K/w2myP8Mg+siJOHfRyXyXkI3tCTBw86E
hIZT0jT+C3J6oPPy0dU+hQT7dTSXdmF5ip+ppGaJD4ZbdqdPiHQEH+FTcx0g5YlrZ+ICnxRAGjcD
9xRTeSLwDB1ZqjAos8FXlwNGF8vYexEpYhpiA5p36lQw4tiDZ4VE4Fj38Cfs55EGXc1rWYl2Tmse
ngdYaF+ep/58v/yUHknKBWHm4s4sGY/tSqcMUODgjEb60rv4lGPyyp6edrAltBUQegRXV34JYBGb
/M4usEiGPhuQ2WCgH3va+FFW5eYHu4JlIf9CiwBEwxvtnb2civ5t6ndcOS07Pn1kzulaweBwKZUf
qN/ZOQHME3qsqOH4Xjxp8V2Q6WRHW0ucjy0oFtKdOx99H5fg1aBHVoJK83Tu3rKSb1EhoXlz3gKG
Vz2fbmA3voWncc0tbYShOsKtZ5ch/U3pLxTGUpod7ctZ0U/2nsloY5fE8Z00Oc9m712XRS+M7JBD
+Xijk/iVXkhKRkB96g5BlhExJICNBxOVIfzBDTLUT2POe4GpggnzJdFpcWdbPYkTp8JgWXJNbp6i
0rWIHEMqaGUFcLnSh9Q9mMzPx6965mLS9ZlL90ztLEqvCCIrHKVKjoVNUWtJnE91Pn7hQDHPIniu
IjbAlLVTFdjMhOSQq2/EQvlu5p2cd4fapSlM5wxvbX+YUHlDGZzrK1q1VfPfgE1b+PcrVJpJwlgK
umv30DbdI1tPsdMxa76hwCiXeObPzmyU6BI7IHsDArbKGFDyVORykzvkt4Oe0B0622S12byBmv1e
lm42Oo36vSPjpwqROeuuXMJRLvOkLESBTr1tnT1onzj5N9f2HB38v0FLdzuaLDdkB/HBfrCnQpzA
bTX8W9kRmGErXIjkkQGKEpq4f+ddgknt1/Ib4Qi7urHhs3sR8VuQMCQabWQHBX9puB2n5QFbwtRx
hufd3YX/IPkfJcwomi1cAuXQGXpyyEcMITWUinyx11B+nKUgXDG2KgOrNJ7bAP8kaQNCFdY9kUd3
S5t//EMU486yevWgL/f4GG8JA0crpKOIqrPKudWQPWizXJ/j55TaBpq9NHu7U2kmlL4JSfcucxql
SaAM9v3yYx7ZAqIT93RmFXYEyiXthrU3zBL4BgUaQCHkJ4SpPCKaYaCfIeqD8664EE4g968e4olo
rszVOIDlcfVyoxRFIBD1/692ZmlK1jREN4VAy9LuxMoEAJPcPAW8cER2AyOeNgE6RUyQyriGVTlI
IUzP6N2p4GcyYfZcHWjaZN5hQJ7UPjm3iUcncdcEl2zpbMZ+1/2MNfb0YuIvCZ0tfF1V/pMgElxh
WPLH3J+sVgPBC5H7Eov8tFwDoUk0zOHU3CW+u4F8jr3w7Ta3P/wsR1Zuxmy5H3OJUfGgvvDb1K3k
ERy89C5DjqzDGAuCq0DMIg22AoXJ57nyjTJiiJIWAJOY4i9FYLbm/WkQAOSa5IWRw/75oTLGt2Xb
DicmT6TPeRs1CJS+rDZafjkCcLwxRbLx0ogHTLNz5rQ7WnwETdrtkCbReGQQV1UBq9lwVW/Cbad8
j9CEurQ03dntU83bFRrNeMLcH0va+z1TYrFkcgaHhdEN8hLpGSPt1/K7fn2qXa4XWnVv8rq20F45
FB1o+FadsfEQIa+WVlm5QEWtZEcNVLUc/G9ilP/+GKdGb1fW0nHvMgOBfqYfeUr8YfE7g5LHXw0n
pCGW+0/Jcc9Tf5rVvCnyyt+rsQGkhYGT458LvDKbA8oAU1h29qGLgx8dwOkj2L/h1/yDbYmeUp1R
yebDxR8dD4F/TM8e1elHdiaydFTGT53BrUNs/MMOA4Q0fFov+VrTUebknIWbT1fYAFqd6QBD01Jh
vLKes2/UcjiDmeNrhdTgAPKg0CzD2T3rTwodZCi4NJ7gPG2CtUxBDFAugI7UeYdKyZpuJXtRjJkQ
THz00ctb/FvX/i+kfNKGMIj7W6Nn3VIAz/JeL8D1hdo9ayWmztI63cA/jVkoKpqpoSIa6+nu5bvC
2HA9+W2j3t4PykM5QRz6UFuIbhGFM6VjvLgYCcnMNbKAs9Tiws2fYxCPis9cWKQWkudzq2J0fm7I
n5tGbcytBBwcuquG88q4ce/shZqdp3Ju200kx82HiiOy5D02DVic8XybwJM94RHUtZTgCGbP2ULl
ojmer96AN0oisKC+sdz96yrM5h08NxuYzzkXydHzy2mKClhiNHZp8QoyJe1FI3OcI1cbCnCRo2Ov
7o2irwCWghZfrW9T85EEWdGnpYp7idMi+phu+ZgdP8H88cH372yicDtb7ZY9Ry24GztG8FLCe77M
HBI4+bYTT/oyBz8UEQI7I5awfQmIiW6m1A1NVo/cg1nU+4wFFlishCBKkZocuLCZsJsWUamLkgEJ
XUZcLbRj3/VSxZ8YRaz2qksCDcrZSoZoTlbbYepwiamFXUCwLZVF5Lorq1hscNQ9BjFqsRVMe+ki
vZXnLFtfSXVtox86ROGIz7Ao9sqSg9uNIpL1zPKjNKbd18hmOwtWhvjPcSJTM/2wvSdFAOQtsAl3
rwalhM0B77EJgSfkSZ9DXukIoVrKzfcIj8lzvtXiFARBtVpg+5isf2Q2pA6FLCxTF3uMhPLCd2I5
H8Q1wCDleIVDyolW5z0ORMNyccuXLvDh3R/NWkcSd+TTcVYUpy69RfXkGhi7/AEhvtEQVQDZE8iv
0a90o9tmBYgbJkzvmIV6eun+/Db4KxSUuEomON22I+RNL0TUNzHiJKmhGQxWvNFwf7tMEr76d7vJ
nBR5lHY7dS4TdfFEMN0FB2u5RPfRPMS0gxwEqNpuU9pjgr9meJblHFpJxzBCgn7/3fJMnPu3m2f0
H/3ZU8340ltN4kzAFjH1LX6XVIXE5fKi4GBZMlkrs1NaS/0Xh3A2ToaJqHw+cJr072oHfsmLN3rh
8Y96xuO40hd+yLEsFyZ2d5QEkqPRhRLukcIP+b4Fp2El/qFsUT6SCVWkXVLaLvYGD+aNkLOComCf
icL99cDZ2XKe0orioY+5+acksvRBdyagDflyjFVTKtFBXWZxUHpjNAbHHlq19efcTE8ejhTjQ9ks
gCC0kGe0Jcl51fBSWxrWV6P1UHwdO3t6jEvfVb0Tr5Fu1Anu+9ceeKnWaf5R6WZatQB3Z/QmQNIB
z+N/aqo+2c4spkOjRtdAdpHZ+hWgh1zLFMP+m9tE+bVDIOaQOLyuqcKYnzsDntKQ4s412kNBEDvB
pW2a0hsYNNhaevHr3ixdr8mcYOBfP4MwS5Wf5G6yzWwu7SyFxBfVAtmm6J8s/Aj4f8t2IqbfpvYX
RkXnMNmLmOseVwbGPJDB7O/L3rgo0k1UoIu5g8e29rb/uRIgEe6wmT1IuHkOgpHYie28amd7cP//
FqxcAi1furLwrl1+l7U9Sd0rFFA1kbKt2ATu++rxN7r3CL69W7zNof6Jq/uMq69i1oMHnSv8aQKO
oJYxghPEZE83Zve4cdaf5BU+7WRxyYG6JeniY2SB0IxHtYDdswSuCk3TTsJ3xToPWZmMIxBfY2qY
3uLC3cbfZn6VfCflGdBF+aaXc33BeNllE+Gzdoa5SqDPFusfIUrqiQ6PJPLT4r57J9q92yITdKey
NZ3WJ2mZNyGoAF2zYfo0m4rOfMabl3FW2244Y2sd3bgaktvlNeNCT+p60h5trZDMjgJWigLiexXf
FxnU1+yymeEEgRWfgS6NWtrKnSQHDhMdJlDr0oKStCh4CpedOuEc57V5glSuTUpFFjLhCyKsgMQ2
0oI+ozQNYjxkUCud27Qs1T+iexakHOCZcqQILsD0oqLqKCjtWFCUxsOtD1hSxID+5yJ1JiJe12kK
BO44wUZEZWXjwRUuRUrw/A+5mUIid4te2DkKtfuv/VT6bg3mlE0TEr41lOOU5Mtq8hsULaEWo+x5
UhcOZqm42opYqUQhueb1esJO05H/8yHtL3jRkm+/bLzE/loEH71dJjGWAPzzjrgMDfMlI1a8r2os
/9v3hD3b4WfklRlONNgmPW8zwTu/thLrNk3JUFqm17DXQBNMr1Rh6wDYt/pjXgueDbjEJNobtTOh
8HK8TMmhVwkWANhjUBOsAeKRik0Ma/F7i3so7/YkJhmN6Ozx32W7cTitbSQh4P2ZFkeNmlAek25a
sxz/ZQXYDwk5ji9hn7owyysUfXbzAvjdb/JX6Ut6kn/k00vaZzQ8bfT88Wcw2HFzOf5prD2o9EO0
pPLgTjoYAHi9MDn2g2vBXm3DYQO25rDkYMMBI9r9cQ8mZMjfvnPMlOs/eQHvUET1JmVaUjXzS3FN
V9l0MMEZPjwjdQSzIJjBLxxuWNOvuKIQYZ4Sva9U0EOseUl+/rjsV9j1T61SjA/iDAXFOg00S7UT
hzZTVsosHsmJLIhS+9Lp3CJfP6vxP0O9ZP+0OH6S8cCRbnMjsGY1nLVdfOkzQMvGCb7SkyEDdWMZ
I3jlGCHb4iT5OlRsLaKILdDwJyEIXxRwNGLL6I1RNRxqz98jywlHly4hxxv3b3HEFxFtRHsWZiBx
2vetTsOl2xLBmrPn49XyqRlNFi9OvsC6gsRbdoxkdcvESzAkAU9xGHuJHbNE1EiSERp/6eqdpOyZ
0eUVYLDwXjDCsfFHQHW7JMtY9VUCpfHqwWp0Bivi5IOFva27y9/J2+/cXl9iPE3d0DczpqOMb5cI
yvwERARqRwOPxqc9G3pwRMqvIiqZgtCmowidUz4hyV54/FUQbLORRndp5LYX4P5qbnp95QsLIWW+
LFhemn7QPhENkXUnLqJ4ytpAgDCnPpQsGr4A9y1YuuXF5zOadbabjirPuDXhdJnzAuSMn2If45kS
MqmES5kSOEeE3dnChDc1NWFd5OenUCkgaiRVR/7xn64C3hHsgGGKn2hGEhM3gVsA/d5oBRjYgaYY
znWZEAjiNsA+UB4TrowQ0CyAgye3GgED3J3liIAsOZeJo8vuIX+68/MuSbVdUOS8w8bC5eSZoEnQ
aVWh1n6/aYhgoq+IswefnruNbkBcRWFtpk35jZPiXAoc2iKvrr61qgFQkvX7emRgg3dPWOyN1gsT
QuTF2VW+iraPosglAgPb98m6oiAVsDjmuErWpIweWt0CHqgz+DdlXQvt4LnoMSRzecOy6TWY7A7k
VCX7Ypl64IWJCT0Wfje0hPRucr1LTX3q02sB14Fk6OCPQHU7Gh0zluVGkn2sUJ4qjf3KVvbBDl9X
aaHhDYICdZzeQoPU9+hS7ATMU2oY0xZPdIb5My8Wk1pU4xOPArXT3AEGUTAe8LsPyZCHwEI1MLlm
DioCumbTa6mek1QxirfjlIQU03yoAsdPioSGruheymg8dffUobTJee9vcwh/GgCbYDRZXdpA2dQo
l8+gdPQmL9bWWPvmIW/6KViYdorqwzs3fwC3pqptxc8u2/k3LxueF0hgjRQVdzd+otYrATZvBzbQ
4ODZaPZI/vS9EpAqgCZD7yxGUrJj+MhvQNQrAXjWVu6gh4FSwBv61vdSqVi7Qhx84x+dYqUtUydd
GUD+IQ8jZvYkAlo8OSrbu//ZD0Y8wQKfXuUZzQJwE+xDQ2SP2gt49Vl9Q66epuSm0TqVZzis3Ikp
Yw97ru4VpZSBf9iZX0C5sovBuHWp4/yxVYj40f6NxKk94kztc1nmKtQliXJsUYCZsnfVSTQi+8zN
m1XDNGpFCT++D54Pena9cUC7lquH+h//NItErNZDe90fhMbxstsL8IszlQSFxia2Fg33KGN2HxMQ
0TaCrq3I2fGYkQbjROy4AKPngKyDYYCjvGTKAbiH8CUvcpusry87quFz24k14Jt9So12AX+E1ZK1
XIGEdAD9sQ469DmZApyIx/OKxUGpNd61iiKxXk5bwnDGPISeaXGB3O3pq6s8iRMYac3kMT1e0+H5
CIojIOul5Ti9hlazK7zgZ/4UtBFLcdrfhw0O4zbMBD9IPRb0NzBhOeJHJ6Kp365IbDF5zrRyt1QC
1GhQkNRffC68k9KbVuXwTa58QOPs7lH2V/w7kwNp9Tqs6rX4q1aqgLg7KTLZ8mqVzyLL2/Eu2MiE
yDfBNK6ngZmsm32rYWLGGqFzrJQY4EMbiAKfJqiH1mHDOrv628hhby3RJCB7RL1UoY4qrwRq6avh
RFvOOiZ5flcDG2WIR98RSTrk1sA2coshtc17TaCtJejGcskFosLj2dknIY+eBmsVfEVB3CXDX2nb
lPiemaepgl2jEaPLG1ZG7uLCwZG3bQpavkq44lySiStIdE3zC7kvZgWGxO5lE0Ev8VfVPnycbQdY
/lP4jVTf98bwfAPdRS/dxAmpIMe2df4T5jmIduFGhYL66AA7YoMJSVtjlBxn5Vg5vJiNOcQ3tKmJ
esyYEDOrLR6Kd6ODmsvgDp09NqJvW7v7Gj75ADYxJcHLBRNwQOXjjEe03XsRh7OZ5J0fiT4BbGAU
MZpAhfJuOXTvIY+OgUnQTyULja2W4G7OAnP5lqMUxJLBHMskBBy0m6Exw5JUGnnXxQaWitZpjx5/
kl7P2b1R7wcM0I90QK6IEX37210Cp1glDXcKWolSKq+ZkIRiQsYUgFPbtLwSYIAUKnp8awaneYRC
r2xcUYachGM0sYwyqCiNZFe/QeyRsCAFx3yIjCij/fEDj6rJ05FwmIMwEDs0fS5/Af8qX+g5kVsa
FF6y95Ri4eKfsibZcakuv5EwHa0wmLcY2Aphxx9vLlEejFGLqYfaZsblwiwK5v9zhBj43Ydw0BsT
hmhTP1w0VJQM5s6/j9MZ7H2qeKPT5wFMu7lzrVLy5XRBpttht0jjsGJlf0ihDKLS/VGh3A1ph+RM
8TZUNKgccSn0ebJuih0THhD3jrz5K+6/xeU5KUysRqgTEgvK8I4a3Ygr1hfJmqSw3zNNzWueVokO
ql4DSqZr3+rfSrGdOyCs5Sc96sBq2ebJrG4MsnDpG+UVZ/vpAsL26XP+y/HM2Ewo5KsfSSOZKtE+
t0CbH+Gdn4KXgV8+nbluREvLA4H6AlKOUuBsRFuUe3++HWrskunPoPATgkFfnedvQTrxpus0YXzt
kNR80BjdToPwineuTOvWepNH3+VoLaQSkyy/iUUnEJByg/Q79g24c89h5yUeUsG0j+qnoqvpcjWV
6+l1GbGuwRfgduh49Wt245VpuLQvzD/eg4pGs7X8EH752sP8R5PENctOgalrg+1QCtoWrmBWuBEN
8kOaL8b809nJsRhc5bdktw91XDtzo8BTT+kj1P/g067nUdeGqJKXTFBTZHEUkumIojPIlh9X3foE
Trt7Nh1YJc4Tu69g4c6qEoDrN+yUfjWszpQ7Tdj6hm8VU4n4t6jlpKcy97tThIgwlQiAbVyIQeep
eDpy5qLtVebK8BqdUTfvOVFZWXziM9bmeIuhkvJCnL+MwVpHTsTrw8UNhN2P1fpLEbu7rxKafJPA
11IudmXVLk8jMNZ2FtetE+oFHN3Q2KXSmmbAHLSzhz6VH2kioAxw51mjcPAKNR2PNfysjgQt/c7s
o90VcjG6Km6IG+wdmtNXDgE+MagsDmIajKmGq3bTIdO4OL4t2hOzN/FoKr4xv1KqGtPlFujM9Ad5
fTPMw3CRrVr32u5sBoAusaNlB8yiCyHnNLfeoXODQq83mj8HZWlYmhNemgR72sMPHGOMYv2gvKlr
noFxO5dhAKurm+1mndIhG1pMzoWZwvm6MYxuwxmBbOXN1VM416/Po9hh6jwiPCg7vvlNEyL+kZFB
UEYzkpsPT4YM/3mDqDQ5d8wi8VdUbmQFtkUnN3RHFFdg+WPnvmtcnkXh1y0Wcq44MQvv0reHV65J
XNdXGwXILFctW9uLCxCCqU6oiXs0x1ydAMFSlItK/0d22axS3tocsxNC8X6kWywRWDbm5WCY0DRH
Gp6rPeWlgrvzZ6s9pv9yeMNmrL5DrbgRqX1bFnKDOSGo8JTgRBPMgJEb2/JDIfGcb7x3wXqEx4H2
aZgcMZ6mu0POTvOjh9psjvqK1XUE8fYkftzMN2SEs6AANRmkvHMdlUrNjft/kmjdY8wJM/reiOF0
i+WkPy6DCKLWjSSU74eNXHPW6DshJ86U0efDEws5qZ0iq8JSvJlJmO/vmwwoyrLIJNKh5zEPOFHI
VTec0JduLQOs+Gly5zZf7bgzq+Nl4mwysn+ztpC6KDIYZdSfwlPQ9ACao24LTgaJ/80FXtIsJgo2
PAkQ7XRa3Lgsg+8KrmvpQ6R1xFtCBmB5qL/SJgdIOA/bhegkjRGzVRF0xrbxprzZAH0TktJN6VyG
K+h9Ih/Ud3ciidVx6hfuqHAL7ME4EefvfWkNKRACF0e0znwzfvgCRDhH6thPvaKCkoRPzj7pY6SR
yk0DNxhPxg/1YnVuJJc5nYrUX4tn0g6VvBf8tmOdOyzbc6+QDzHnkk9Pz1Fus8Dj0iwtYpZEc01h
8xGZoe0sSdPhlS1oq2kOEvMTE/VKvIO2h2nGOH3r7HdEqikJi3sEnoLEY0hK6611Ikz/r7btqQHa
4hZrxp5qOHKmcdvyechWYOEdElpR1HnV6mi0/J//JoPPhrRNXRDPLvAvSszvwa7hXE4wedqldHbM
wYmhOzD4Ce+h0YoHtPEVqLq6PsH4LqLbMxc8E94yfJeUnucO1ajFnJKCBa4i9gRWzox05Ucvwpjo
rtg85OO5ATOEpkKlsysLrGy6dzxC6CQnOKGLyJ97uzFVszz5vv5aGe15VG5fdM3Lj2f+vVBETwVd
ESMZlovFTpVOZm4LMHkyhTbaPLsZrU2EwJrLDmRx9i3Q5T/reL2aXclXgTZV/FxRjVkHhvgAcGBd
+hz+4EjNJ8hSCe+4eAablk8STnW7xmPhice/RLqYjNR3JjRDnNbmJgISnQ1v26jbD563HTyLKbCe
ps2723hVyaPYDX5NSX+m+rcf+qrL3dRsls3sCbtmytMRPgsm53roLOa1XywEmOx2qe/kPqSffozr
cQ8DYbe9itjCkP90ejcHva2LG7smZuG/10j3UlWoMli2++71S9tlC/ZrV3BAp+8oR2zhlliEjBdc
hjNupEiaWnhAec5Ujwj6EpzaW7ppnVqftW/Oo7Ljtt1EOwffOxqM2QbxThUFjuCmI9Ick7ZoDUdJ
vPT1BVL7V1bUWkckVx6vu56+U0eI+9hoqtAQTY6nyGhePU+OZUSNnWc1XpckqkD1vGtmw5t5aANX
YXVruJ4QZWq9vsG+xI/c/fdt2he9ksbkQRUHbd6EcP61bpSqYrSZR3/so8y1DRtZt33a6DWixl15
pFTFkOhTiPK8RHA12I9F1cHgJK30/6LebfMh68tg9SYVycISgqqzIZK5y0XkdUWn1YWALlW6IpY9
zJDZ6GhFov486vXP4XwHagsf0t0Emy0Y1YoQ8XLUSVcuKEyKMD007nUtZ9q2ppskiqemN9PIIYAB
yz1Z/tPnbNp9RySXTtJ2uJKOyaggNt7/WF+GM6x3jrlxgb4/p8Ie2Z00s5Yw2hS0YdrnKAb00AGJ
w+o8qx9vsbTvRCj5lv/LylLqW9FgNGZOOXwJ6YtMwt7pc9e7eufktn13aLrRRQs9mbrmYudKQBqI
djZepN9yqVc4SmWnY6Kx8LSfWpO9hl2XV3TQTMG4ij+BnnyRY2EhvsUU3T9hB9s=
`protect end_protected
