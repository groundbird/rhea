`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Hpzw0yuekPMh4gIVDJLyDCqeR9qmCMxSdTHvotLPB0OrHsADSFUUk4cvnaXTxlcNUfgTZWLtreP2
JPz6Dn6Ffw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K5AD+RSNzChCqQ86wq6Ux5cPGH4wsNYOSud1gimdrAVCKMo8THc2RG89RarPqk7WGnbumYICvVTP
IQm/7XK+YY1YbxqzsAhm/czL82YzgCqnTtuyc+AcZIyPOwNKXZSlSMHIGBRWSMrjAbpCRsaQMK3J
KzWkX49fDAlgDmH1hqY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H80cOS/i7Jqen8bUY7hYsMwUR4eiUmcuQqRvD6Re7MOGPxqBsM/xuCCy6RVLIDRafhind6F+w/KK
Ys7z/hGr/rtKFZVMlbClS1/Qvh04S0qxtFvi4VIXCt5h85SZAfZRWzkHNvBYdnv0OZcdyhKq38dp
CjqIqpQkpZPf9VmG/NHMxW5woMLnQzr31X8vJQWBH6UozXTONLt+rKw3NjJwvSEJqueKblnh1ix4
IoJDleoqoG3/InRZLYcGX9nyPWA8bfbxB2ohZt3cdGZoaxJpu+Hi4LIy/UD2uS2zdoIJrtysSD5u
GnLtaScpZyavWfCvn1WO+g5X357tbUr5D4uz+Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t5RQujqOO95yZKgYTrKeMKaOez17xVVUEpGSXDRVkWRUDIqLzvConfDl18fDK91uUbpvKF5HpHPD
i7hGCZ+o6qvt+w/cWGCotAFazzuRr35udxLbntFKpAUnRup6W4d4iu/lPzbobj76kXOo6aL6yq74
pVG9CdcUIhZGM3aX3f8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U7HdC60rTWhAGbdC2/s1KlR5wsGp8cP3a8J7gM4uDVATK1cF+bE1IF3paj+AYDe4XEER+ENCD/A+
JO8xwEVytsWPFnJ900x86AD5Mn58XrvrqSzLga++D2jOjmUccjUfvXXw6Dmub28RjHZMgxGz80R/
a5IYD2yu4TM3tGx4tlYXHD0C3TuQ5sSqu5XVCqkXy9qR5WQ5HA5Jz8ksTNvpviFC9MmAs28G6bZq
5Crdl9T7S/5GPalszrhLAqeHchwlz3foEHS3r/IY50Wnu+Gib+Xikt8rX9ssswxR6fcto4dCDcrZ
qSeL6KIDbizTUaPhfhxICuBvIDz4FCSwOufWug==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20448)
`protect data_block
9OAxKFAqLwbDVSVBK8LOFFsfOCQWN1Jc4eq2VRrH+iut72Y0qwyFkEGA8iFa7U0kgRsoSg93A8ZH
Z4qfLC7XusneExbdghXgKcUnCBfGlTo5LhDb0pN4CjqiFYEM4fgHGTj8j9qyiO4eOWtyzCUgvTwW
J016rsqRwZ8lRdhgy7eqFk8PKyaPwg5q6m6jkMQ6Tz4oO2l9/zpCohLY2QobG9W/83arYd+wy4n5
MStcOcsJHjAj3yn+WFQEDJ2THq9BR/NFHc5e6PkbKqA49KGZmAbotNzo1o1ku4YS5B67l00+sB6B
ATE0NVEULYoRwhMgvhWf+xCA1PmdXSZCqGXlA1f0ivHy8JybSiApV3NhzTuA5VRpuKauuvpgdArk
/KvBST/4QROZmO3fIhGEhFaDBcwV+fSyNYxsfRRTYt6AcDpdRax+O667uFwhXjq9LbIkWqpDXwKq
RKpkX6J7yMm9r9nB82mRaANKXxxvk4iORtQEZx6UzZXs0t5T8YIumxiEReXA48TFjl2q8/ZODham
TN7wb3mJrW9STsSWNB0rwt/1XXn8vwY4TWGqHo5Qep0rlw8+bNuMs7bFv095VIguRFw8tMk8bflK
tvQlCBfHRUG5ygQdsDOPYrqALM4yaWfKTAlXzV/K2hGZuGCXWRbUQ9cew9ZlYU//79gsBKI4wN/P
JoCZ17ujAn+6jVqOl14+G/GqunhvVELjPHRTwRKgDl/yPesQ5UyBamaocUS/BpdByU3UQCdveLUm
EBsCzuku/P3mpKV4ZHVPGVKa8CK0B3rzz4TnP+wk2nrMmFla7j3br2QKXsNR+UXkyB1Ehxo2enbg
c2atajHIgIwg+n/rc8haUKhOD0PHKP/8FWCh0hnfTKxHj34WSM/VadQg8/EUb7ZUz6YYey9zTWAh
p87oyqY47hyVfLpCgr4328bzJ0NYnQU3/x6C8lzeaC7xUcs5eCB4vh44ZegrufIGTavWsZHG7ss5
+dAvlf1sx0VMKA3W77y2VGn1WNIgfwghjwtTuyhKYgdhDMV+O7Citg7Z07pyHRY+FGrP/TNH+MvL
n9tjXCKptkhR2UdvkC793bwKV2RmrpAPbtSCpp7Q3L6e8lVRLdXinjKb8+FjEs204qeYEot8G897
yjnGBOPepAl/7IJhGhxX013h0u9cgSgjWebj8wEYFg38c0hEbsSR4jpL+0JUunek/ismd43ViTRW
GPHFY3cxL32l6FlOGLzIdZEzjDeH+QbpJX6cKBU/wOMd0b4Xxkr9DVQKL6yHk+Z65wi63R8hDBnm
eqiGVuYFlbkzHuVQG6H2JPGmN1hQQ9O2eXGJFy3sRivaJo/zxnclR5gC6leLjd73RWKeeYKtyerf
VfHKtUZPrkC3gwvH1kZQkvhV0Qncswrspj2nJUqWj+y67HkXSWsQ5Pnh6zJ33jTayhLopxtWqBGg
/Xh8m7yb5FnFKIx22OooU/UEH2aLGG/Zx1VqKS0ocJX0inQpGygOq3oD4BysI1wLlddI3egYD4j+
l3vWFGI3CVlqJ39ofIUXg+5sSp7wSq38hGrXrVrH/JZi3y8Eeb5RbNszIbFVfFAGK7WQJkRZA1u3
SJvePqcME81IXN9+AExTttAODrGTmRiVBisNSbIzHNGdxCDPg2Y4xPu/YsFfr9SpfFksMm4U5+ur
qHrJwojlAC8MCbFzy/Dmz/Oet3gjwPLn75MXBnaMqUQbtioY0j68nSIVBMnAlEJ3SSU94N3CKtww
77yN420YOX/ZSaSjIxv91Xlr3w16X27WyupLz9mTBIXj9ke+LLKErEkDOor+KRXczlItOPC3prlL
YrC3+gK0yyXNRQpnHBQrSQgppy5dMqy9VSy3YWYwPHPCBVnrhEU3UQvx+SKFS9HwtlzP0K+H+Yg1
KzlxCYVUmrqhfIfxkFZhqfnzI1EiYU6rBapbFAdE1XacmjlbzLl/xV+8VtQTgkxyN0/sT8JiFw9l
Ps4tENAd5FhLHUvIk5vJsHCDvMJMmQwQCeeZM3rgJKdZQ6oxTfge3DJ8p3h43eKfS41LeoMrJ14n
pfbonfOM9t9af1M9IHRF+1pNJDYXUob5x4+xTrNlhMtGOsdo7RA9Hn+3+vUHbF9rN009YJyUGwzr
VWcpPdhvUvJ/N/l8wNn5joq1OjiLSMFWzsAtx5nh1/ndh9CLsL9c5n2MmFl1ejlr1OFQZllO6FDk
IifVWH9q+SvduJ5XMeCoYqgq0VAmSaGNH+ptF274Z4WrUZ81VOPch1um/yyvzdt8PJmFjjvu4TP+
LThPAp6YOF5+yx2xnUpBC4dsTimBXg35cw71p1G1SGJxe/o1kExl5zACjQws9a6MxjDd6xYWKxyb
M9/J/6tFsCxMfY2nw359AnnyX9FefxDZCKbLwO3DdBE8+wxPyF1E6sQaktSuLPw2Q+WuGdDwwIww
rV8gBkwNFiqx6drFpp7rKcuKjms7sgXEHRdtfP0rTzyguBdlQ0IY6V3lnelfjHRGI4lj5viQP1+8
cNnHaT9QIu/3AJTAgLbUaRlEbZWep8DFMgEyLPKHTEi8w/BDdEd6FaDE2ukWWRo8qMvT+K2O59Q0
hfwbHErsN6RuEEjLEf7OgIAY+0OjnyEU88kAi5KejXvGUN7ZndI6GYHRgOjkHw7A8wWt0KM8momz
jeO2HI+SpzD7BD2Otokn4MYcj8gVfcVAufmjTgyGFxjfCEw0jrMWhkNdjOIQb2a4Z+JeKiOSBw2S
CWN6ULVmQra0J4qiTv4JknP4rgDLWIjew5/odGpXenK8cN2GQotFZUXVPWsnZy2UlKxCcQTKFFQ/
VQMEync2t3wJxdT4pqdGsEy1DuuZCrvKzO6FMhjhFPmOb2NqDTrSnhUqdo03WQAS1c7NAsKRwdQS
bXd4PAVpGD44z6w1ygqnuHToAJrGhthpOwQj70tEi4dQ2XSUzc10tjJBqtI8NfS8HZ5grwn4RZ33
MnrKaztY5/evAibDNLGAKxvKiNxRCFQnTmQjndzsduygakN4HkmGWD4VX/rwZg/4aGV4V5b5IoyY
YMclpGOdR646NUxu43lbz5VZHt2N9Zyn+CvH+S9oH+9jOaqqqiFlpp35mdAAq2pFA6tr9xpLwZi5
ybipaKFPKFcGIgY68HEOhxos3FxaeuG8IsVMFJ7tg8Bg2ttBaRVfkG9vDUWylRCywtizsgdSMEDx
3y7ECyALa8elN6/4hjrJubHHY2s284avMSNgL8ZspFG0gpQmGag++3YqtEGYNrgj1gBvMMEm98iT
2uK4TV514ei+xvZ3dIjU9l4x1Q5A8gXe309blPLuphn+5e9uAFgq+M/KBL1u3kqhZgFwYM2ulifI
65X+RzGfnTdQX0uQUkK8SonUF49VM5BmE0VIyik7bKP2xfmZQXyThF6rPY8lYdnbrdmtcDPrxFea
0c6owwmvzS9LhG4FC5gIjrG76pdY1oxsKDCGeog9nzq1ZoIq1RGXuhk8Rvd80AKQAAczjGiB2HKq
M/+wjrBgyTZkMzrsVroNsAArVzCENPiajvOnvtIehHberIC5HlQJBfTJdW3KgX1y0TIFM1YxgGoy
9goQrf4U0gyfvaqu8ezWoyf6PPiXhC+0MlaBjvZO38H+l4KA9V78rjeosVp+a8GRqbwf9LivOM2o
b6vM5FnYAu3LHHVrvh4TqSYxBqZURapFIb/+qgXxrTe/wtoLI6t1MIqzcUXd4GpGyZj86Y1YDq80
y8l4ZT+UUgNOfHvM7uIeLrdQyp6NQ7Cu8bWcDh2QPSSr0RETGBQfHKBzpYPblBmJW1vZD8E/UbHX
VrCGi0Kiq4PPSsp1jn4HNTMzvsxK4RRVQZatyd0MyBOweg/svPcMf9X1aPwbVYpsGxG5j2aL+Kf0
+ZWY/RUtnohB/ajvTvzMP4xFJSE2ZHJeAFiecPvIs5LBx+1rI/CEbzGufIcVfyTM2KB0MW46romY
o+LWFvuvHgDCt6JClaDMgi8csm2KXmyUd6Y5GHuiA9QdbM08DcoepjLgQc4sn4VveyMJsRx3KLrr
9sY5XDZCif+wwQBKqHaqHMLsNn7CySpisPFkonH7AGhhY+k1/+rzsMOCApWgKJxCZL3Y0o2tyrIw
h8gTxLF1Xr0oO2tHVbrGSA2VJ2Dg2CL6b0NhgnCu1utTSmSCvMnUC/TwORc7ZUvmzsVtGzHLMR6U
0V+G0ZXq8KqwQw8609nuoKMxkGgG64GvbR1CWXtXtUb6powKfadLDG/oteAenUxwfHRXFMGgqDNS
c7RGv8HoTraOLsMx0Y2XKmpUTrqfSSWWDbWiAu1Yqf4KQZr/dotxSrmHhB4C2OBkWB9WHzsYinWj
IB4QfBeNfFamRTUZupmRYlhvo7yzFF1RULCqrLL7ySrmjUFlwlDBRCahgd96CqJa/6KVMx9NpqSV
d4oinc1IsTyXp2nahjX8FYQKIZORrlKZhXFY8WjbAhAaK2ymlz29rGvh1GkHXE8+c3dIv3PYjnKQ
fXr7+8Ii126U5NClNEuz+kWqOMZ+OhKEvex4ukeIja9B+uJd1n2Szoi3ozs3lv2EQAwT00ooaZsR
62Ry9bF6M5srIXkwzeQLlUXfaiNUd/KegqrXnBWQRrI/P8LykcmQCVsJp5EFt4SOultW0taLEJDw
B7RJWWarTXKGR9E1/7AgHP0Klvu1KNzyfF5iGkOnnIPvwRZ+nDw3yp+n7mdG9byDNEYfvnCwhK5A
dOvHk6xVxFp+vnNA0KQdtOJ4jPVGhEGb4AAQBVnZM06b1Y1+07sEn2MKKcp04nNTBA/i0XRhgi8x
a6+JDXWrm6HVGGyo4hHCtNQxocyOomI40tbNuvRXcRqTq7yQ3j/mAucQ77NzTZ+N3J+7aMHH6Wfl
64cQ+8xgcFIrc4zCcZMIek9d/3pjr61NU0wT9012RYfGbGqy73IQsiNKmWdONgUE6hWa4fgMyVe4
ZnUyMLswO4BxzZElWa2ngO4afMN+U+9yPS0wB7Wj58zsZ3o7q52pbYKZIuaBNU66ZI6rrCJHQ/yR
QvtMqADqFFmEQy7ooT1S1WfKZ6h+D6yTH9AEdpa+TIFBxZ3x2i62FPq9ECeM3U9QTrXFs01RnmRi
QV/AfDDi9N9bl0Iu0ijn+z9K9wLbfgFFY1MYGZ4Tw7p374So+kUwQqZnsYPUhB0UcCwzyLQuadqa
4ivGMIY7GU6pbcfCz/AEcvVqubrvD+hrQFKGO3AflEHyjDHnQxSdWgCN2W1c/0sRRp0p0l0haQrW
4yT4IdKTDc4ZMx9bCoA10qNbFperUdHQivH4TNpmqEO8QzEGp1ZQ0ZLmLdyMSdoUTtB/90poM74M
X7g3swvr8bcPO4ZSutUx/CkXxnDNJT/FMsxd2F0I1hkAdqdQkv50/OM0PrNdDk0dFnGh3Frq1pXB
XjNAFeXmKCQrYTf+Ow2R4Ba+Hyeh6LhjZpFrzd/MdZOUJ0/wUSuw50UD2IRL8xdHIoQyNZdmKCfU
wcPACl4INrNy3myWh9bKk0iesieEnD4whKUDrvhLz6T2ZHPhS4O5pW1itjNnSGGStq/KNr5LJEGK
prN1JNUg/FbVj4UqhoLyY7lTwADhRxiL1w7WJeb5mFWXLQUl9DbXDZhadaovYLNRH9sS0KvutuSj
Cbv99RatGatRfzdHDxKMcyareck1BlK60Tqng+Il9Z05N0yrkr32SBn6gRrul5ANOd1KcxZcJvRa
I1dtNrE6+y6h8GhsPpRWww8coi/zq2aF0B1WpAwDNEo11ZNwydXmVqGFujcbRCK5QcFpE0u4wZwL
zF0syyd1ZiCZ6apK6nLC24t45RGze63DzwJs4O5+WDiz8YUOyOOWkGCCqt6W+u0EWn5Y0g/slsYu
NLFn8N3laVqRVzCuoIfgwQfQnPLkStKgPyp774PUa5x02s9H4ShWbesNDBtYK3LDWuKxGQDeu0MB
qhUNHvVKRRGUfkr5Zkw6lUtb0/0j1hRwOtt+1LuqCQrXB4Uzbz5SS1zrtBk6glILpu7hwYF4ea6u
dIpmEOB23aCPNtalP1W02+RdRu9RcfMKTipwY2PFJkFElQ5YYnjkLh28a9/B206gcr0//W2tmUKc
bguq0E726U/ugGJQ5ly9bFLTBLnMz9uYJkyCvZQdViA1BAAleHFzRkCNbW7BQ3tsLhv+n2eVAZJi
0R+lcrEARqdWoRMje7Lqyeb7aBm11HeT+WPUXRuISRdalV1XpSqjkSJopOK3AZMYa9O1Fo616VTC
SlCVxhISUoD8Da2Fn3NVTYz7n3YWeR3FCGyNbO/Wz9sbJl2eSbZAPCwO9ZDlm++zRFjaANXdTDs9
bsNcLNmxjE9rB22o24FEqmd4xzsxsvZAwFesoOK82fpMlc46IfmVUCLeXkPdxyP0f6PQpahx79at
jkE1EoSpgqTSQ/NNJReHxnvLsjZzdfM1S9+oXMQaO24egnHKEizABoMXwUmaFAv/ZYdTuH89nzup
PwpNytfg63EkijyGicloEmOD9HgtGfIsDYXaUSKKwQmtVrlunIiQ2q4j+St/TqiHYiEhbh88tH3R
gDaMa1QICqMhrLAfdp7LtREJ/DIhPTv81/AwsaAIUo7skptbkKq44ybMXKdABqzUYGiwUT63Xy7R
I+DsYGTJoo8/LTtG1s4yOANNTwc+nt2LE5vqTX0DUQiQ8/G851Q0wJXXLIhcxMgsDDfM01jVFOUD
gHZCPLOLs9qPzM9CnbRo7uyMhjog0fiRLXxocnAn3+wbmPl6UrYJn2hgmqRBFqRmVvV1/wkBxO3/
XUzdmLZtOpcxOXjV31dPm1R5/xZ/H+eagn1SKaYFJMRXRrUpYjWoKreXH0V+3XvNm7Y2LeQ/euzo
VRnIcaj8pLSST6XG9T8Sv1GlT4XFV2Y56xoX33dgFrJoNFItvJkuXvoerrcczkpf8AalPK6IE5mQ
qGPd1PTOwVs8jvf0r5I0DC+7cQAi/cEV/yEmoQHLA8qTbpxFKo8DmU5wAvxUvKX8lQIS38+OM0/N
sMlNPPoE1Rs++T4czsrs+Fhx0VukPHcd7dT9RmkekJWiZYLdlVk/E433zbO5Aom5HUbzX3gfG9tH
Hjrs1FJYJQs/IOYdjMAVAlBTE8Yw9gqBJHd0M9eGibKTcWWYdNlP8OtuHVkjzYZVkkvhV/WXOwOj
OERNLHc34MDZAd9FQUYrRc9AURKyLQQEC72upOvgexq9bCjaq/whcBWwDb2oMobaO1S9VfCPjIa9
Hvh7lZbtkR4fbhxRuHI1qzzjEMCpSWAAJoev1pOWuZB2n1gHiLVKWlOGsroMfv5hOkyt2VuglhXB
NRa9X2xfJgJtdgMyNwHNFsDK7iu9icoPHuc75DdtgH9/wPGQystvJIKxW3rwZm484u1iDPCGPPKM
YGZmfv5sOdPozNqcfGkIb8i7UO4cs42B4uZwMW1IbwOl+Z8kHElJXZWj4yD9M4p6diYPCpUdzqSD
TS8UBjiLrt6balXtKXKp2TP/aY1AEiHI3yk5SR1r96MNRKOdgZNmEQixmEeUf0ddD7wUu7KI37gU
aLYzbW5fyh96ZvavHD36jRon7K0dEb1BAgNLWh/MLrOGGKpv1+Udr6BMHXm7mxyzYtl3r5jzt4BC
O3zHR3yS0MX7TeBmedKGBkgtD/dLVJhB3kjX+aFJbFILqlwVLdYDlqLGnIQRyQWEDRVmqR+h+gxl
ZHxxr0Q/npq09dM7Ky1jENgUXxwPfSPUkiNl/FWeJGxS+uQq9FXDWpHXgWVYuWELgSaWOoZiemdl
dUynb9pJc8ENWilEzuG5uz9e49xuP4gcRU/gYtDec5flN0BpvOUIKPj6BLlByz2+n/Aoe3iDKRyE
FoJ1zjy7QRf52W60kwBEDcTupbQT4yRMSfSCFJeMZJUW/NZoodCsUmix3hUV5bt7gjf98JkE/Npi
V2GiWfoM2ybEHjxo2Bm/JSixdMSO8R19lsK16bQF5w21kcIKFQLLgXOF0r6zG2eYr7Dxjs6yfXcJ
QlhODb3Hs/vjCPReE9vXwWpwBk0lvyfjWmOjPQoWI9U0AmgNwWpz2SlNwydns9KSi15X2JL3VWYy
Sc4AM7My9brXwYNVATYUER3eJ0xgqHmrAcEmf2bwPm+m8/1krCFhUh0PKMrmMoZTA87ir27AkMMt
5pPi9XQYfsiileE1vSq+y/rUuCi13UUW+B8oBEFtgl0Hyb6iWPoqkUgIpxNVDnH7K25NJOLdyia4
weLAnBbzF1mE9u60SUZxjlZUAizIc3/tuqWSOs6njHAG+oUFT2f2m/23jtkaLuRWzksyRq01Fdex
P2b+U8ZEBRhUwQx0gqGPNh2LCP+cqGKYbigF0ksZVET/GImHjfMgxEE8R85nAwJaffJ3grKUKGoh
d1j90KePwIPgX1fmhq/WA67b30j6zKjcTxfapVwRIrU5SgQE0yYAg2ecfnFKyFDWjIY6/xDAM1Z/
hgngAHvGxHWO0L+ookwmK767Krm+4ofvcJaucw4Jdygutn6ngpuQKGHW0uuSLxmG+4Tn+4BfZwzC
eKz/8zp/bX+svrfD63tpyOpXKSrfUVICzX3qlc9NKflQb7DL4pcwPwvkaafisdfbNGFyxSzizLi4
i6mG72Usz3Y+AyKuD1V9J1v8r5zF+srNQ6AX9v6nQKQm/nePaEmbuqlhedmA30cFwQOWoAYx9iKm
Y9VCQnEvqQrRE3M9g1A5LNMyAIMsLgrlpVD92elReJdyF4LCY1NxIHpuLQwyZ00YSEYDCiEEGhh4
np6g4QTviSjgx6jO0Q8Q3f/uXtUQlG7dkAgftfNRxEkkRCu5unT1MYGqYNnaoAejgRpjRTH0sWl3
Nl/GwdmT8Em5KNdccyifUSqLK6lQFFp+yeO9dnycIeWJ/s4mr5lug9vyBNb+o2C/aLE2D8EFaFMY
Q6+sWjI1NDawJEVHNwzJjp5zVdF8tzCVR7UOvRSs7L3QEZ8nilXylwhzp2QmUrnrDB3dn3QBM/vV
d6892Db+ScpjyIIPwfkGPIBYHQIA8zRzKmlmmKfDAcSEemS5u3YLbEpCVBWqGYs9PBkXfYIr8yrI
2XXiv45s13XNnX2GySYZQeoMhTGBKTDoyVmsDirxQhtdvSAU0DBhcHHH9sBKAOBkzfD+DliLlFR5
7YJBdlmylWaDJX8JrZnSpfZWU7dOsM7qmBUqyPnQpRfu8xSBAJJAJvi3znqGImqLYonrYAK5zO4h
LoOIPCVNv1GbluIRH5oezRJhQ/ukIjJ4Mp6rhtBWn5wUurKQgWUB1IfudMuTz3NQfPkUuvTiIEjp
NPH9DvJnnmGQKDoBb5fhL45+UH0LgvJGZ0xvd0JneNxp2LOjxf9JAaYKhIPyZBl7zkPHPC2tP6Ae
ljYBXQ8moKzCFTK/4P4j59slBv4C8ZWg74u97HoqllMGGbOSUbvZz6XJH6YmtWAgLKLHRxdAp5AT
QtqsdjCBS70vMZKKRP2mkfaDuJePZrK6TFcIcGMIyijUe/ddlfsL5LCWYN0vj89ptbv59iGCM/Zt
KHExbfLzgazt68QKzF//CcenBk1xoLPU2rGXmJppdiJIjsVmmFY2lEoB9w89tQ4LOmEWn5goJIDA
y79BSK5QRUaswxUan3ZV/NyOfCLmydz0zi/4jjfNXg47Cid2OdMrM9kQB+AueBrB6C30UaoaL9nM
DpYAws1rJKtyYzVPbp0GI3eP9DkOFgqgJCfSk8140HGLBGmZ4nudEEQV0rG3Cf8S5iJ5SMH4c6c8
i3OFx+GZUfmltW7N8ZX+tAgQyAeofThD1LLpIKcYaqDEYyjGr2MN/frbgn3ZDlCuRoEuSgC3qqdH
wsegLDDYIaLZC0NsRU9kWrk1KRsDw4izjNnye5QVo+3gV3hggT+I7mUWniELf1nb58wU0vIwIQRj
9/NvjdQwN7VWgsvD9lXmfqMM+oPIjbNL1dN4feZG7XtWTYkvK5gcJF/KCxeYc/sG+pIZ5aKIrMSc
ltcygChVq0HO4hnRgRCdVbjVk/6/dbVYYf+f+jNR4CBvwdNVnVQqas9HaHsCniC3Tw6f9oYqLqw6
bQCKHxwfr/Un1yh8C07jwBVYQv5xwp6UmxjG9CP8+pQ0WTjYkAH8axOJcwGEc3jRMTgqyEudzZ7G
avN8ijmVPbXzPBLBo39K6UBRzacRCsKPiZtpGqdgQ2LddAJDHJgwQTUlXbnEg5ZXxbFcA2LLfywF
xPu5HdNh4kd47UCJxR/H12zhbEUSSYEtFpTCmckvNHenODntdbmfyZO2c4EkDp0y0G0MxFE+SBd0
sM5rvGe+E+qUASQkKdL37TnaBMSbnCp5suXsUXDNFdqrtYW/6Pw247wHwZuCwSCAPjfpSnbrAXEG
2EDnKnk/8gIE6YaUSsp0NMtIlF8uasp5wGZ9mN4IFzekjl4W4lZnqxvNEVpOG3bhm+dpE0C4VpNq
U3tQeO82oK3jgmknvghFpTXaxMqQOyy5p96UAOzFTQkUAzHbQ32aOi2BHEiQ3432qofYtA+dlsh3
sF+dDY5OWPYQcf6+dQPcn5suO7YbQ9cqih2NdEQNX/JLb9ofhwtpvkQZp7efyQXGlvUU2DdAkDrU
PZ2aETMX6Lz+d9HFHJLj5Il5+TSodFGaPZ89bpyLPDeyzYEhzI4I5FJyFbYsRUcs0djjKT6LUqds
gtbiybSLMSPsN33Xu7CzZj2EpR0+nIwUxvzK6f08+7lpj9CY2GaA/9lebgkNVqifgfn1oLiYSEcy
ii2yFalR+m5ZFyh6wM0ce7XEVQibky81W3ZpoR2tn3Vm28gc+AuDuJri7r18oeeuP/hc34aJ/yQ4
D+ZVA5wKncU/J4kUvXfQfTWmUIsG7TkHjcRM1FLlK3xhvXmpSkofqWapu/u9HCEDWlMfLIZNkgNh
NHhJmt+v34eWCzBbQLk5otj7Y9v2N+iEPpsFADb4CwL0jsOGwPu0K/cz+OhtBgWSPXazaDwKJF+M
x2UrCKCqjXAPXKoLUgHz/W0E6SWnponacP0GEt3DWCBpoJeDlUzYEb/6T+p66JpsfLdsWXdwKuQn
mASmj6HMfe2TuhGLETADhZ3f8PdXXnu8H7LzhOYH582OTyKt80NS3bIUpLFK+UxmUWAQdhjlfIL+
HPzs7oWCF/qEP9z9tOS7gk0PJL6ilPN7QDF2P3Mawr1digdv9hEcsgfJqqT6Svx/aR0G0tZ+O7vx
9YNi9YLvFRUUo78Xf559+182rj4yy8qmx4EkY2ZMIE7LFFwPedccFIuIDr1Sh9o0i7uD+pipcuup
XzIuS2A9G3Ic+4UO0RZo7r0N8rxQta03jKwCrHHnc2ouyJFB5YD8ubOpUCyvIa63fiiIjR8xQAmJ
zSd3eiiamh+XZbaLnYKpMIfx3RyKXTs92fHcRpOPcmh4EeMQvfn3O4gB3b5bpCtgk+QGmLkCQR+f
TnBKtU+BI3iR34OJ8gbZ1Zxcqppp1xkDU5AlrPCzmSxSz6uP8hgLOxMEM17fa48wpOz5di/4RrjH
kLc6yAutWw28X+WROMrkCqiN10AAzUEs/6SavfbmQgCzz6USrHpEL6EHyiO/DFrpNUlbfF/cjoHM
JjkPg2bXgcvsY40iERotHaBc8DWEhWxXxnW/9ciNyp9yrzS4DOSWw2EmTpGX+Df2hgvZZgiLj+Vj
d7fpdoeFmiQ7MMg0PJRypv1YoebXVxXhOw8fw2Czg1pzIL/puHG88pkuNdrYC1FOcA5/xNNxGe6X
of2JqBJUcTZb2zmTI0kBZhe32f0QYhtiI/5KmY8qcLWzOS/wGAJcW72SSzIWDAKQ9Mq8A8GE5CgO
kfvn8PAn2cEuPhhx62+gp3Hu5ctC9tIwoaTUjS9t2VvAizZC9StwGhkawdeUtir+YXrxcGb/Xlq3
sRX17wxcem0fyuMhHstah3g5UWSCsyuDLIBfftePIVYnP+41UgmwB5CghSefECPwrL2xlInSceyI
dJhVUIH8VYUmXtOo9S4rNGA1SxEyKPb2tRyvbIPrbCp4PvfZEzyuEYgxBBSl63rvLHq7+uaEpZ7N
t0jUqM5UdBoPuTmlQ7vD/AvGN+WLfsQxAsO7wYYFuGtZLJ2acIsZtZxR4lwvUyv+MlD9n+uRr7/Q
E9ilZStmL6bbCckts5OUyHNwjy7aNK3k8V7LfxIXowIKHgvNzOlUqqiTNnknVOorp4oO2/qs/uxf
z4OS6ej2t3FmpjG6ZzkX6IYzJzc8PAybFk0lw0DxFEj8UAG7LYbEDEaB8ngTFMMfWuS2wP3Cksf2
OZspBrHAvPcdbUb2RP4SLPuiPMFXrxCHznVb4BOHQdlDXxEjwqltdGUIF2x5EPAs+Q5ELXROsfY5
2dEM5zM5YVqnrgLd2mg62E5nsGfkdFko15JcQWaoSgt+caeocPT6ynoKglW5Xhbo9FkcSUzruoeH
OsaRlBgitJfdLeCDBGK8fvNPWk3a6c4lBf3ob4gdSXLSzk9zSuocys2Kns/WpRDjQL/e+pG0lYeV
PzjlcuMPOfvwQvfUO0njlp4AI2C4ETloDt4UvsNvlqSQsvbRzzcr+bXui+s0539151kX2at53+yr
WttRJCvpY2qW7NXQdayqp/F2NdVERMrvUHTfzIfNLB2SQEGQ6GF9rU16uO52lOVoTuL3pSvSQdyE
T77SKETOs7X+IAbgKb/dY8jC1wYjmjpztQ4tsEiusXMsTsYkCsUJYZQoXjLVH2FHq4asnKrVBUZZ
mozWy/0LyDahnF86SHPSIT4/w9Kd5WIi8QyYRmFnvjmFqzSVezRlrFWPDFQ0MyE/fU9ZGfuQSVr4
1ODahTrZQSCbeMTPv+o0mNINQ/jWNil6IZJzZNEXSUhoOXcayxdD9sZjxIQMd9LEaGJsoAcaAH9V
qqMPvoWr2EysyOK4tU9qteRRAuOdRDiUxSyZeHffVzbfsy/BG5sVnFiC4PX2xArufj0aAUZRt3iI
rIXrivu4Q51lRlVGV4h8h3KIsirw1PmKvMthxNxHFdY3C6C1eXs4JDJvHLQ/4p3r8vaVG8vFb9ci
J558C1AbkGudln+LDkOb0QTQ7upKo7KWHXyenqNvVwOM4r7rCBqGpWPrCBZ4CEl6p7FPnjSlSBOc
nwDWfbwWJU55btdZ2epv/+/pH5R+84g6F5L7xNgJQj64psba2mdP1XBAqDVPCdvZHYbyS+P/lAUo
H+uMSw8Nec6QrRYeD5ZhJzIM9Fm16C7+feDg4xWRxSHaizs9qgQ9ej1aYK6NVzENCahN4q69sSgs
8lWKlyXeI9uEhpTBZmS3YhOhaPAyHQhDAWGrxZlfNU0RNCf175/xUwfGg5Hp364nVpdbtnpHghYg
fxHcqjhMKIJ+QZJnhZlBcfioymBdUs3ddePS+U0A4ksawHc6NRAM4gRdvh4+87895PH4xUvaDR6y
0XurPzJ99U/jtcMeHWTNNk6PNZCgv7Vfdlp/jApcaCRMUhg5Lr0ArLZCajLL0RoVkSQcCMmgikDy
dLZKH2Zxp9MLZ2H1HtIcqEUsma6C+wQ8BV7CfBsxG1q6fMJHvybgj34/wYkD28lL4Ge4c0Y66OAU
JzR2vKZbaB+p0ju1HGmKaehMxA/0ykqyhoOFB9DJa/QhHJl6s9QTfgEOUxb6l9KsaTjfLis8uXXW
gnCSwgC/Dxt3GSMM7lVfNFuCj8mZTvI/qoysrPLd6DOhCkZ+wS4xR8Fl6BgMqNcg2E9Uast/I6Yi
zsP25cFhDb3DGIvBguYR1w+Q1duxj3ZttiOTes5dcvMY/LTFlKAcATJqfvIUTlSXtBGIHx4aq77D
Tx6X/xUHlqTnNSBGV9fKjHzO9x4UAeIwwUI2jEA70UyoISP7lfcZWjiVOia8YEoFaENm8y+A6C/6
5gGGhZzDm38ycftk1sI9U7nDPgYzL130QS0+qOBh/+VxYslr9+XVvhOIKoggzwAlzzmj8M6PU8rN
a94mBbRB61ki/u8sJK1HDOBQYBGnw74R/w7C9Qkb6YeY2m5ZSCjknNDt6MitwO+3mzKETrfgcQAb
L3i0tAC5fIgogT3YvW3tGyJ7nTrS5fJhb4rGsLuVoMX1gz5cKLYtMgcrdLtSG9JiksY82/H8SHQ4
cUx+YAtqHLioCSo+yzsEFlMOC3CFSTQsToQNjKihsEcJ+uIpe6JUh4Zjb5BoycvkzXn41+2lSYyn
uEPq4R7Go4Mn41TpUBjmyaPYLDEZBTdUGkqx5fwlBsYqh99Aq4MaB+z7AIQAiLP+DLasT8cViQRR
eYrhYytsVMRzmKA/ePqr6JwAltWgQ5VyzDd0S2wCXNuPRjsM5atSa67RU1dTTO1TUCXx4tN4t5Kh
NgvqmiddgxHfwABJidXC2pFDvXKwOFDqJYIU/1vLTumW76viOj9G5ZYzYZnrFzXfr63VBFpDAjVS
Ve2N2ybKU+vBtDzdQ8QdDPNbzffAMjDXQH4dJfTUFPNMNKtjfS81H0F4LjKgyok7/DTkmhOnd0Qm
+UZPZHOb+kHdS95rGcrqAnjx09VPf+6uBuoCHpa7qPGeyy+IgojjN8adRTlMGf7eGfvUF6mpvLNj
hu2e5LrziSExSH6O+3s7pifOYCIaloYrCSbHQR3W+wlMLUwsK1R1YbYTnx2B2XiA9pGomLeo1MF7
QGfV720rELplEsWobB0sY3lr8NoPD74EBnDGVAxSnqCXx2nAXOFO+wK2lc3lfrGss9WVrhQE3CrH
SGYIsQBkZmsoEA8Vm3Z3g83jx0sZ7ogrIO829NzNq0f4BYVH5h67DA4TpyPH4Hx9m26XdZlRJxJq
/fZNvdYyzdBfsktpY5ROJwTc4YtbAsfRltI2SPoul4pDbLZSg7ykfL42eYTxLpwIlkYS7CasvWgP
+43myLmtXvxzvYqomVuQPSBeDUYpxJ1XcqTlPkLtJ8Y/85ervNikCf+QH5EjB04+HMqXZmtRs/J/
jWlAI43B6UyedYmUDr7PC2VAYH/68tYpn5kH1q77Kkzb6VGm9ONPr/eem/Vio+fGtGzSRSCu8R/p
ivNQxDt6r6DxKPvzF1hsCSxeXl9UBwW6A29Egx4lTWgFQpBhd3UERL0PNLr6wcl5hVryH0dH8dBu
Lzkky0A9lTCU6J2xEilWmoTcwR8dNBRKzCnAy/o/e58ZF8wSSE/cT3EWIO5v6qsd9Q5X6Ez7AJkI
T+IvVbqO5HknfMYLS8eWAMeDP0CU5Sq/ASaQY9fKPpP8LW0SMCwMXmpF9flf99bFeYEo9J/5QfTf
00ELw4dWCR09D/RHh35DiUYblOIzJ91EBdRwra09GMfcm0itt27BosjOy5U40h80TfGFvdUzBhdc
pwmVV3o8FXIZMCfAfzRr89DEa+AtiEFEQg7moMQVkiBUBQRRw95dtRYvirTlc+83HCzZlCtWwziQ
QUlqH1XFQE/5fyETVyUoYHJ03b0m3lHFdaQZVYrER7qRVxS1k4quZPlBnqHZJkjgvTUotvgBC44L
4totry26Y4hKkBoRfdjoTxwqYVwCqdryrVEHbwafO8jAhC2cjwHBvJmT2J9A3iXbeB0MCKmsMYkM
RbH7fQ52lLYPkqKkWoynTf3rqo/hCDLEg6pY4DogHklmpVlrYyvr2q4ODKLXDGYGRrCBJLJYmmp8
lILvUrJdU+xPZQ7hLBCobny0BAr0tph6BkscxkjpjdC5ThQUpD3ReYQuYVlWoQuwIflo4sHM5J6R
4USTsFJdU9+FW5CkW3yDBdkW2/5ymU6ESNsaJxHg6xrgZX8aWPbN0/wOLM3qpG0R+80IirZbbO8V
m7BEtFR1gaV9dz6gXlQb+m65stFUec5Kt8kWeR/RQFyZ6LQam9UcYA6Bv9CQ3+JvfdQir6PoQGgM
fWrPrqwMJHlficZcU9+AnH4wticf3sHDTfVyUIFxnl7YSSoEfOo6pKFnk2nDpmfx4PCqm9EEsdW1
lHRFYNFu13GUryI6UNv8fRXTeTZm/zeG08f8phbjwyvZKiUxc/I1v3tYZFA2ED7+fUnQ16cdkE4S
kUt7HAapex4xD42eQE5UCSdEj++vGur7ojFvRfFMBG7LyIT8P+ZSoRkIXIrCCfKDJF2h5/sACx6a
TSvUHTbe4KowKy4pH7Qe+cNceN3gfOTGH4Y232MX83YpmjioqxQ/R/ovSqYDrk/rzIJPSx0mz+Vp
GgQHidymnuvH/ZIrjlnPVZCjR9lS/5pr9z7966ZFpzovbXmGLncUPuUzcBzdriQjCHWZYl9wIwlc
htVbs9lcHfGD3FwofqwhVt4ySQoHtrmd+RAFwo4bvJ3a7XplbJcDyrjlZigc+lKokMJk4O5DcVVd
xQTSHv3+1+5tV5CYnqbbNyLMFe7gRA/vWfCL25r9Y1x4jgYIDrXV+mkgTXI9+bKNqJh7h5ICK8pE
RwYNUPsAyR+M3d1a8SFcH8MOZG5eThrK6YD5VXWNhuICPZKNmqHpU6PC4kMTO6f9ovATAXw/AqgO
CL7SfhTtW4YElPdh8rnXVoSyY8y4Nvw8BwNY8vT8syXeWi9GuKkYxa/RojOMCEO/qZMTYrM6Z0ye
TclullY8EQ8m51u9245GMYLC/WEmjCdnHVrK42ASY0Vy0adWccZQbXAKQYwcIY+91Y2CEPDf07/b
h3yX8555IAAVFcUvVoivD9iKcgDL9Al7WRDyjzSD2NNcGVmTvx4I0etnMuPm+WA0x/uSzjNNuorY
QjzohMw5RFWti0DW8mMkuoF9WpqpFd7GrhhM+E9WLLqbsrEdHZrQDhG1D3jZILAVHKfntMqeeDH8
kmdSjXdKH1wyAQUqfryexZQbfegGX2TXxY5XrBT3PpZwL+dX6WogsT4ElNkT+iyJin8D+P9L91qT
xZoGJ+WdgHSAMPLiQSZfHtKcYs7kiR47ODOY0MjzHhUzmvejcd30lC67KnXrnFcYi+aAbtePNB6H
FvvifEcmwwRHFqWNqY5VABHhl+do4YuOKnaXqzCbSYUY36SYnb5bddRgCEjafqSgr1Ke1OkrUn7y
huwy36/HkSvwq8qvH5wVb8lgCbGQquiiDEmlyDwvSidELx/SPAjDFJ9aNtc8LRuWK+fXU4BMMEKM
ltOs47dPfk3/FVWMfkEuQiW7AGuAiU3nrDQDgVtQmRALEbJYj/nfLduoAnhhynyrXDX0v84q26Xi
+UYyB4nMb/2L7TUOuL3mRJtXhB8FgzC6OeFfisKNC5TKnQPSpplCMQH4crZ6UHlWoUAyJnRVc1ue
s4LH/Rp4vM2A62vrN2z5xLYZUfzFYJOct8AaiVu/XwguqeByxiLYQ6wF3rNnDCxg+0dTefwmbUrS
N6RJuWEOdkRv86jDkCUP1KrJ5cgnpQSYHhjJvQ7lXqCJEwaw28nEBEKvCCydJ2TFDBFffczxpVX0
BpXFHKfP+9dAdidfnRrNziUv+2BRGdc0FgYpIZLsyZSG+wL4MZg21QZEMuPYh4+XLFqdtGepzJNj
BdUgkVfjitMORkbLxgb9kmPEmInfgac/vvOYl6qbyE80JsAGVbeMnYgEvmDQ/Bt7D9wJYFBz1PQT
QarzZNThPN1tI/S9ughLLuPNGyBv4+I+Pt0bysqYWs+K6lomHulrRktT9TYKFIqDF7IOByQYhf+j
NBLTLP2MiwWKRtiyWjU3DT9ceKnkbWVm46bM2wRaqvsWAja2qvG2QiO9D6+STHQHxKJSM+ba15IN
54fEkBnkM65q0HG0YphiNQPKP14WRdRXKT+T2SU+0yQ7hPOH0LIy2s0TWdp8+hgS6ixKBdfVaP3J
ULRGYNztvPlMDYZ89tIn2vvuhOUl+yP0acuKGVuTdiue0wOqv/ZaUx1pSqLJfsvqJrgclEYZ+rZz
4fMhxO6T8hFXBGK2FsoKvGJqCKujp6qegQSw+K7TtDmwosJfzDOyGuchayXy/T22IDS6QOjfSOea
yFoCtYgiNxrXTdJ5IguMu5yy+22G+qIiCZrV2MlsP5XCkmiO7rOajqElec4PigvFGu3KFATXlX53
gzvb/hnZh5TPgvFW8+zINVTttV9xxymdWiD17Ju1EVMf/ukl7qiYtmhaOCX/MhzLTWhAQupdOvhg
O4XKIGuNj7bjkF+ZnJHTUT4TtlfV994+LQ/FQ2g0Dqnk55+vYctwsdnum1U5uUOqoqdrA0lxN5gw
mimMeQr9R1jHnao04f+UCI5ICvJEMHfcLluzCTiJooE42HJS3KlVbwcylmRvONLmMsFApI4+eiCs
huxpPqdxEvfDHxrQ71fBiu+1YCSQKAKQ0wn05ux+jq8sWQPT+NTRUqT5Sf0XyX2OxkOV2T6yrrKz
IFH3TgSh5nvbSSS56uLARsincqcM4+Rb/mn7Ly88VE0aSztB60IliPGm1rKLQC9kJsrT/Cv29ait
76rEBr+eUtOTqcPjcJcdHQJ8m6qJ4/oUAuO7EJVxbRasxZiw3D7ltlkLONxqzC+F8UpakNERwhbL
nZQ2XUJ9Iq5DAZkp49DKBWApMBo+2PNA8fmeHhwT9+2zevJYx0MmoCkrJQLYdisYvFBAcM9IxWif
oA9yf1tB21QynpY12plSwKukfwhBDAkRLznwTKCaz68jr4Qto83lps4OEzx32KT8ILqML3vL3Tmp
MavjdLY8eh8AXHBPoqI3SqtqJZ97NviC18EFM7cYc8c8SyRgcXwcMq3RQlXk1FRB7GNvZuHMvzsa
WZFG2zxzDUPbggv2wAspPk5xbcIlSVt7FUl0Xq4pwnKQLaAY+5FMuI4M36ObLPnnvp2oqlb8/V01
sdAjxKLpVzksxmvxQXbXiWB/R/hmw/xt/IgBoLgp7u3KH2X6YKOLq6FH0Gi1lhMyQU1vUNcbk5W2
th11tm+Nve8Z6PfHBQeyV7faePJCRVbaMVU6Eq6N/xwcCxzuVbjgJXJa6scSgmXdZGlcMkTCd+8w
581mxul1onY/FQT33tvovwNrwDggHTjO1g5kAB5my9cO2SzhClmpWySW3sl6TdQnxEU7XdJY6Vi8
MFM/5AH6gEt368EAiWsciNjXG2+XM2ZLp4Xnary4P377mxsTpD5eHugL2pi1yVVd2PKqRRAhyKDV
iBe7CfQgQfDhUOzTIMpb/WQl7nAwMbOScEXq8nQXSKPoLv6UKTMBUgSKWyBalBxtUb0pTQggozTS
A0+aAhoJdSUN5NkwZ9Jx/JbolqolhlRK62eYQ+svCrxTwjon3YE+IQiI0knV9YJ6o8T/ttz7hk/W
S2gvqtuPETGRUlYcbRdsqAr6ve1anj244JYfslNcNro7g7LGaUg9QxOkmKpwZj4kr4dN5bquzT6f
ojZtxpCjMb7vNJDiXi2ZnqT5qmieKDl8/D4VGI+Tyu8yTgfxvhGv0/BiyISsNLQN33HXvDPvocyX
yWpMUiZwlplUzjyVdNeMktVYW7TNiPlT43XP+gH2vuv+tRrt2hEgfnH6+iVvCy41MkIhbem3SasR
/bVqePwAMcaleg/2eGtOXO8t8wJ+I7TWKNUHpa+o6eJw0mvhReWQ8RkZN5jLjl/jE/stArHO/qPd
s0I+CQ9BkfjHhPuLrsnfU2h00f37BHSGCPO87Cawu/60jBAWTCxXVLtCVyA1n71u1fp5X/oFJu3N
pOgI7MDuyB6ZFjZtVcGLS98TNICooHHVoNZxkmCmyxEbx2ty5fwgG6gZle63PCkr7oasJhqfdGWD
wEgzu6Z8EET95WvXpnEAY3q5f9SMiL79pIV6pzJNRlh4qu/EKO9UOFo0MKrlSEGQ+rmNZ8c5geiR
9akLXBWfMY4OjBuVFL102ZP3i3VY4MqfNHBh6mtc/WZAUOtauSN8cNw9a8sGSBM6HDYv0u+l3/b5
iDiccycRhijEy5hqndMXb/IVnKLrDxWCTWRTQrkwk3h/oKe8uqLp3j016Pj+wvYh1o3iK0rpKsjf
me9Nffw1Dq/iokKnpxNx3Gbrwkz+4Bo+k31QnZnvxNDXAtXUYDBIWwBwCvjbo3Vxf7Qn82c2kWhB
e1IhizpLe+b6sZi68qWwGa7eIZtbb3ZqeuHLgBgScG0e2YEZwiyc37nHVrJ2aZow7Za3rpO2TdYQ
aqRGsjXQQs6A0KL5CEJAIN8OjGfzGVxtLY5xo1eCEC0qZelZVJGRoZMzdwd0J63CJ9x/QW46DfGz
Rd3qf7gHVQVwdbUDJltlbjXqOUudToRqwmUPuRU1x52i1tIjf+vAiGFvDMHHbEybMSrNleGefPoF
rtMUgs0Ogwv2L3ZJwPhU2wE0mKqCBxwnuXTINY48g7nwv5nGecq3WlROu1At0/Nl18fnNmeVmXcu
FbmwboQZ0ebscSfzUth98bQmjhAr/rsagpWbTSDdUqkX/pazdQkCxzzeuTDMcdhPNDN1AYDDeMSt
MBE6C3g50Bl2YfYV+fKUaRyvRaS+zGiWNioHfbKQf6c8l7EWtAjo3SYRVtDITn6kk0pN4TQ0BK7o
4n80V27PTsftf6aneRDvEe9v3O9iJ60shMJmWRzCW1vj19OeOu5/KdBAbmJGIaZK5Pu3r5bK11za
xeo/gtxzUMVSHdV3NMlxHt3e7Dbrdypvzg/nr5sTuPT6d9xiCvUq1rfLIXN1YlocEX+UDAUcEwO7
pCw8Dy6Za/KqmTHYdIB/Bluwh5j8lNwBF4LIoLO9PftNq6TRXWjYZch+C9t9dmTVgqQuQ+QFcMfz
JxWtwE80j1y4nU6/dPO9/oyJMMF5w6SwgTAlyxdYmMMForWhOM/u9zjG3OunMzhzVGnck4oY/9tc
XQpHFVr3QzT7Cj6V4YdD8a1R1bCOjU47LhAU1yecHBNg5IvkYr3kPVa0G6sYy8M49XeIGytz0EGw
7RavIw8xyT2kL/CUgvt18jzIQpMOVsK0A+++CM2z40d+X6dD70yjZEc06WQriarc6qF2di7bzu6H
8pxVlHHulPctzAZan5jcw9NPsgHorYuTmoYlAyrFW3cGBDjYORk1GThmoaFjECCYmFacZngyMNBD
uD1tSwZr8q4FAtEIYOqoEBxhMPzVocc2hxj7sty7IKMPXVrzIAVNfmuDRr+8b3msIFADYjO0QQJw
v5tYhs28/fbxLpCKt08L5SIyvhZoq+Tb9ayfrAzoYshJkMHDxX7FXugVMFWPInkMPHv3a6TiO/yC
1IJ+63ghj6CeYxz55p4zo470dgJRVeOgdsXqr5cmPF28Zu+KEOWejqcKXQjR5vJRJrrVk27h/tEP
zuTJoR7MWFShmQxBWASH0TmT/r9ST/mMTuwyLwzW5lDDcNTypHpVvhSci5qpyznRprUh3I/PYe+A
7b50istaUBijSQ/JKSJWo+8xNf/oSzW+WzKxbFGbD06qjZBBBj6YsWCQICjOC2vqoox1HNh4Lbaa
e+/oMAzfv983eMOlYxrYd05t74VvWfN8QkMSK2SmKF6P7AUYbWD5/+KBUDfIgICFNNZF1MWUBIdk
M+xdYGIqIyfLCPulJMLN73E3++2n2S9JyyMIp+vJq7sLbeZwuMFHLc3r7Z121WnhdcXrMcHIp7WD
AWbMEcQcVobrMyfzDk2g27rbPnzaangI3kpi199QhPglsz0PgKoM2ZgrEMfMYskCs7ZAGB8of0gi
LDsCEQ34k2IKIIzjtal6nhuEZC5e9fUbjZNfpJ9vyTWUZ1uUNTGEbzPP6SOKvxSaQ+v5J7W+G/Yp
g1X1NXShta2C6gQXTeG0aZ4O969QbZBbzdxPJVYKCPtJvJktkN2BDFtXGmkjo4S+Dv5YfYkZHR/H
ox1luq5xdmcWo031ZqvsaB1uBVJl8SAq6b/GMZJbi9+BVYJ5Pc+24fJS18nXqp87HMmG4XRQVvQd
Cop+3gNZW4k3pugW4O3x46q0IC0lvfd0bNOo5PgHysVzfxQyXLZtkrQGgdrLMQUk6Sb5alwUajyK
587HZT11lQo9bSzpKV1stQ+dhORzPeAxzq5o4Y313cECodMxHbni9Kq/6+hI9KdymaI3sC0Iknpa
qfO1fDN7vUgPlX42c4cemGOEJsafhUUpK+Gp9B4CPRNWJdnxBa5tgaHGPiYu9zZPoKmHYg3YXPGw
5T6UstXjcsZrEJUY/mmVrtxxT04GiWJPOm45OWdLN/wviqhnogynlWMX2rPZ3qfSW0/r+Ze9eiSR
eKgyvCs8zfNF4EYapaY1v0aWk5Ahu4Kt2FA27o5gUFxF75zABuscWRglMRlBjOg4zGxo4WSOjxyY
JodhnDehkyEw//5fucsQ+S27jdccQopd8aHw1UustQK13kC+G9k7i8t/jDPP93qKL2y89g+2ZPbb
04LJjEwqr7dQerg8eOIOyEY4ZIxGbTEgvt4GAceBH+MdIUAgw1ylQAXRfbFKAio3kb+14/OlXAEJ
yJqiS3SNsbBN7wLE+Ywl0LL8rPqy0BXoOlsL2UdkTLPCXk4Q2CBMRtmU4yIpfA8XnrXVckkqPuiG
nt6b5U2ICOYwfMrfcnaUVnD/7DLnyyNEVm28NwTDjGM/9lw5UlQVW33MtaDTsl6WmkARnhfO3dz6
dqedf44fkg3uV5BjzQGn5VV9Ee/rBqKp3z6mrVu0HUcdc7sky8Iu6geJQ5OOPgyP7H9juDCUYQ3w
yOONy9gqgLd2L24rpG391R7kcIgMUvcr380QmJFW+eESd6VQBQYFMaAHgAje23c6wlDeTn9CId51
55poyBsiaP8GSPTYZ3fwq09OvP1+w8oP5ndWlOC5cm+fBj8LIoUY2tDXFm3Q83fiLiR9U8Ec18gh
HKoU405gYaykcPCaCKts872OGkkwf9Tp7yYzQpzGCWpOFE+hwTOdnmvlEVetGlG7pZY8U35s6itg
NkMYllOHwSqVHjIbREwQO+2TQ0S4jgnicMgDZvW9x8i38nfp+AhEm/gRwoBHyFsZr/0EI8cxXSiq
Kdy9m4jKrOXCAXmL9fLJpWSkXHm2FIZAhlqQ1cowecARXUjVxYiCPO8JdZvdiHhpvcxeIpg0vU/p
NTJuza3IkAqBztJiKtqVkSqlQ1A438tD4sjff0pbUO1HCSTxDsiefSjmkZauKyKhMpHSVYZXytW9
lO8UX785iuKlXHjOCfViHWHBNYsUC7emEw6GTtUGskjNbhJePb2Dj2AtOc4h0IDYaHaBl//J4l61
HzUDYcp8NMz7qC+AJmwepfQArH9Wl0gIDd4G/2ESdXhDguwSJwzsYueAG4OaOBt0FOpTmsrQqJVq
nBdFgRkG4cnKAq3IHOApaVsVlp/P0aY/x+bMTQJWFD81H0IulDZS09iJUWWlitw0CUYhiZjEiDCC
VdxlkfecWiif4BLXtZreT1qozm3YL+6/y8qJswuB2+p3tbaukcMh/2pYQqH4ys7erM2SVzSmnlSK
ens/uF2KKPzY1WQitdKvrdc84M/5U6JJScUM4akO0TZaV5JX/IO0bo0SSM5TdpqCRvMdwnEDqVRN
Jjpmh985omEE86tjJtrYqVSNZ6RjgqMpyikApqRoDLIfe7qyxtDq8Q/PPbRH27YGTIGsam11KIM1
9uIAwktyNx1u4jArCZ1tyXMZD8BfRAbF3x6ZQIBcjZw8LJE4loT96AhX0ho1bc7OK5+8JhMX9vRK
N8LSH937/+vYJR0B3zCxC+x4enO6tDTUpc+dN69sK7MQg8FpQoPb5wrTkKncB39ry2cs88KsdEgw
kkVxTASoKXQ6EGr3yPpLXHKthgtMilAdTkrAvmRjwM7JjE/NwPrmF0pAF59Ab3o4c/bNdot5NGwN
POoq59BGWHzTW0odIDSEh6jBr65an/LS0bZcmgWq5AM6cTcCyNjTXIq4RQG9MR5gEKOIuJoqB6h1
6xDrvWSrfdAqWdS8G4vQ85ameq3swyj2kWOPykLlHJbrm27wDj+nYKWyCp6zSDW+sWG6kzs3nUh4
BQHkkvcK8kMIXwa4vnlngaLL8YQGOI19F1rtoa3Avd4YWUTzzqFuFhabMqGCG6SOg2Lu5aDIrJkM
m5i6e8/PiSi6FoYCJ7BZ8ftXvr/KoGmHgKGolMfW5v5vduNdHkt6gC2QphpiAQKzvcznTvOVHaDD
g9z0IHGiIkUPSVVpIdPyTuxI9SNospIFLmKapYCSnaBjrnBsZtwWPMbCRB8U31RHavdRAezG5HpA
jlLGXC8c3b4DS7K3vBTMrhlZKU2QVVV1wt6EORVydE7/QCahA2/clnoDiHUFaxC6Q0DIwCEY4Gmo
Ml8wbmIurfr5j0ijuDR5cmb+FZJTjCJubg7LquOsH66XH0qeRGrhoHfJ4ZsVnQo4874T75tZr9nH
+m9hilY9oK++xTXkcyt0jlkxpuOWy5EB7/ZZ/xhWbr9NLUSvxFhgCmYvprMyaTXhfQE+uyM6IP1a
dCcuP5hbISaZw7BxyAKySQU8CdJf+0Xhjx9wx5FMKtDLfKETKxdzh2sKXthoh3c4ldyPvvxflhLm
xOGiRAjszi8Vs+SYNSRVOxAusxKV8QMzmeSwb+T7EXPtMap95lI1jAi/VnDom/rp3dNIN36qSzXw
TnyAgA5/gFlIeXAQ15oZct8zFFierDphxkgJ4kr3M3vxI1vKMeQN3quDhikRFxgoDjb2++3MVtzt
FEd5ZJAADdBhz4vd7t7OB6lxFT2Nfip2y4S6/uWhHZw3E825KJivT37awBOZ5GBJwZoW1Uxu9xdh
g0UaOMIfpnHfxl4Y59hhMue1w3TqeMvEZtSnevP1ibuxUX+bn2v2ZZDIDwBTmLZg0lmGuVNHfu/h
EuODOrt5f7xiJLk8TZtxqRSD/2L2BXk0nEeWdLuKRCfuUoYRtu7t6FyNzRJlo3VrpcY0JI0ty3bR
+09r2UGPsTz5ayss+HfGq+O3JkQFKqPSLrYFlLJIzNmaXHXdDkirXksPsvJgjZ8JLAYTNIhnd0UV
Vi4+0iLHnYkZ/j6b52Mp53I7ziiouMaZfklonPxj0wnGj/NhTO+LrRr3P5Cbq5z8U/wAnld8E93F
EWVg2+DUe0qhPd6VEtSXAASCx1hfH1+joaY27grrTrw/JLJMQ2AU3UljRDoUixmqJg/KACoHXzNk
I9V0QUWo9Q2bVE5Fb6yzooMC/TtPR6/Iqzd6jhFAOqfDX55Dsau2ekjA/OWSVxQXP25tc7TRkR1L
u3oKGqf8fvOLwr1VZghNc3P0tYwT75vFZuLRQTCoIcojHVbOtTFPAsx+k+Hy9ZjNa56LquC750TV
qipH6KqMaCvAMwKgaRpcXnwVSSSFbTcL8aAXGdfNtNNUmGOUyk3CHaPloHLStFF+RmyL92kK8quo
IIegK5E0D0TRKI+TdbL8j+pi0f9krpxOsB1gmmjID0e1fsnlQEVBwjXO1ElxZib6Z1ENQQurcp0D
ppqJLTJH2aB4i9RX4x7zjjtxi/PE/K1ku5mSDGqR/N+5Ncx2MsChwMQySOLS6IuZVsshgBGTnK4r
sOEhhPVsSTSGyAWQpznkhJn+1+Wz4NpTG6NgBYFDdlwlKXetUr1fE27OVcjx1NshQTY4yV2Z4dBN
qVjN0dctxz7p23WpfvjwnahK21ZVYNYwDhMKvkNhZAaooR75XQW31SRMGN7NqEqWwWpOTnPlUkZd
kTVhfZxupPrh0fGbJiHyWUUyZXvUx/Gqp+9lOZoPSpYqbhKr0e5QRlcCYqTP3hC7ZhIPARXfbbKp
a5qg9uUig/yGSi/00T073SRhtu8K5q+Vvc1Mnf5L8kCcIg5L+MzGYY1ekapCZqeU5jDczN2LhMUu
IW4q6JKKBVBo1PA/CC+iOI90HPSz0so5Z/xSUZWcIOIqDhkKxcJX+QR5CXkcIPoGyHnt56gr9fYQ
fnctqN1QDjsKX+SAP6Bl3FnaENxM9lmjEPOh3IlTpc3J0CU6RtTa8+lNRPw/itq+vYtE+ehSqdl/
Vr/de2zheKphRJ1LOKRpJD6bSnjWT0XQ0DS9rTOB2Q9u4D9NXxzJ7p+3tmNA3H1HImoCXiPocRtl
wusKsVvzCZRN0ul7UcvGm0WINrhEoi7xtPt8EUOhnRkl0H3qjekO1aOsV25BQWjaNuNGph8DYP6/
sQYfvtMWUF+aOQoJrB2XmlqiYw5YOlozE/yrwnIXQ06qeUzpVY3R2bb54HNtpOeUZm7hcQip+ibg
0BjC8PFjPt2NWNu/41ZeYiwwF3WsgkaPFEMpZjKN8j4wj7xkNU84d6BwoW78iLU+Qk2CTPyzDjxr
bGVqox2lrmgd0oSLPZ8Z3XIxdD9KFTTyqrUu+EVzjNotpK9ikCcphHuR8KVhCxwq3EVgU0nyDUAO
8dXaW1eudmW7XyT9+YTSQG3/npdiCrajklh47FFI94/3QpOzq3D4Cz5mImHHF2b7vMxhqijufL+v
FppurJxlDTJm2MschXn+C3ZccYKPVTjFzi/AI/aWBlywAx6MmVmzgkA0yB8Y9MPm6Zmwr1EObMIC
oQ22h0hw+gcsMADOSnx5MYam0LPRoXu1zprQPdPsfM+0DZm+wmC6zOPZgCFj9XzVu0WHF3LL36sx
l6OPjKf9nUMhAoQ98+ky3ATGKX6rRU3q7xO3sgmCjE0PF2MmJOtDy4R2h5MYwJ9AfGV8vXRhTosJ
2I7SIgFDE+8LOIhyeY64+CdLHH1VKAH+mNUd0ZTiTIqQ+97BSO+dfGvUzRYy45+nETFYewd885FY
bOWJ6z/aSWWG1UKXnkBuojjjUhZeOJMA3xNNZ2eU3cdxoWdIFEMnE9H9M811C29arGXvrtocbm7b
IaCSBWbpgwafDctwl8GivlTVbr43ly/AG6kfbDVSF14X9OBwHbid82kt3SQuWsTZf+MhuRAF7uNl
PfGiSNlewr32eWYaRWVyj9XbWQjf8oPkzsyhyGfYNmcPnKtGzvu2HdKR4GE5lx2GAaH9JlOCe9XS
d18cTIwnJW8fE+B86EblWV5xqCSTP3GhdFeNntD03LkqloOsEEmqnX+2iXShLFzRya270n2FxVap
tr5tpGlEbSmwrknuckKsG5Dyi//lbl30KF09lCTTTuX7r8SVwIXSsgjQQAQLRHsA7cV0RXrrlXBm
Paxr6R7FDISGdtY/mtS4Olc242Qpnoq0YuS4oaa8/+QTmvKXdvsC83/f/y0t2pYx9FS0CN33Xi3s
uOfK9V3M5UTbo+Bg9QOvCJJEoxzrsz2yaekVlyUVOc+sCPE9cHbimZx8PQhiqEPmVdTa2LrySpB2
BxEHwrHA+6j6Cbc5bQhhB/NMXYZnFe36MmUWIO8YWnao6UlbEsJU9qNQgDtqtKItW9P6/TK9S9rN
7I9M/OKMEXgMVjaxdTO7AUqNnwDBXaZtqEEIw7jSvgufgkA1ffK9W4tNKrAWEZPhG5vuEOXsFIla
c1jx3MHdIhgo2SrS3R+/hR5u6o/lwiNE3WPTl4X28Bla6xocatadvjkT
`protect end_protected
