`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oY5wf0WWX9TmZJ6S0zmqSdysGyQUSpHhrO3uYHSsbT/3SPJV1MkWxovK6CWoZf4Hsx/8no+bh9DC
GOWQKFd3xQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DCpf50Fpo6D+nZDE0DuufMJylk1AQc+gPV1fpqvFhXKsMv1xvCP5UgMfNL0Fm5I9A878fX28Y+IE
rQjqicz0zU7oYdVlQ0WQTWGOiWON3Q1Uss2feP3lQbEIpVTI0B3v+QKFFB6hWsHyPS6/KyyQGsLz
w+EgHqC16a8wDqkEpZ8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UKzEP6VqgTWsCFk58axOjQr+0vN8abAoah1i9n8tHxDcQkIPf3TbS/oeFZeSn437we7U99Nicp1B
G8J6uywfMMUM/lmA38lvWCnjyOHgrvbLnVCeGhhHId+PGVozdAsOle5B/Zm1QijVC5eMIjM00Mck
6A0tIHQ976Tl+CU+ZD/klqYjT0V4qP5K0JVK6IewU4Eg6wNHJWDuJdFMPLLGQmwk7BVpSeZG3/Zz
Trskdl2qcBE+aG/W5ivz8xgcG8vxWJ0sWequwRmaw0gBBEv6Il6V82cQcEjCemDIWoswlggzQR7z
0IIAHpObzStT/t9//lg6r2lnob2G0o/YKDDlFQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xuFaXI00isIavxltw8bYz15xYSGDD5xZIJ+QnG+BrZce+MyDA56rxkrHyj6cecEhrUiijJFr1Ljd
mJqxbnZDTRyVLR1aEd1blZji+q0ABi606bV2PY/eDVJztlQgdKWqU7v8imTnSTFFNcqbsa6H0D5a
2tLeuK/kgGR+DVe25hs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VqGAq2kVIbSpn9FUtgdAhOfJmfNxQ3ZC5nIVSOgN8SyaueMaNpm4bXCLdDSWYJw/+INp68HGY345
hMAqnGQObmw7Tp49btnaZS0kwP+RjOHHJ4ru3J0OhoPl0j/RR5+VUHOuq7dqJ1HZ5Kdpfur8Gc/h
AMrvDUnk9ThH8VpOJhsH2oMrN07LPbv0P0p7ehQC9NEd8qnGD8Ar2jLb73XVuHVHGt4IU96j4NJ+
XaLwbFvMbjz1Gs7yoimBbHheDTV4GHhp0IR6mqj0ccJGu6xUHWUDCDQ6Jd239hBD9T4DRQIsuktR
Pz0enByNgWmJyw+gEeGgjYFJbBEHMRxnnBKTfQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5072)
`protect data_block
N8L5lQdYG6OYemq1SzlnrXtvr8pnDuR9vyC650ZH3EDDDN8ySgozolUQP5d26yLYafhncHIWKJTM
QjNN6UAIBJsT81X5U4mksBVLprYG7km8FDZW0QXtCpdG9sgxhSeVru66VWDOU685AsoItp4msK1I
PCH+92p2Qi7fw1DCEVToizngDVQqR3ANwHtNnrbhUmti/VP20280SD3rrkIhQaMiSpUS0m7a7zOo
Zo9ecJ3Gt+wxUJb4rWkNunYUQeUDL7GTVKLjb4NpsXDRr2budPQiU2u5aJi+x5IPDaw5npgyxMq2
xnCAdzifeRmNpiJ8yCg0cDCP9tbwJIc4rL1XgBF+ifJ0tkJHYBbxA/TDXwvyb3ToEB0kr0eplHxJ
wc17R7XXZEXbHZglW34GfX5JU45KP0DSltJsfEg501D2cslOHo3gdRLnLLERG5JQ+q3jYnDADbMW
glWX8KWIHszzzjvz75dyzpmeTXZoWvv6HmYPriFXprPQxm3UT6+6qDL5w4pBtRgkpAxqT8YfDHY0
e3kwsHvT4E/KhffUhGunoW0XZKWpdqrCIwn3zdUSnqHuOCzRUNJl7Ke++rRZZxKm1QPlCnDy6yla
SAhXSfstfGtbWQNMFeg2HhFvJknb2mtALIqKT5Zxy74MYIBqfuoxDXXk5kPKdSxpRZSdGE9m6dKo
gxywvrn9TTu8NAD7xgVuL4xPFpNuOdDGF0QSEOIgB4F4VhUfsCJbqbSzKy1Q9keRO0D8MMabUn4S
YE6onAsMyT4w0yut3UeHhuM2Yvm2flo+72pv9ZFTEzwpB/8BRHHeRAHGPQCv+BGaiLucMfvLx8mF
59Sn6KVtuWlSjTb3IILuLYUyvmDQgs8fu5U4Hvwe8q7m3Wtq41Jx4uOssM6jF0hZcUNlBLIO34X4
FmOX5WR6Ld400q9qnvE9HwnxxGWRk3y1pymDCJHEbibI1WG6F9Ab2Vi10GCeBCv0QAvDzLG67LhZ
gMiXgRNjMGYA3pYKwbicU0BRSWnrEqWsqi1gxLAmVKaDdyDbhCAZjWqObTAPXiBwUsdjOAgEf+DQ
RnqeX7zOMCrXcU97qrQh6ZDyRQb4J/G1s/vHECDAo8eOztopsSnNKGhqsbuEva1bRNL1rX8WvqqU
rddT7q0MCO3T/6L7My63OdocKuZqg5lG7VyEjo4rnyxReqOu1NKKz9cdIh/6oRDoL9gdQMMGak2f
V85r1cazoOQ+8zHW56YxFI1/GSsHdlTV+dQWDDZyQ6zqA0jgcm8pEGtMpUzwHNZLiRB34dWg6BKv
5bfheQ3Enf7Se3leZgQIhpdfIz+oXK7QvHgUsaZvd/nwT6CcX5A34WRHIHgs6+5nRNODbb5xIQ7j
8rEAhyWvj1XWF+cnnrA+g1sij+gBtRprfmwD2xUQpWHQCPF3yNgDg592UQo6tYZlsgBZdlASiRY+
GZDWwi6094xsMExcNdmzmcqtxUqPpg/fPs5TR9NVxPsVTYQR9bVYJ7+x2VcP+J+hQXHOQgVCla74
OZpaLYeEtoxW4WVTLI4YbWBCMq+mziHHDeQS+dPJpkz1Mq0AXkANGq12OE4UWnSK8huidPR53mH7
ABpQHYfrkY89KW9peFDJR9g/9J+SipMMFAwGf1FQEbc0UfNtAkckRDr71v3iAP+53yHGRshCKgkj
THVTdSIKLLPP9/LD+bZ6boXTOp73brxzMteuAQIxEvkPsgYYYdIiAa2CT3ZyymFmCbTWK64bOXzG
LWDdy18Wwjg8zI0aMxs4YPwGa6ZZ/+Fc8AttUJQe0+hBa335cz9ENOCWwmS7EwxS8qGWCK47V+nD
DqK52KP6nyOZz5D1sRggfRYx1Rpn2EQYebJxJJH2ow6b+zvSIDyqG+jSEHuZ4GT+j7HGQgH6gAVg
ZXMr+j3MjDXLwApAyDhsoNjEo5izM4YUiHvXe0yIZ9CCnyA6eBxLDdXUD+8ilH5ljcCINhkcu9Zh
/67DHRRaGDvmVetTgurdNujhhW98hvhd3rCAyxRzTl02AMuinzyy4qzLQgE2XZrCjv0ZhyfpOA4N
kiN+q9hLJvWkAdGnWWo0SmM3q/K8ASPmqiMfLOhPmrxFsE2iLoJauOZ8F44bWL0Wl7f+DTPqovJL
0PvrpiCBE1SLLkhohFx+8EIKBdEF0Z0HVqJ1ARkSNUIV+P7UQjIaGv/t9sLxL23bPFhyHIYIsl88
VBNEc/zp5Dp1orp40NgfjvEKOktp/9L/mY09XXdvQaSUDUi9dq5/zp3LZA5oiGhTcwUDftMTV4Zm
kblMvO7Ty0hJ4ubjKXahXTo2lxj9TFpTjMcNkg5nOt7Pg8IteS6pO+NMg5mcn311byTP7fsPdPVd
+UpxNVRk5Lh8i173hAzgN51lpshu2vFdlGiw93xQ2SIgxqX7wbeJImublCYCM9PC/PXl9KJwHN2C
F8qwMVmIx+HKWwjHR14DUkVMQN3remwFyoAfl+VC1HpdimOju9mhN+bAFRuWtHYUfyB5MpKMDu4K
ctB6h8Zibc09sSYDl2RUHB2CwE0v9r1Wlzv+Z331+bJrXn6t7cUvz95H2d8oTiFyb7glz0b0c52m
T9LJY+gzWH7xW+fPLgIwbD86kSMPL7la1qShww2GXFOfbZrVvqB4WOff/duSKIWVDMSFw4CdlGON
EgpXBKfx8KJGlgySc394mo6guEOn7hkqA4mBA/KbGzOwqERU9kDNRRWNKKGRTqWupWDw+4oKTdFr
r6BDDn8C7o3z97fLoVBA186JS9onS5X1QkgAFTTiK8PlZiEbDxsZzaxuQcKP7QsM9Qu6Jo8Unzxz
QkPqGGVZeglfHLgTa4RMN6n1w7crc2Pp+/7PvUlrEAN679SQQzumkZvIsQCTZGA/qVcJvYie8HvJ
egcEQ7Y10AI6KQ64SQkUVANdv1xTpdQRBp2jA/gIooc/cuwS8mnVnAIsJPLbB88+WGsNPnrfq/Eo
0E5FwnitxjaXczu8H0Eqfrv5l/wID+tti4CTDgvvN3EO6fsfaxWGTuPZj5hglK8RIFExV4JXyLDX
g4W6ZvFFsXWw5w1XYH7u/03IxRBe+xwyc23uBQSZ2rVRVFdEnL2nt6CSmCVl6bfdKgCk/bCJpOap
0bW99Yy3qyQwiF8A1xnWj+LuNDafKg3wo1KZgpNa9lRtlTNfnLonPpgeTd0NJKaUqRj84LYUknwP
62DSfn2zHpKJgKJSgKibIMKyGaTW1Bk+bVkgOg3fyWgETBzIf76rQ50XuYwz/cwv+znTS1ByKGQe
vB/CHB68BbjmRHtTbZgcC6AhellwsWHwmbRKrMSutOsMUK9bk+PK1N2XD2rCW9Kgykwd/aotaXpm
0ZJLIDHQlLH1dXcpT+ZTpn0uQp7Hsd+BhJa7yLcT45fJEEeQYdFC+lpK0PHZ/N+QEFv4QYrgSugJ
ntgO2EvP6HF/pVEMpNvaQLXa/czfUCHHh+9770gGp8Zu1DONHEk+YlayZsQONNri6Per4UqfdkKo
65D05dsyzwYy6kgEsqwJ9Ie4DG5dpA1zPI2GggYyhuMmqK1ipGCRku7omSgt9b+DuWyIMEQAOeq+
zF2oA1fKn5V0QoF/xEEaaCqTexO/33rN6f1DKMGH1qsucbWyAZkw0VGtQeEHiZk6bpRMgJee3Zeq
3+tBI/cnUIRsIwC7ouWueNkD/XFnLzFn6f4bHXt60Fsfu2o3ekzlbX2m5rMxXcAfq8mspcdflYAA
SUFtMXdSg35oH4c4NlARFcvATWkavWyetXfXCc7A6wA66vpst8qiB5e6alS8pOua1mPFjTH/Mghm
0P0udeOvMTWflWa6IXxjd2G2g+CbticFOkz+RDtAbQ4QlC8OxUjS2GeMgrsQRISM+hmEY1ZUiB+4
9kH5uM05TRNOXfrS0M05mXXLru6Bc5uQJvpeIQFUWwN1Lv+TYCAcnjc+1JHkTx4jeAD9ElNgbfqN
vAxjVGiu0CGR4PvkUm8iOCJHRvNkqBIrIBAOl3CahDhgeng3BxU3Su5APHpyjDmeGxV2pWFDh+Qa
rslZ5xO5dlkY5UWn/xAuM88Uyd7xpqQpk1lZIU+o5Nu4kSQRDd6JossTG7StYUVHuflyPT9IEK9N
CWnUUOziEIggoEg4Z7073/2hYtOfWYU81dOFuaNuoCEJUl3BB4m3JiWHCdRN2qJ5sWPpzRCGriWP
zuuCA3D35EghHDLBiSvBGUmx1d3iGe1AnLSoi0SsQW1uWUQpmKZZ38Bol48WrbJhpvK7tIuc/vBM
SEO1q6Rvq2SchjUdbIKrybJhoh1esDeRjIvLg/pF7AIvvaTB/inTMogLw/hQPo1qi8z2P/fUbsGK
lHiERGnIjasPx6DlqVqAHhcH+qGqMCVe5+FeBxrjQLYZJAqHJPtI17+OLnzWQuGqlGVpW7TuH9b1
C8qk5/ovqu7XsWgJdHBh8NuSWRZCqA5AhNT+9tsjbvnGnn8S+15fhShv56OZyMRzkNIeSKgU5CH4
b7FMkZ0gmU2MTExlmlDC2mYuXuTRqswmqUeM4zx1RouKg/FiZf9a9AmYO29BfZa96EdgVKpZ1CJm
2wNy/b7DtGkHFFQHdO86g2ciXtvVnDOTq7Ue3y8fZVc8+OnF+e3Zz2EYx60dJkDiLoHpUuawlWwJ
k8eRDl3Q7oXf/0ZqXKfZKfC37zlQWPWHwYoUjOvUGyNM1rBZ6wYdOtGjQ23qB4n9vRLCl2sj4Ccy
i7Zxh5SNGyRagqgeLZG6g8P0BvapmgBm+bKV4mSVqNkIgrv1j8c1p62bBinWM2WIB+BQAnoPVu68
G/ZqU0cs1zzyjvuwHqbYLe9PbmIZf04mn0J+l9/V6L83UaGsZmYSoa1Prg62fUcjlpT7ztbqPJXr
jepUo+GUzKtklPy9SN4vsEBI3uF/a60r/SZ6yJnQdl0QtODLj0wSMQ4UeGYDX1Qy1ZxQoBQ7yXWN
HqCsZVfAnjm72tbVpaCEqI2zyEjrtTsf/1p5ahCXJMYyumzvtABYH84v+APluDNrj33ejbOVEHG+
u7ouURI5UvZ93jDtJ2Vj+m5IrLgHS2UgNLdy6GxLIZ7RpnVXoK4xJfBrKkZXvWE1sueBrGcIsmr/
whHm1cb5Bb7OwXBDQE9ba9n6s7kpzdqlnOkdkqdCHEE90XkCtQFw+cLKe9fUIQe/sIh32iAD4d47
J8klRXK8C2Vwu1fKe2prJBjFWKgpLDvo03bLJvFPGpkNzgbeAfy5pf/k3MzIpvztm3TRUU7ztiiP
sLGfTUq/gt3/OoihqiaQ5zuvLzp1ZTX/tEG80buCar8ads84kcg4UvSld2MxKBTr5+210O4+qkxr
9FEsJFoE3M623NUXEtXRKGzgYxMJw7ALfr6BeKWH5E0uMv8tbTvnwxaazVjKU0P1uIJEuqplj1YP
nHuz3h2FOeMJyXNfHtUhsPknV5Yt9z+6gCF9XvjMxGsgKLYRT/6PyebyHcG2/tr2OucJpGa+nbSn
gTDiZrluTrNHA1Ipvr/6mglucEVIPfvYHb/jmGIBe/gVHvtQ9TkG6dYOdfheImzaAeKyI46Sz2hV
68h+he7SjQeJJxNuoR58fh40LUpz+qk3hXwlKhTfOfeg9lQ8PGs13hvXnbUb+htNu+5X/suHJjDw
wpuAIYdiSp01S69lPbvVJHnHJjnN31Vi55FHocMKAGNLDARyRveHrfjZxwu+2wMlpI0J6acnE3QH
sUQenft7sWRruEirelEw5giAqJu6EzEbdUe/pEX5d2Cs1jZof5d7nygy6X/7OJOXY0HwestI64Ho
0lztl+RxxVfZ5jRjTA2Lsl9lUQ3hx+TK1P6xagqZyktkCygoR/8cQvBGJ+LUD/BVIv/krnBTsTcc
QxLQJI6N/NUghvgE23K1/6G2EfbGLeTUEdrKvFPL7Bv3m1T+8MxiuAp1NhDHEPsPW6cK/U8NXb22
sQ3IoCeDc82uRoAhcbFObPaEHGpPOtAdoqFj7/qyYqNBblN2oaBIHxj+tPmg3RThr+364J40XFEu
3KGbLiYRLu5VVWdhCkvadm/J7eJeMo+QOV/G2tyqQiyS8TKe9LBiEVGBHZCShi5Z0MOkBz+j0Erj
JyAUqtTTMnwil3wXLBLiPRRZ5E7PbTvEwZPZUP+L2+KzG/m2CNGGdblNjij+h6pLO+/PdvUh/yaH
NRxkSQ+gF38+jM37XzWffLv8lClx+L6zu5mzeUBexw008YOfN7VSS2VtVtbTM2j5C1wZH0Zl0np6
RRljUXlUSzyRuz2KHIvE7PWxbfgb6icxrsQsF5a3i8cS0i8tsWD536L+wC+PFHqkywWUjeMaWQEy
N17QuSGcsnIrAYo7IeVEJ8F5QYcDuYslGwwsRuGN68eYm+Q7jtvZB1viZYDEZjxIYT/LSdQc5G6X
Wmx2BWWbuxEMvrE93d2wXx09Irl+AXbB76n0VV3imUDuINH4uyChtHi3B74Yz3Kbr0ijk0h5KdD9
i85XUo2XtXljfrWJbbNUmMIHLlxGj/+3qQLwvmXCeuYEUrZrQohcHQ3lnexk/gZCbRa2BM1CfyfO
TxSs1LDIWKqSo1uMXh5wKjJ+ab7/hK+q/LHVhxT88/qQZZKa5N7UE/V+95lk+nGNaVgw1263sm6S
woQ3XcOyAReIQpA1DP4wUhkty0koMJlj7HwDKd0qEQ0o7H9fMhKPr4U4NKaKJlPqdx2n3caZQBuB
OXU9KFISD8GL9JPIung9P8VsCzisf465qRmPdl9K6xigGnrqbx6ip04ZUWdMsOYAHvrU1lPhiMU=
`protect end_protected
