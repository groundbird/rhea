`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SBfzr4OG+Kss92GDhB+efubXS5uCzjiib40cGZlEFPDPNT+pOpfhMHbdHG1nbFM9wtj+9CQrtkcD
h/8niKwehQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mt/Lj8iu8VFQwXx95kTY7IBLbVHL9MBZeQUGRd/H+QQFpEC8iEvYdwuls/JnSMmhOJ2iG5c6Aay2
u1AeM+iLROD5Swu4Me+XK0dNgExJRPxxJVAavNlLZ0uhtWo8VYBTjvIPrVm4lD/13tPSa84YIMlb
64IZtXVHxlZ1xtgwhDw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JCLsIFfMYTZz0usUN8rJQKev+ydw+fxgYmK+qep0Wl8QpcdmqbvncpBh7rLw4TELgLWM72+RX+Cu
IWh2h87v3hLIw6LmzAQFs3pjrL/0oB1BXefzEQJeeg/c2TQCWNKiYvOzwmNesJQoo8gxzTjOc2vR
AQzWmuJ1lN1kT7rnF6pB2QdNiQLE24OI+tsuorPg9wUb3tgYLmQMPMt0LVvXWIo7jDuIMeMc/vgY
igu4wk2k3ml5YgtywiuQrDiCJWGH+CgGvip8VcJjDM8KZvl7shMcsH5B19/0FCqZFx4jBCVThVvX
5k0pvmikEwgIRU2DfqHnZ0stWzvXcwTm1ZMPjg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FBNdP+IxBwXtudukAN/KtNbUgLpqhNXYu79lLsOAhlaSkQCJgurztMExZBUZHDvMED9UZio2mu51
WlDl5iYNVX0dfqy4tuChJN95xCdto10XoznCsoayXc5ve3WiekjTQgULj8ldunSD3AAK8twCgP9q
iFHJ+EY9e4UGgCq0Pbc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gsuz/gMQPMDdtXyFHgCwtnMRQ+kML7JVa6S0X0TJd/CnW+9xdzZNfBrWdxHj6SwNwuzJwJzhNOOA
3pM9d+Mi9ZxN3f87dGEigB6Qmi8E2ql7SWoHZsLJK7TjgaSz91SHKvnP5M447Xhu+bJTkJwPdqAN
0twRElEXyfYC4XFxQYiBqsDv2CAc/FE2T0hZ5ZkQXCwudML9MSj0DmEfqMD7YIkHbL+39Anw37eG
fPXi99Lmxn+yqIGLwMq/lF4tajdPXAXPrdrihJrTU8MTm/76qUl8Ix/r5fL9tL7ONg1iN+cqKNNr
CAvu3g2+kH26lv/2+EGOeOkPGWRS0UhajpqYiA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
Fmz+ILi3ywuy2TrYL5y9scZiSDg2ftbRP31Zvf5oj6bWemEX7lYO0EiJ3IIF+9KI+CzYq1VRqBuj
VLBggUub4A1TFNzOkNW1HuVwTxoZco4+2zjd9Y6J8ggAwaL79rjdRbZD+siIb+cdg58CFrQIVhiZ
UCMdDrQU7qXFRxcB8/mfSHv2Qob3hswWIIQMAdNj9O+vDNxLYaY+y4y5QZbmVw44Egz42MIACOL7
tVFTCb5eLQQMt9CeuQTHmhECAgHaNWzeJW/xL/9O6YJo+xUQVU/rrrEm04ConicWfVQ/5WlhtRZQ
n/g0zaE3WR+Tr+K/3+I4iqoqe0KmfvYc09hWAxFViYYBrEtVVN18KPYSwpfvF52IWWa2wPXdmd/J
uOhYsR98uisNZsj5xLlSNdrkRS50yWNsA2ojFSpjJhlqYlR6+T6di09Zs7viN7Fw6afaYB/+ceAg
f4u6oI48T4LUJ0TvOUwppjEqlXiubEbhuBUgR0poLZLK6xmAmd9NnSqWnbJN9ITlJL32w7qdv780
vsO1cjrxhFklX5h2t2Jrpuj+8GMF4lDIpkt1xHHWVBSuVnbN7Ww9+yu7XrbKj/E+9SsdfTOZf80g
qtVzLvyJEWUeFTcfeLyOPPJ550XSTqWWIc84hq+g3VCN2TamR5G3WEF0yG2eXYMPjqisuI98eM89
xgm0oF0rSa7rdNthN5Jssf5CDa//SXY3Ku9glsTKXNzkYXeFIb/ag8r7fLstCksuvxsI6TW8D20e
/+d019WDaIR3udaOi6S55+kUpFb6X8MpegewQNlQnrJUeuTUgwgr5I87E6prdXmc8STkeVKJ9tYj
uH/I6aH8wVEbYL0v/h5D+sjpRA5uUXmYNfALdJxUOz5xG1xDaMU1as696ixXthfOR1xDhg90YFi0
42/m5S0LsMoHh1Q3vGGEfkLhfFinYNGj+AkspawqZKT3WRrQsVluhvgvWZ8qIirW3SaO+JLRfAI0
k7fiW3LVqIxHivJ30Lsye9QyhWtYPpK1bd4X3ScHw6LBzJV6iDe3ynzPm3vBLo+vczMjd01zw6Iy
5sFD21wWDqInUhp+gJOyBxheu6rf3iaVxBxuWh9zLDnyN5uzeN1X2StmYRuqoopjQl8mnTVBk7Lj
E/DuZpxGzuvFS2L2EcFlk1BUFkOiGZt6Qxr26X7av+17afFa0dJrY+rSYM6vojbmsoNdm8GrTacn
KaaXeuWFCfTeFDnpxHBRVq738b7PNNps1i7krlfYRxunYLTzS8WGS0wraaaYBZukM1IkQA/C6q6g
4u32ZknBQJK37icavKrBwjZ8kO4r0++ymA9B42GTk/6DQRjXlx3OsCfh1MCKtl+0mlN8eZw+UDCL
D0yIbC/PW6disr8LJPw4oNEDj3A6z3rFuEz8jxJiBJeH69z8pjHC4WusXeX0MRzo7hNe/WtpZePj
R2BTBQLrnn7CVq5eP+tpIyTmMZ+SBwGNPKJamSHT3CLqX0wrCBjvVFi5jZOZSdM9OtMOEyCE7AGR
WQRMpMUmofFWlQJgtsvYhmPQP7f1+gUp3vs2vwwsLKGUKBkQWpMKXE0QdmYX9VGHQL3374eW1kfh
Ye5YrtLX31Hx5LHY1/X3RFS6ewx05t3WJqXlWfi4f0bDCwc0B2B91xZk4GkKP7zT7lrphA87B/S5
dwgi1fWcgMoaKPrUXfLcMOyDLwufeCKQKiS4nw5mTlMhTf1GFoYjRg7GB6YTUs8icGC4DTuFfqOZ
DC5aQU36iNmGTN3DX9Oy1FGwj4xh0ct8HBiVd4pTGszKlGxtsEU58PG7htHmAv/l6F0yeSECD2IU
59pwpZLaETUfMinRxvFLsgxvZ3Xo2Hc86ackUnhOsKgiYToYABbq+oIi7U8KM/e9oRT0yifVbd4P
F02WGhokMuObHfEElby9cbjrlEUIyWAd08tDEJgiStdputOo27bxv4D/767xHGktNkxVt7sCUwqH
ipO3d89Ay+8Fx5qbAnuKjlW5LhPvnZny6GJ4VAKWwFhmrFaKyMCZY4preJttZBFQ0ML3wgMbbMpa
nNpvIyA7whJ39GIC/GtL0RhfWuWkEVbeFRLithjcaM0klfPhYMyLgIiStOAu9DD1/80OFjLSMDNa
xAMWn+Eg8nHbVDeJXMosGiJ0weDYr2ipu8RPOHQEjcJG1QD0BNIaAPf6apxoa/lhiCzoWEeLvCSi
w6+HAvtPBZkAY5cdZ7wi2iuoqXfuHDFzJV8VXr0HCOkCBlzIRjbwIoB3WGnGFqn+DFNNeCT277q4
nWaq/Z/c8lwSukmSUf+R8Lo0756P3qOpOTovCTsmy++NUVzuw+CNvI2cQ9neiqFefmCxYnAhdwQa
uHDwlUfznxr1JAkXiU/unxU2AQ7XiceEBkGiZc6kSeVFheACABb9hTN30yvr3PeFbfigmMXRjZPW
G0+6W1nFWncfw/qgHHiFswQd2lkkEmdfKJYOQHhfEkZY0AYz7oV74jikz7gZaUT3KThWOPNBYOzF
0sS4z08XSKZc1ePFuCzg6ngC+o+bWh8zD+3V2GOlN2UX+LpczzUOTNMi+o2D9l0ZP4srZKTJumdx
uDag/2q9a9g5lahtlz/0fB0xKKp5uSECQ4iAHX6F3r+eRtXE9QguH7t4h+vImigLKlpOrhFeVC48
3vpebTB49CdWSJHEgowtNCWxmu/odyNBy7dmBBVFh+3RGAKrRQ65xaH7CCxwQCjJqRHRb5ZO9ipB
vzUAnVM9mTTazTWdkQU+EBvFGbuzK2bSxDvHbQl6YD+j+NVH8f7Ez5e6oNhh0UKqQnQH1z47JFKT
5gDPM2dxPuygPNPRUqtY1uDViUnxIk/60rWGEfbXMH7jVKEGyRz6GWKtSvXjHpsOCXPRm1Lh33Jt
zafN6Tqqy1Vlg0M5EzyzhX1JzOJZ4Ylv2GgFE0KKnDaoFEM1dUmZ+gb4rmGiTSxBhffTMuUgSGo5
ZRGgD3zwW2Q9GTgR0PRQs2eQwK6U4AEh3Gvi3hNLKxrXzoG/T17TTuJOD5orkBSyiEbFjVhALGVG
gSkf/3mnV0FSB2ghjzeyGjm/n8PuxLqh5Q3PrDVvTJGDEC8VtDSk+U0qCp8v/k7Ml6zXYHCrUaLr
bAW3Eod6SlZu3EZ+inV1H6fHX4nkJObI3ZODS/L34mmNahpI2ikC9fCCjmiy8+gG1hHTkGNCsmmC
U6U9YBzzf2AcWgebdTUtutnLgWj8ayMsTFdz2OPIDEjsprJo5+EDfkBmSFZs8yXK8vfmXHpWw/MA
dzGueBZn52Di2NbVUyRY+kh7JbqmqGob3u+80/Ot6FedKXO+aVSMQ6UhGaskh3ROIitwDIRMTn1B
jufHS9jxO6Z4SUXuLQoGnrEHes4HFyquhbNFq+6ZQ0h47asyJsaliveh80SjVOdn89UNBkIyjjTI
xXdclMcJUfAHMu+ui/3FHP74uG+0yiHlHBrqRs/XnP+hGTxzS/V28kouO/is6nZrF2sewQfXi3To
0VolK9xwtkvK7EYFWbeNijrZITZ+oscBVrVrgLqZ072Ai9+Hwoja8Nz6/4qtkeihth1HG4tk2DTa
a8JAEFmUzCf0lcoqGUyxBRWI5HRoSiQ6wvWNCUi5lmR2QhnH0L0iav1IXj9V/gDAqaw0wky7nBMl
bPlPzVL890D6bgYT4MkDsScT0b0FojnwAKxfu4rr+ddSqjzVQo4D9+XILTSSPpFZh4Wcl1kqnef6
ekbjQEUytV2QnSrIKenWyr7uEVwhoEkDg99Ij3PsUU7fZwt/1aawe1BgwSdjmjxpRaiLJDsLwZhQ
z2PpSMUzwaQf9t1iqvZEBmMEAYSNgf5gxjZTtm6EVlUW/1ikjrc4HS/hzAmnygIvQoyVoJtP2g5e
LO7JNdyepa47xwfP83STVARiDspJtZNsfjqF7Rbm4ZpWS9n5oGuSDWHPnI98DOxi/tgxW5Yt2AhI
pSOavLkeCB3i4ZoqVI5WEDLO5Z3xKHpvXzhobzKL2YmDzZXdG/oUrfOhSWwJWYSQVtQP8gE/Te8z
a6r8fgT3MIQPXeqVaS+pUD0SEvrX0WhAYk8XB+jBQhteB7YWwpoM3qv2Y5YcRaRUibKfwqCHPv3I
uoDpiVQwfWBoCAZvY1843Vwz5UELLBxhgmt8cI7Z8x6RFe5l0gWgZMQf0eIdBS+AEcPy45cM9s5m
DjTDQpuS77In7Mvjt3lDUyavukTxnEgj3AfIIb3Ijb/Sja9o9SBQnOyBjiUkj0+hcIARdW4Uf1DX
AEEngZj6E/oX8o75Rqwd1x5LA5PkuY+BIQKDD7M9+w6s80vVoVL1xJjq0HSHSZEdlPX4kGUV5CQc
YQjMsXM2XgkNL8HUauFN8mtqZ7pKVE/UXZff1yP0lHXu+Y8P9MyLrYcdEdTGNaP5WEi2iunlICGG
qn9NTl6O7uAlgHVBVAPx+jQRdMz/fFDguE9szkZYvwyHthp++yMPuUBuRiCgvO9B0XmBijrTdcN8
hsARoNden3ntijmp4nMUiDW9wW6v8dGaPnjMGcG4HncsFHRHitCFBsKW57puHbJdyI4jBlR810+T
T5TU/1hyUEuiSi7nLy8mJyE72ecfO3rmHDzxbkEe+E8lxLCqp2kf96X+CM9b5cmt4sI7KXAFVh2Z
bUPtcKiRGU86sqWA1vpT7R+LlAv8Mmq4wcnZer9uIbz9RglJWJK6TqIDCJuMMIRdNQ9Esf2AVybP
f45CyiyLCmoohxi2yzhz2hJ42TFn0EPgRfgOaQEpigXb+2L2tWE8pFHyxJVt9zSYoPjXCLRDqdNr
cW6qxrWtGsbaNq7nZEtq0SpvzxNxTzRofcyrQOUVAT62pDk5vmWtlHoC2VGoiACodtdSD3Zt6wQb
B+zxf5MdLFotjViA/FNWl9Wh5quJf7J81+VZzCD9JNklhK88LXyV9aVIMjM0GFzaZfKNJNvqMPFl
0jv7rfUHfRSFdYEZq2KNrFeoDNQyoRbOGvDqlug6m5P8QF4mbfCDkhAXJtxSQJFjQpcW3/B7iBZs
PtHLekmpY2092qD7zeLo1GkdBLrLaFv4O7r5NDWOJooTKSunLznfIHgsEBdWRbvnG9FDWIw5WDyy
kyT6I1kkGdkRwzRwAnU6WTH8+w2cQj3a1piuG3JUu92745BbUQ6ZJBQXcG30VZHzqKiamEcehYME
5itpohxPxm29YkbM9Qho/em+AH6TDf/GN74xcvE9loNXZIMeGkXsv0E/OxUXemqv08QzgMIyacbY
tPjIVnprhgStIn2TZScUfrkl9aQnMqI63uuzpsQ2TjjepakmIV1fAm6zSDgiW6CV3Xt57GB4maOL
g9sohWkCXevBAZQiYf+NfAyQZ4vHKDvqYhndy0JZVnWv6suglRzakOHn+qkYJv30bsIKZhoH9Rc8
eZiOVLdqgGp1bLWlvwvCYBBuvZUM/lDK56zxBj/8tWGrBB85xjMA1HAGPCNvIsV2gZHgFlR89Vxi
MkSzgfCUPUvTZMqzS65MyqKc0kGo4BkuOKjARpXjeg5GaYDqJWDm3JICEyttblLEkkJzHO6xEKcR
uOQQEH9cQntjFoeydIkuDWLkFWFc6ggiQYdiPHzcBvwmuPwoP1GK30w7i/7fCZRhX8Qb3yKx+bgY
Usv6jYcKqqMQWutkFZP0N4ld74DhUvajjkOyXz0++v9Zq/B3kgZk8ArPM2wKcg54Ifk3PpWGtUBu
oEcySCumP+gjmTVpz0Xr+XH09gjCkjrphF5mfVAxqUWZ9ySyehi7xQfejH26LQPVu013qJBQtig8
AEXO4T9NcPuDTMNMQO7T+aFtOzR+FBOPtENY9XQ4Ibg7bg2XlEvcCXdeGWqYdqiWzT24lRy4Iqug
eGTniRng/BM2g7uM141vK/2+HVmwi3emOQGGz7K603r0t/jQsS/hOgmIJcmTqAIbHzekYkFvQwNB
VrPu9WrAgYU4p4sxSDiXHhWa23cdPeVgI7WL7Za1CxqD7zYNhAJaxYW+aNqgsvULmjc1HyHk5Nut
l7HkHITGbopUOsqpF59m8xGW23xhO3Ktr2IOrHhiz4I0FD5cp6RfEiceXNfCuWsvmsTYZWWmoZlq
ixbeRb6Da8dpcfMY2DM1GMBYO6jAjiaOvH8SR117/AtrHwVG4SKPotMEhrz562aKXjauaZ6LrgwI
sANDvpgGkw==
`protect end_protected
