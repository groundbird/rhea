`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HBqAuq9hcxsmTJ1jdxaQYlC3OLbKFqXfPdvxa2exmonb4bfWg3vqN/vPhykq5zqdHfzFR8CLSYLR
GRWjFJXJXw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eBOW7G0dqoQNH04o2KCJ86uBUy02mV5VeLxpOmIvdVnPCO+04igTlkp8KnBXz4gbCVk7DSTT4FET
cRo8vW/zJaEFB4RjuoSmVokclG0Rk5zeqE/Msx7AjluredU29LLJ3eE60GtcXVg6fK07EUjtADyq
XrAe8vOdfHgHwSMnUOo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HWwI0Ny37Vu0eWsjjGG7S7GO9BL8MriBXrIBTa35RxbagroL/fZkV8ZFCTJXbemrg0vQ1pqNOiHS
OywTAln97eaL04UuarJIZNQTXpZ4P3Q3odcywPvNLIZo8kEER0MI6AQQG+tcTTzUSld3HkFOJIeU
e+lahPy5Xju7OxF6S6weRWHq4RY/pWLpcYHzR+4N/qe2SbSR/egOHcjGAN+M6AGAM2+NZibTJ7Qj
Z+7fEE374CC+rSOa8qGuxEodS/SGh6YwlKg6v1l7jZy0dxDYXnxzpagz3Oo0ksLJzeQOV1XMcJNG
5c7YTvStqW7p7GyqwDVjqxfqHIu1RQR63uIGlw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4ppDYKBgxBKOi67zIfJ+WtALISLrfIDtUMoq1TIc24wRXVHuc/bQTgauSmhf+ppPpnTcwlXZaZmJ
FBwlx8JTdllzZGX/1OvdOpG8rtjvnJfeaczRSlMeAgSQUD3fPk17AAAdxDxAmMfrC3wLlDNLXLnj
UIxKu3DU41nBsT8F2cA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a9KhQp0xA7iIs/BXT2jIPm3JBzZ59SXezpDHLJSe80IHWKvCrsU7uFQJ3I9XddfuhojQKJwYpKQT
beUF21mNSi2fTFZVhnmRApunL2FG0AfkVWgbHJgbi8Z9uBGrttFmlc0MXTh6SruCvh/Hx2rLsHSP
xXQSli4FjblCTN9Gl0/U19BwpwJo+0YXtfhGC2OF0DsE/3+AXa987m0okNuAnG3fvsfeEURGHTuS
24+GKkV5ddJqXA6RHD28MF5LgRTJd0hbog/MhcvzXdubhTbHEYlNVJ7yS0IHk73rSWy472WHnxyM
KaRXTkt4eJ7837Lrz2aodRO8oWiswv9W78vTyg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4432)
`protect data_block
FD7g6DTKpLS/XWeI0qi0qiP9gYFvJadNiifnmiiAo1iU+8syGU2uA/rvVNULQHNsaVM5GwJUWT+a
IkzT3AuUHokMgw2bo3bItCUTDFj+scpcJMwjF1vhzc4mIRO5evdFVEr+8ql1pJ8A5dAJDVpgI1vg
sd6BQpDpIxVh2BRlYpWa9TLS6Ur3QPqUzuDZbyn7b0XSjaPQzaI6J8xs2hyTJ4+YBHSebjlXZJbO
U6mr1Lz08DHLuRN83gQ0U6udua9OAW2iSkDD+kqDMAbxaTSkeH2VTW0uxm9fiLTXTXxBdOIHNf9d
tET7/j0tE4NiWqchcO6QSWh2SMo4Xqz81cxFVkGZhLoqxEZq7gUTaDck253BBjo6apTy8IGegL/t
9mIGIqZ60o6UzyebyuCHiayjxeSGPfFzDH8E+58473/ODh07ZeUpqKwBZG8pZFqJ5iuQklOWNF11
uA2kb74dAFsTSMKjToUrYiqw4LZ+8gjJ6xrg/d0ou9rj9PECeYUZiWgyrkipXk8Ds0Ni69wTBKDF
4TKw4k1sFDcTFLm2QaE/YPns0myprzBrouDUXKGp/CyH2EEL9oe6GGsu7ykQxdnAzBfatW+x79FZ
/ytEhVzV1zrDoNVI6qSxhha1wydPhgbFoC6BVRnskxMCq9j3WkA9QdSxVEfvWcQUTrwh6SAXMT4d
uM44UulowbGMQ+0N3blFn7kOASX6W7qloo0sxi4JcTx531ewf6YGRU3goH1wac8STqs7iCzWsDx4
yZJAzvL2Bf0GluGgVAKxto8hfpTEu1jJKOuxT5WXPXegaxPpozw9IZsnHpmN8wYlzcehNTnUqydT
uJ29e9ZkeNYUjtDeThxNDH+aCS96CKwfLvpcM8JmvBMBB+hR+9OjB3G1RcRvoBrPN1f2qBqU1lpL
8MXU4bv746zb62Mi7y7HsJiw1JkgSXx6Sc63WT8EHvGQf9YixVhBwceHYER8cIaQ/5Gejg4UVRnn
WfYW4dhJE4N4QcvKNUD0aSwc+ZM+uWXy+aQ1GDWtY8v+TnviFkf3lovnrCW0ZRgYF1WxoDCPuApC
dw7RIkM+AlWSDbSzcXuJWnFhod1vy+5RNJA2JSyzr9dbUaUGchPwLoVGMHP8rw/Icoqzr0UHo/Kq
hscjS5gR0a90lknEION8Kg7+WnjLjybrhcesvLX/Zplpw4pRnSIWk+dfK/oWZ6d/aDBNVTsER9M8
5jeeQ1CtMzyiZuugrjRx5exfurbon7dt15KZDTnffkMHTLj38qjmCRjuzWIDI5ywaPPqB5hTvK2t
8s2ZirqaYJg//hO4zHc/0LzMYcSE6lNE9c2ojuhqWvhs0+QDQhXUzXElW4hYLrDSgV8+mnu7b8BP
gOtymc/1YO8DYmRxvupAYk/iS2siFl47GgD3qWzvb1grFxy1DRPZGjawqXQ9KGkemWQMbBb7AOm8
JYhZQibFpW/E1f+mlZReOzBJON7Tvbv1kUnBTx83Slh+tbn2Kp3pPap6ekKSjhwXyRf0EHhX9rk0
kKNUfUIj55aBdTFimoWbxPvlekPbqcSBlsMiUdjoTwC9UpAz3vDPideV49H67ZyA2zEF8h7wpxG6
EnllbWN43TMCaJ+rzUin+ejCsmudA/uIRuNvnt2HDnRTYhu0u8ilS950MruQpSCnSR/NTaT4v5DR
Wb0uINzbgvWHYtE6/oqmfcchMfpE4c0JGvbCX56xUX2MzV+JvU4R2ZlTvP/CFhcZiqEiFLIFpxWZ
Cu4PeJqvBRhVHI7Tj/xrxaFwFfNsE55A5m9cx7WDD3mo2XSeq5BVn8hJBmKZOUPUlFyDBMnUBfoh
PDzeBO40Q/x5cR9WAJ5OZsAZeYybGO+S+xT6iHUXYbwOKKQ5JDiiU/Lw3i6F5SH3tlj6JC0WAtqw
AFVyUIqPcG9Zj+zCjqRJKOia9jrRJ/cfOTPbzilgbRihuYpi+689c4gXTZXE88iVVMaxkmsXk59o
l1CKxIHmj38/A7Q+ccrzZjVR+Jr/AYHKZdYZmkx0imncP9TptXjOaYiqnrK2c3RGPQgUlsERvs+c
7OXhT0PQXAVb1MorFDdVjv7ylN1PbFsAndOb4i/0y2Eq1LTZG4Zg4wW7iGbfBZxM10nDQ9/kOoW5
GArh6RNboesN2Kuotvpj7jJuSnw37nBpjd2Gwsq3dVlIfolxpRrmNZHmyf22hMBz+m9Fcb8WV6XS
boI/CRfd0I2pkwKgeySnTYP8lDeRzX3ItK9r5aHDY93l0WKPaVg+/VG1dWQGxD0m+CL3X7GZhFAo
vx8YItwpQnU8b2gZFhEb7NzVcsGrfvhVXEnQ35r2vrdZ3m/R5rMKWHVcUvk0ykEJv5QAMBhIDsLu
7uKCjKlFJXiLmUipsuS2hwuLHu6+WhJh1jL5HVCPkvy9w+uGG9qQociTORl8vcNZbU2y+vi7ntdl
Lxc++8dTtpnJI585ui5mH2h0DmfJFdKBWpUTHA5EgAoS9wF9MJGtzgk4NxVNPU5zd62uPzArOayi
qFo0+RoYUrdGSVq70f8qf5sBAXHUosr67rgCdxAsZwrqmT+L9IQt3gVbuMhfwpfFgww0AGBBV2Jh
TC2JSR19Hdv4UNe/jP7I+Tnbl1d3Cbe43SmB5qcd67ad+kIkOxE7qDon/jhREJlhu4HNUQiK+M36
3eHF/sngdjg8xRpmk2k2IBWmV10XkOb8w8oiOosJN2KxG9OhDER/rz1tm+relaZ8ZEReIJJjDXKF
qu7JMlHWfiWfaJuIhhbrchG3zrSbuXs3DY94Lu8fCKw/SekmgBHFxooDXoPVriUlCfWK3eii+sqN
Q+bMDoxDy/Cbco8gVCaMeAYvFUp7z8inh92qdIWWVV9sjwcXsXEFYMywotHCQQSNPvLkxXwxWElw
1AwSQD7zEtR0FTEtV6dJ7MKrEoVWCNgBGptR0zyhWUQLIFMCAiMvQIWfHS7LFhcmbAgvKBTRC1n8
YxFQ/aZPycS7Lf35iElUMskR/Ye3Mjl1uFDfIgxpGmFn9RBgYLd/Rild0gzKwQs1wDrjKD8h77xJ
9sq93GbH9Yo912EWuwlIVATZKs8+BIuF7Fkn7pfM1pU0nCz41q3vIM8YEi0lFgrEOm4YWqZ1ev8/
KqoBIPc6ZrzGRt3rjiP1gnYaCnHt6JWFhx1nlBO8e33s4kGJpJ3da7cZ8wSGQH9jFrAenteWc0g6
nyHhFsFPqsCtnNJSX4LujFNMgT/EpeqqRkrx4WTs5pMSUb8sBPo6dvFsTqg3s/AYhaxnS19o2wWm
6AS5k/DDmvff/YtR3A0YKFbg3n8kkTjiOibs9yqq72lqIhYbKN450zsBdW1v06y7vUnIWyHOjjSt
TG0a142XBZPUJ4/jNGC8ye4Eq1qX5mmFiEi8uhxPzH5N14tm0wvGipfuJXHk0HKrxnLeBO/+adpG
XGW71nrSqfuPVxrGHwKnNw66PTjdeAnGyGKeAxha294zTAC1CEzuAmVlMzXQJAqN+0Bi2dYsk0jn
a4tX6MFAHTV5NrPnV6vuh5Y0T+eCH8nD2zzoujrLponEUatPhhBBVSXQ/aHeLZCWAnz6SeVjq5PG
hqX/MAthZCFtQArm56K+v6C+Hnwxt8OLbFdJd+KZPt9U/PazcIGnAg84NNZAb2zpldChpk9Xs1L6
ez7tfvRtIrehSWnoiXIOW0pk8rT2LZLBom4Qy0auxyE02l7G/Jm1cfntK67Kp0QKTB1gFlZwAzFx
2oQmfWvvEnujbpumbyDHLmL1dMNX7DMdv/RcjHAhmP3v2mmyzWdwV23wUVdGK9hfLmi71JSZht0W
iXlddJEiv+3fITicvg72giTC/xEAPNyQW0RSjAx7/r55mCJPYT8j28d86nrd82aM88gOLWGv2fnf
UWcqhZx4A49xNjPMMtkXGO23hx41jetnc2ukuc+E9mkp8aWsoCXqSNH/LrwHPQiYlF7ejNqtkItq
E5CdZ/es2sCQ33o94HWiJ6bO4CvQsLkGt2MVfKVekH44JyngjfSl8/VJxSvzeKkU+pvdlHOiTmHi
daAiEIPCGN9AlNfNl24KGffHudds2Euyef54cVZYvKam0gCogVKMSF5045OwcDrKcjhXyOgco3as
6f5iy8MeDHlA9MX8N2usYaSFCl9NHVdIap8QyIvXs6wZGVjSqD6XA0qAJwoiJytwcxi8OzNc+VB0
A7xGdeVYD2srkP7vFTPEyWnI5msAEFVlYV0gf59sHgUFMgzCIBP6EmhEDIh/aT1HJs4VURjnTn55
TWawFfv3d7xopxPVFg9W3spWoYooby6+DXS1qCHqlmsP1FaT5QKCFSDM1e5A2f6s1X75tbtkCX9E
UC8NBmomdB7He8E5eULTQRKyQGvQe2Qe6+wBiJDtrO6TVENDgYA9XcZ+SDMxVl+0D1ewggbPYRNP
HfGTq6L7JCB+pd6a+W0TJ3HOMPRrbv1R106ocs5KmVymcEfISpJhNpInybK/TfPEfrpN6QiHmxHK
8cjPR69SwZ1dhW3oOCTtUvI/p5McBbr7zypvvvE0uNtqne/K0v3IOGflMgLB600HR1QUhX9fB3l5
/hpiu3r847shQeuDfUgg4/H3XTY+kjuJuofBMXFW4rv3EntZ8k7uz0ffYJsdZHLA+V6/BpuP1Bmu
cr3pi2P6p9Lbgw2yuTVlZD7wMZJpckURrbtIiaTKCeJanwSVBeQqwLpjHOnuJC3wyw7KJObscB5k
1sMVMllnnEvEUWxT/LDK7Rwgjj2Rsk8gYWx4uSzSS1Xm1/UDHXPliWiNnXv7iBP3L7pjTrARMQDU
025+oVNDZeCB96o9wr9RUI+k973TxkFSJ0diA+nEqq0z1/WnWP+UpI/vAE8boxd72d4Df892PG2R
o2c9AqSOuKxwJ19rbhavaVkGoOWEyEQQB2htqvoQKeadIpd1z3l/fNUUODkml7jqGQa5Ydlfl5wz
kcaGMVjYXtP8ys+q5zYRk2UJSZ6NldvVWnEYHDcqjCLmGKmSid1UpUTVi3q8Ylp+584T8XFSsal1
btt+TgSuQwpRx8rvLLj7+Yi49vg5psDKwQ9YTPJiMVHbYr1BnkF9ucusPnB+LHAOnBB7trGEdq90
oYEYjeN0aDSQUM13yCLKzu55Ebf5LjybKUWoMaxDv/N017deNaTtQ15XyA11P2vZm6zU4/YOWR/F
a2jIgimnjk7AOTcTZfbLvlnu+cGa8Jiv18//SyNH7Ui03S1QNuj9hgN9Zm/C2ccoLGRDibl5BcrB
KBiEQAaInBZjMrX3y1pMUv5TiYHYx+Md6jwdR+LixVu23b1aAVXSXryofDewKZWvtCSswKJYK18H
BrHQZKetoYNu56hqI+aHlOmg3In5UAmB5nPeJkP1Pv3SKMbjYkNIUphNwU8AbDF66pYaKBeAKiPc
5fVJ/1eJ5It9WLDcXFjvJdCJh8HNnVk7z72BSHtVTK0DUlQUPlwqhNHg5M9UcL/Vnl8NeSq/Bnen
6YgC1WOg23WZatE6lZgsuhVsNiCrgObEjUIZRfSQFVF4R701Etz9g0981xPJtAEcPfSkIBHyR8Cb
uulcgTFn9Uov/ylJ16TDKaY2iWrAY1NYaUUtyi07EwByhsNq+nO5Geo97XncOSyY7tidP0bqsN2J
PEk7BsbPZYdoMllbRt3tz24Q6ZHI7xe9g5q+X934ZbUVnCcA1obI91hTUolAMCTtir+s9jDUaBpz
QsZUeZ7xqpH4+o7H2eOf98l84ZaBRh+8jDu7oscEwizlqkiDfZ1spi25ATSLJA1LchKnChn8Yt3E
MWP8uyKwg/cVPw0zUKm4XfvQsFeQuof1yocDV31f61FaU2+zIXC+f1I2yx2ZaUKbi3uC40+7BlBC
x88CS5Kn+Ho/UD+ftCXYPsRzBt3lYFKMgAKlCcNbos2Xib53LpkhlQl60A==
`protect end_protected
