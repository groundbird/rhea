`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pNnfPxwufKNu/AudTnGtUZ7FDvQcQU3Xs99vw+eIbG9MZyA5oCHJpIFONkSCpe7n/3fcR0SENBuY
SBE/3xHZMw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PrKn+EX/XWkCNN9n/chnKmyhdTZAmR1tGfhTgcuDVSvcpWEMkUyOySDjtgLhrMifRnRYz01dwN87
orta1O3pBhl1t8nW9RWJaGsIRoOr+m85dINBNtk39aL9Cvmg4qeo8pY3ycVNsBHz6Nz24TKmLp1P
FxA1X5inwfn7bwn9PY4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AVLy2SfXFJOgKj9p2e5xirjKDKk2CQoXQC1AhwhkKld99YJo4xmmQtHkK4d6ulhKijeOwiT2q70x
IAzkLdpEBIjXVbUIYWHlFHcU7CKNg1eIuNABZXXYwZZFp7cEBsaW/xJT3FhhgkAfDmrPmGeh7qsJ
nN1pdhGSwpe33inSzaPoupDDy/72DVVRveir8rwVntyyDiTpL+uEX/srQdqD4/9TE8LEoDevA+XC
9kjjOZcxx8AIJSLyrYJtwml1dKv5yEpq7StYQwlCET/MgiCF5sZgY21soaoicuWkTDDi4ZmdVUpG
3cLtNyXZ9PRMlaTgCfNvSWGlkzy/5HpZco9jNw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T1dCp+M3yNsXjcXqigODAZ+wsEFeLw9F2KwaatfKJKpPr9RYXd4mg4fVfm8dTkB3IlbXfyHXq4gn
/7OEOVo3ThnqH0gxGEQgn7aHu94WfbfVLmpJSMi3ENnZk1pPLLdqXU+Ed5QvfUF7mg4498O7gpmp
TkJxvjOATzKh/dn98S8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lFzHA7Pj8zxCgUuROH/vFtNAHHQS53dfvSkVyBjhPY26IMNd9FAD6II4LvXbAcd+CMjTuEtxjWuh
C22rYe/+VuLn3aez0gp4wHSP5foGR3Yjya0pE8pggbU+UDyAeTP3Qgj7VbkXEJy3brJpbFPK5Mpa
icJ1BX/Vo9lMBEeOvkzJjohuXXePAjVn4msiLQ2Zt9ZtKhrfrDaijFeYlG5TOT78UtdzP81YRZgn
QEgZCSZKUmwIMcAYTACvduvbiklmoQItVFExzMslOWN7Tqqbmkfgoj4+NNakjb2RGOdar0z/Gwfm
bLT4vVs+td95AGOjxPhRI7R42CP5FY90HRL4xw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9856)
`protect data_block
+MzeHd33A3YU1BI0GZV/Siw5wQehncgiPgrAPFMm2woSn3TbbHlsgUKwAHkpt1uZunuAj4XHzslW
jike0wHDgiWxOIyUoyBLmaRZNcjj73tMzMAKc51Bar1c/Paw93SSG7qnsjzlgqIFamqohtrANh9A
8p3LFtUYbz6k/DuvDU4NmOysqj6j+oqhET5Ko5yaze6pDTX7gdikzFFmc99yWCWaOk6jKphgaLkm
SqgOoIJFnhi2M9WGx7HT7JUfRbFLTZQN/tA194exTyGPVa6JwtABUSFaRWNnC8RyKWXzAzxBHZLr
00xjIMGQno31zF2+xjp/wWfBpy+sYZ+wUNyev9BuVZz+zJ79IC+rucw+BITSqJGjZRhyJmaHwW7g
+oi6afLLGmHm6JbYkcyVptAhvL2nw0cAek2sA9yb2nlfJFChoklDcJVKD1j3VWqoGeXJoc3EeHmC
Hwxqd0aPq9ZROzUrdxl+xzLqMt568N+q7loYiiAVW/rKcvLrYwtKCsYl6p7OoGSPT4Jw+t5+LvDR
wGVNTRuz91Z4IkLjp/0nmNQCASVnYKE6ndFw8Db72Cxn2UcALYj4XwUQ0bZG0gcwpke2nafqUq2V
keKdTCu2BPn0CDV+Uvgs10f1bovQx+f6Pm0s7AM8WMTe4ctuUD2vBE/4lVNpl7ME0LfuMK7zU/48
nxDCLb3xVnUBqTccYJVBUJgKu6k8mHVtHPkJziD/uEG3nL/JcURwZbHZfmpDrNfRIIJOqeSdxc7f
eWHoUVFJG6857MnwJNmocgTbHPmiZ4XvOCfUhCOUL1r9SDE7AWrE0gveKgK/jWk/DaORpnDVu1Eo
HJB9js4aENb7gd44dzAoQfvOcd/Iy7SGhyaCO7tQH3saw5CF1Wa3kHmaCXfH8nKeuz+MWY4DRsnu
/jE5oao8d6I/1LAie+BtjYRVfh8pv9C6ghqp4PUQ/ZHxCg8pITFV7CiENTEt2q7PuxiT3y2sr6z5
R0h3GJrKYsbWFov9uyb1tZOvIeCG0aeAKdLLpaW/CMbsvTaNoyHkKPD8KbKGrygEJXmH3nQohsLx
oJMkIOIryxUvxE6Fz/AHVfY5+JleAZFAuMmZAaruSvorlfGsaENBWFee7H0iiUmoN6e+k3CFLb+Q
HYI6nMi3ZFbC35fkN1E6G+Dg8JpTuQc2U9uTXg2Hk809mFUWczEoWLzOq6uX7A7WbghgqZZRTJpe
Ye5igPzc19uZlMbA68/a+J9qrY4PiivcyW3B3oUGhNfQW51fZMEih11ct1ZaZEgbnWjBZoBC0Rx/
jEbCJLMi3eP4crVBNjnyAtskEKkLFZcMDLQYDIc2Kb/Oqnwf8/zvFbPkx3MKj/fpj1oaIs9RWGpj
LKEXgGSJquardi1NXA9RBwBAKk9K723sKi7GfTM2OXgfhRh1M+GR13ap+Aa9u2APMDfnYK49OBqy
pci/m+w93Bp6lZEx7gn+vObrkCm6G2083MNk0Sr+XCCSuCpWnGPCXj8nImkV21QbEEEToUDGfMIC
HatDYxc+msoQ4B4fq2olFaI3fQJq8PG37JXTyOz6nqrl3u9K2/qcCMsZ/YX0d1izm67blPun+EWl
Z+jJ8JyjSXvCHBy8oy5nwgJ8FmXOaopmBhYwgqwFo1yWl34zUXIDNGLwKyd5CaRWJAcIeFu1bO9O
7srJq9guSMg4AjecWUaTPHL9HdOXAgtTCF1qpt9R2c3vVpI5gWkCu+ilcNMu2MpgKMpN8JRmwALx
1oyeXxkQbogi3gie7LHQ9ibHvXKXWxXkYb75BNTA1hJQyy+2zzETSncNTYAnSEnGGh8xYNLJPag5
eDXIO/20LFGxxYChc0Q92/hIJwIyaKVAHEQMolKSkCYB3smffzo/bXpG65I5IgcMLheeg3u0yNJa
D1Lxz0kQWrVM7wsMHRpwZ1xt+MoS2ewctMn/Ci9Qrjm6iY/RU9oLpWYnF5i0GhCBlyXFuIDmV+HI
nEmZXGCPYZTRIs3LN6AmFQ7quXiFNQ31PRlKcSruF+upzjscoOCGQgM9QA1a07p0+NQDgVdFQ1TP
kH+CXv49SSA+CST4u+8q9hc7wITesgaJHclIiNCyxhU8FgPvfK+9nm+SCOJcNdt1K4aypkoeoNHt
Jab56iSgr3HmQUibf/YkKIp7N0IyRZl9+3udn20QMkd58NZ0MxZKe1BAiUtiEbJylOoY4ZODlS+Y
UmSkSD8C7eblHvpYNYdu2UPrN4IeS1UGGqNera5Zm4TvQAz696gdfh97I+Qar6wKt7qmeCEdUl02
eWK1ObuvYQj/l+DzgA0R74m43rxXqWLYGYNAVHq+WStVD/3RLmPnPfSrfJs9lPXmip1lyk1W7t7b
iPP+7TScFy/DbEbjKSzCbAx9cFsZb4ZEvUgDJ8uCXCPK0N+qxJuxDPsl4p0qK3HoNcBBByx+QqHs
56NmWsynFe93q2flzSy0W1BRGcwxThcloAUxyiZoeOA1q+Zd9ZfvjHw0tmGVq0YPnMpIUsPUfkbA
OGaEeS9nkqJJHCrtZ1h5usweC1x1Whaxqs9j6LFEwjkZBUJWDnStti+AzS8F7OTnfgjbUith8/uz
QNBoiWfZQbjrZtxCP2uBLQkminc+OJgLo79UwQuAelF/9x2PuIjpAWPlvnX6FnI0LqiAgNOoKBPC
qNd1jegPk5jQAvbdiySlcKL9FsnPgQiA4Ak3/S1KunfMKjCZ2t7FqOMQOR2uWkFUOlovKRk0Dr3t
wbvI8we6Q5T/ARh0GpKfZVDvPPyokN45OkQNn+yeCVq/pi+44h7t14dRiLdsKoEfy2QezEaV7dl+
JMFByCE1UEquWEuJYbJLCD3U/9G8OSDYe8VfewvT5oPHIcNVxAEKgM2hjT2wfv+AUrI/qKDUsioU
KERuDeFTnpXMUCtg0F+vP28ZVSsJ4t3oPq5D6uw40aqh30cYYEm4IRrB0UWV2K+/GeoDXTVmeqoM
WCzBaEJJoEdXmDPVpXnCARrEDsggr54geePZGNem8ektjo8s2e5obd7niEYVpK8UDEhr4CodFTeT
ELKRYr5WVIIpXzZCuf5lWq9D4njBgt47SXyXXWpr5HqhsHDmw3lVRr00HAvmz9uUNC2FaF1dNjcS
rgwc0hxLgfNDy0prpWnQ3FQJHLoHDkjsN9fM3jm3N/Z1oCsx3PCVT1j5s0+4JcnhjHYSbauTkaGo
DFCtK18IzGt/ixEISS/QWpzlhKyWlFj6jwDXIGN7er8AnzkCxSi39rZiBAjMvQ4Fszc+TaZpL8Pf
o9JXe3rGg+sISQqioiozjC8gCEJJPBxdPSbSRqke7ZtLkCQH8cVuxKbv+x7/GPac9h8VUeaHnXDj
aNmFJ5BI6p1/NLbfoIiQFJsLv+esR3VhCn2xLrkZQ+UbRa7DUs+/rtp+1jarLcdwAL4wdq3VA6MJ
MI967Jr/36fuZr7q+E/s/4qRoQy5WQ8G7idTN/Q6Tnq32/QWtryCwoYhG0T0Vz+6SRobpDMzt0To
ijVb4e0heHhV6kNAathm8D/YdSNyOdKmHITIO9YGbL0FSB7xB/BXZgq8DaVWjeuv0bMwIXSdZT62
vQSvmTjj8FWbyknNjpj4nv+qedt/o4m6t14pcmYgyhtNIa+CLEs+/9VlbpBX9JNPYNaeXzJ6A9ou
FrJ9Xjl0OfGj5iEOU1nbw6Jvn3AQtYwNMMAWE4LyMpbC+uzia6+fSyO7eRnCwgQT0TBJNcQFdtZS
AN/HZYb7LoiLM/oveuCy5caiAYxsrnrC5p0LK05Xe/ceFsWk5NyeiSm0FvCt3DeeGFuI9QfypNTK
LcY7Ud+PTWeH5OTujq4FXld+gCRtMeRf4PVSGOrtjMw8DB4rJrA3Xz6sgaLu2cA2Q/57hwA492WQ
tiDsr7tHjrt50c0anwJnROtMmGQd3qZQVPF0s7jazE4P1uDiy8NpHBG+6w065mk9KvW7UZiOfkIP
YzXPzmt++SImrVXjVFzmdbomErkmQTfGx04F4jxI9rS3rmhWlBc9wBiLnxDX8P8QOmXckW1s+YRd
P6Kovg7q0xzSCIwlm61mzyV9tuuKupSSO0Xv1ouEqj+/+xHwxOXFiEAS4d6t/8Z+73E3bwqkXtwf
TFARy12HbzUhAqNdZicy0nhHZD3SPAhMK8KPk5fhiRjvvf3rByZWYprJ3J9pV/RLs2zXPYptAjdm
X11MduWOjK4YwiU3ttXxsmX3OvQzyntsHzpouGA650r7UoxV8qJZ/1l3wjQx00akXM/hm+uGSlyi
bsnaMVJE5HU88LZ1X0T2Q+PgdoSk3dR2ILlbwuqSpp1nvb9t9kh0FqFhT+VVOiyLFbbB0xcnqC2X
1TzuDVxk5ZHH3KiqhYNalYNGzMv01rWt//mGTAuIw8uy0uLwlJfMjvBpnuPNqk/ZQelc6Tkuy5qh
qZPkENuvsGXdcHXgPet7+QxTkAiigCIOpgXlKdSFQpW5HmnAOqIPWIZjxq8Zn2G3wpGqeLeKPF71
UgEpAqOgcdrwjx5IK3vELJ/MQDDS28kjfP3EdNd/QIHpypx3fvJXcjmYUctcIoRBKXCq0pZg4GaO
R6KW7Cq95IyQF+646635/pYR/Vd/ZPD5iIQDYiUBzEp7ehHfETZUF8BvcuL54zVwhmGzzzAB09nA
iProBkOI91ipJxTY6U+SHLPNEqH8+Bl4YEpzM56/Rd23X2DryKsQLEyH60DZkTKVEtqke5nRRlQ4
ai1cfQ9mAhCx/eecgmk1vHXL/e8wF2DWdt7cssk4kJVsHgI/3YhCcaJAe5FXqIdWK/FFo/J316an
A90Mm5BcHve/4JNKzuzYJCLO7tdTqneRqV3MfuRDygjp6V5e2lvnzkmgEBgwvatjKU6RrM0NVNEx
VNCoUBAq15X4psfHKmxmVm2nWu4M8ocdkj9eFRsqvGDyTIiyj5LH9QU0bwyvy61wn8ebsakvUtaB
uE83b/Co6or+eLbCrS9y/AxwxE3I11YWas4+oDc5IGO1kuCK8s/SwJTE0whZOKEGNRyr+FLcFbQG
PK4UzYfoSRGFazR0nJ64Me56D41NxFC7uUaCB2TiJg63daoWrH2L3wBRLh+c4C2t4TZJTZ7N4Aw6
7dMfuNA4iwAtPBptQRCNGOHXfS9/pg5b6n9YM/DNF0kQzfqExUCVMzBtsQEZzvgf4CCEgzMmbcZb
r8zk54dMqNFfy7eGe584xr8zATy6c6HDBMrncSLMbwAxNVzoARTcuB0amtuW+EsyN+osLr6XNt3P
XSg8eRyTY/JMUp9PWIjM9jAihUf8lILXhB+ulJd0RdI7DuGgEIvvNvazSATHfR32pvnebeouJHrn
rZPNLGomI41RmTLMvW+mVIPTF1Yr/msZSGJEzy0dOhFO78f41vVLd4u2Gija22d7oiOc2hfWgcer
Y0k9jmc5JN5Dbh24BK1R1lVZkrY/5S6ekIMSX6gGYPQnjkTvuNVduRlC8WT5t07zZZUXgyhHlwt1
86jm+vzQeI4HrE0xSo0SqgzCUl0loRdCActz/+RDqW3FgB+bE29sjDCIFp5+Mry9e/BGSP/mBtKe
/Nk5+haFNwyba9leFagw4ZM1m1iJui6CJI3DodGh5H7Hdvz0+h87C/Fd0KIROWTW2jgicYEHWOSR
3rz5ByVsJH+zREddG3sKleBZFMKRtMEbrs6zYmo+qjhqy8Th7humXd64peOlaN/xgNY66nvkY3t/
AZ2uUp9T5ZDJfRctw0lDrWeBewMR7MYiiSq8qaUebHc5qxKSNl+IiFqKgc4dbvcuBvFH/V6iKZop
wZf0z2JxcYF22M6v3KmKd9prB9+fiypcxGs/lenemSF9nTum1sqtLB1BF1StSiPE//6sfTIAwN//
lt/4IncOMGX50Na79OE8aKQgELNt6eQhKjrdlE2YJMmnXanwPdYVIbnagnF+Ri7NiExGQLSITYYe
3J1jtBXJdRaRlysYIwi0t+vxV8c10by6Trk5l8hjnpu3b7I9PXG+9jGL92dimZ6MYXJOtuYUxLao
LcadOVAQUY/BgaDa4DqpaU9dJZqfHUhaH/9fU9ArVS2Y6NorMXvx0+KVzdq+A75dl1gjjqDey5Wr
pOERXxbioVujAFT0RJCWPeJcWRfPTRxlAVUVppeKje9scDgrFeycoiFupeV+pxyNiIxVfq4Q21n2
w1TbmsHhCHlFVH5HtYyKeZp9Kpy7NzrcQab1o/QPw2GzCBUrewh5pvhciW5yDI1KHJYDh6RT8yqg
MDpEmPbPhlRffQg5X+Gxm3FeG84vYfpeyXe7gz35nNyr94QVNpQATEI2m8uhDgji+w5f3WInK8Xj
VvYlKnUCB2UK8iQqdyYPN1yPI7pIVXp8Qvwx0r870ATyYIfFaBwHlCfO77hga+DpuRHATakh39BV
NNjPF1iU6tck1Lh00p0yu90M4lk+KRbaI/JRUlJv/LLx07MuFBcc4DIoPuCyvSRzriI9FquBJxIJ
raB9wv9Cv/qHdtdlgQCypF7q0BV+gtN2s78mwi9ls5T85tAWEoLTiBneBDHrmustzKwu877d0oy1
zQVh2bZTCn5uRmhsHGQ6+hGT4fK/10rzb9vCfWeH0J18hlFS9gSRb3tPnsdh91yAftndYZp1qME+
PUqBn7AZAvMZpVPtZQh2CXj07Pbf0FDneynVm/ryNKvLCx/YNsiEYTxNW3/427BmVkcgx1lttgFS
sNNeIsIt8Uf03Lj4NXdrHVFMcjFM+LNzfTGxRWFXV4x4boy1ELV4qfgJD7lsufrWBSmKQ42YL9LX
yB2D2wX/f6MTm8uirCJssBjlritHVqVUM2BsqE3N3Ze7TvNUw/UYQwKkEM1NONYhJJljzNEt7IDq
ppVqWJJc310Xw0bfGeIrEDeCGVh/H+FBqUIa1UBVaEODRUZ12gfNCcyos4KvpmEbGwWhSjUavq6b
xwVaLpA/Iui1w0gHZu93EtRNCeVjojpFc2Cn2ey3UWeYm7UXMmj7FiYs8AcypqBqZbRzSQY/A89M
2zissMW4PUHGlZkbxJpI/tlEGkJHEH1GSNGjEd7+k+7tXGPAdTJxbMkIks5ZzD7v3F6Ja+iqQpCJ
URd9NneHJxIMfDc255U20D29Ko/xOXDGYKDh9RpY2b6NeM8wsRQ2rPO5lpCbY/Q41tSHxbuvXXxv
6MCyETAwPEIU1lk+QMKo4ytN5Gdo9FzQJLE5rz483zvLAsfBcKt1/lCXBTz6bYUfoIjKFWJLSsYG
O8vPftQnMsVqwB6my1e9fRaopZky3pDfUIDL+zx2DsOrJx05rN/pkDFBzedkqYQKhUb9Pu43P/zv
/jWuRYm4Kv+rotgjbz9m9bcvIzl74OHIFK8p5xp3xX3WcShnQ10EzXhKfZeZckHtphBN7nTwKvEf
2k/fZKL9sKQt/Hg6gjg19NwYRb0IB4zKVtg6tnjZuYEBfKj93Nm4QlPtLJS+rBnaz3Kk9ecs3gH6
r4+cFkCI/nD3U+IHOJxRhQ2qeeqffjNRbnOXL1NpaF4WfICk9SGVHNhLwDhoozyp9SiEjiE9vbLH
/sIdfOUVdX5N7+UfW+f9sMPpFZyntrqfC0jaoeVTmUomRQtZQ2SpkPfLOfaTOXJPatYSU3M8o3h6
MkEEOMGoQ7LYB6STgMKs0cO9fD3IzFj1a52rZWViHcgG52HYlmneVrPtlCQpWhyQCRMd/GrdFRAe
WhXnCDVrGvkkH4w0aJ5yqMCMlS8l/QlcYwfhKii3Lzm5N5D+35auAWUWQfAecgFXh/DN4P3XFQ9K
U5YBVXb6VAN+J5QP3NQkpQNnm+g4mJI5Nf6OBlELP9/RSUZMflKNhJinTwSw9HkhrZoy+yMrF+Fo
tWnqPiFIxwKODxTpPXXQJtk2JRgi2v1FWM+VSLNyIQ4zPBqva0TmmtAi9nfclrvW4hrVJSV/sBAS
zPUxU5BPRrjZoEhmyXJ/TIYhzRW6OBa/uC17XMLOF9LoiTUbKYaC/MytizrLr8CzKn4DLoiWmoOP
R5ZmGwWLjThQLa0X+sycW6Bcu/CA6GKBS3E6w2oq9YrV1edlXcD7jD/VlgAd6+ardNi8lyZ/kgfZ
DE5SjrxPM0CNLLGvs7B1x49W/Y4Im+J6oVTFXPpRaJysu9NGga3WSLtJtBnb7h8Heddh7ACrLOAT
Qlo4meXly7LRy2uHCozV0jk6dYA4RDyqtIE09EOjl2hvmTmoirj/gDmWKNWB7q9/fw798oSsyzuC
GZvZUX2bgrhkBV7YDTSV/yLmO5MzLQhsaFSbdFHpauYPBNW2VWIaYaCfWv+aONwe0zmIHgIDkC5g
nd9SZLYdU7v3wAMcJkIu9FMzDbRdI23zwaqeC2CdIUhhPSoYZ29GTonzCKE1+RuRm4tGuHtQfISL
MUvNGH5hNX2wa5H7HgA3NeOgtYveITOEJOuLyiM6VSZGn1lQ0IcpNxdtYp/hHk4+oCTf6D4H3IYz
8vgpZDmtPdoZSBoW7rtoPCQa6wC5MHCCVvjYTXBN1ir/zopw1JCqILp4uzlU3qeSIXjeOVMmOp1V
Pi0HcMHYF6w4GDx8JECptu+mzJ/xgEqioKWtx5AGjo10+LqjCLwwc+Ny6LuCRMuHtilQH1PAD/1h
YWVQxNLpC6xdkQjRphsbWuC6IEXakas2p/Yp0Bp3JjuHbXYK2EJiMJfx7pgSmjVoiYpBhx5nTqDh
sWgXXjkH8jPviOJugLEI/6chlHZo6li+WWegTWZVtW9+bfXUJdEthpfTHrxQszHn4GNDd8BO2yep
411X/E/cfJ264pomJOVZ+5H0/DOAfCidccnHeDlwileY/PLISf5NdnTJLVoSt0084t0Nt4sHye8c
FN48h4Ugw8ufUx0iKTvsTr3P1AI3q30bWDtxsbFB+hdhiqY74Fob57BfX/g6Kv1pPhfpD/O4kER5
QdhV0tOVxwnMy/+wDjfqmk8QChOw6MeH+cMxWwcrAvTPp+jkbWmNbCnp6fYLYiK+p9igUr43w1fW
sN0KSOqA0Id1I19TmRfwpFJodZQzdsOInrJtC12z/5ZPi6OyTJvufrQDoqBAFKNGRcm2KCyIvEP0
qmjG2T8LPHAv5ebWkgbHrN5dnmawjYTS/b0drXiIi967hu8NDzwh3w7Cv0Np/o32ruZ4H8H55WMV
jgkIN+t5ZZ75TP2y51S7mFoKwLxKqh67vnBswOOxpZlyZDuq+psV90R49Oi78wPEQfEXHA99ebjO
1UZAOZyxvvGBhZZzwE1mJqm2LItmWZmlxR77qTwLPbQmRFqWQ2GOo5JtM6ZI7L+7SdwAkcUK5z47
MZ1vuJq2ostasb96vK6nOwJXCi2ILBuofR7i+kMxa60QEQCqZdM+KNTVjJesXg28Z7j/9+Z96l5+
T7yDMD2J8wkyGK/3Y+5LYdnpeaj6dEksQyFBHsFK3hrDh/uiJG1LcuoFYMmZCNJUYq4H9CWgeS2V
2WNnIajx3wz7fkcWR/OUoX7JZX0m4w5ObgfDeNc2J05WMK46GF0fxXndyrejuy2ckGSCaeetyc1Q
eNEOQKoajw+nOHJZcdzWdSa+RDFZloW9yv6qIomA9QOLMN9qi0Zl366OHb0EJYMgbeEHFYkondY+
JGr4sSULUJNUb3aXYSx+OtyKlQIoxBU/uPDVZo8mvQGadyZOvb9QojsUdbmjpd2Tu/9GKjiNZZPj
z4aygWBGB6KdBG+nCA0W3LGUyvNvtURYdCWQ6assAXlmqjNv6nspwZR0oJAB5W4STj16E9e+yRMB
4Uj0iivFlbUmXHIrK4mjfvGgn6H+T/7vlbbK4njQkekdcay/XhB4BPPxXtHhcnggTvBO6at94dVC
SoJa9CNbgo3jE49vgbyrLgKqhRuut+i0PD3/18nk69SERee88bWtNNXZ5PPDLmCcI2GLe85aQa3q
tRAqq4HjnnpMLVV5R+4EeSyUaN7m2HJpSl5N5EvxTxS7bCrlWrheY0tvN8leVLCMY/4XRzeMHeFO
U7gWM/k4z5LFsHTiyO+P0uMfMGmvJCQibEu3ltcBuUHM0D+NlvOyBuebozm/V1VcLeLJIdIyUuVM
eH+yarJyS2KpUGW65leHX0Joa2KK75np8rlH6ASJB/jP6vApSLKAv84zs14gjh9Bu/azNSpZuvLu
YLcOmcr5r5OqcL435uvjUccPDJSIkqQxEn4oL/NSvLLrb2CDy8mfBI6npTovUyPhYST2i4u6a5rP
jF5awQBObw2DvZCOW5xhFNKmWhDj3iXAb1SlUrW6n7UTbhLMpSgiJe/aKg7Xn7vIrdJcjOkvxYRN
fAONYoCJdkCO63A92rGmlhLZeZr1sp3rLHjxcPJ7ccXGv/fcyAOXDK1jO6eVEoHFWWYVUv9lN1jQ
OkPWw8MXt4dWYSiNviTCc74pHk+54k4gFy0uGeKT+RRgbOvJ0iE6kORcq76yVM9gmbhQAiQKPGOm
w/jVbmSA/TFolWpIxQfTok352vGItu+RaLLA6c5V17TXnsOKum5TBiRqkqlZG3RKA3SvYrFXiwzU
JlZ5yo+cr6H5F4xOSVaZTTMWlOGaR4cWVWxL8Du/G9qkHSJQltwkqEYpi8+QvhNYFErRfgjGXQpn
ZQUqHUurZ/7UHFJvcgtHsO1uIrSXzCNF7iZy7fCFGwiJ1Q11MRZTE0bgKcESzUL2GvHyDTaqcXnl
YHjw4cuHefGsdwHiUDhlTt2G1Wn25bxwqzOd0/SoB/QtXbNuWp3fgoHaXIbd+htq/1eTj1nTtC5w
dVlSeLDeGYeKYGXON4fBm+JFQ21/EbkK7InfxQ2is/xDzC4a0Hv4FVTO3uwDNQWTVAxUoj/fysrx
bVJTTLqS0crMhvSwWRmUiREKQ7EVVPVtA0ogwysD290u0UXGqBEznH7qgu1BKLZ+zkl/dw1wd/Wk
tNi475Sy2VsXEeRBmgY44OBCbvwNBB2Z2YhrZ5E3HVgk2+Jam97iO+2HH66xQ5Br/dRN3QrNSoXI
+AQlNvCW6gphl/A/Kx+MGzuEDDEKkAVNHyBVTtbWq4zGGqHAnoi1hEilaa4Bb0yMLcQpP+D1k/jB
CD1llSC7YPLSI0epIavMbgaQtLscaf71g9ZPixmzHi3hH945DB/+Ewud3JKH7V3+f9DzD+HWlQf/
RG/Tsu/jXTpEWNkPimLooFHZQD6/l6MVozfinX6tQM4sBxjdaBJV7RzIWnC2qUdJ5DgyUFxta0IG
f1KDKCxVUFDInqmYkS/0/I2HyUBbxXoWJ/Y1Kgmt2/3vlRaXDokQ5aKf5/MKR8Q1LFw0VYKv2IO2
RfejPR0yWBUFxGBgFhVM1riMRPqvR1yQcB003DZ/sAbRw5MiWc7a0MqTOUwLWiSSlqFfofNKcqTe
oIfJ6MOWOcQa8KdlsYegPhhzHQMwQVewHsGiI5Kb2gZWC9jx1BXSFVozc4PHNPbYUu9kBsIzJZeC
WstPMxvXAyDBkw93gzr6/ZDkTbtat73FrWiZgGtFE9jC8WIOOnUcSBvyqZnMvLo6zUJmU0k7ebCS
uK1VVS/l+b3gtXUF0xD1lLn6fZWH3hQ5sY+9417v6Q9vBKpPcJSURZ6YPmgwnLTRFiFju5/KziZ9
dpOuP6WvnYOBZOpvgLuClhU9FaEqRQgvf5Qb+dt8X+0LpMUVGUjIQhNG73+gpFnz+FL/i3XP+57N
sGI7RZ1ZDvVywE248/ytOxZ4NjSyayQpFRVLKZtCbnWnQipfz3DJjJa9QV+7xxTWFref9/jwLvsg
G/GmLdlPjx2u7dcdCtLgdVPz+ijZnzmSUuDS1GbmKY2uTrDf4SZOWB1aqaStM7QSdIC99qUjvS64
HCj3ddL7SU6vOiv2C0p3pIVwghpCB52HlU3a2h9iOlFtuv3Nc4zQytFFw/zCvZBNeL5Yz82kEmfR
gV3V+FcJuvrfWfyVb5FSG2kK3FQuf+ApKWzQLyuKzJourXLp1I2FbWvmr5kPKDijBXOgfBJrf8Qk
7ozRLj0nGA3x17yFSahifJ5Ebrht1nQFY+rhPgITAeCBBRyZCt/fyQ5BdxoVUS4WiV1Ej3XA78Af
MF5/B6ilQ49LNorzN+dPqmmy2BibBdUeyc1DkiYehEf2OHTEjbBNqOlmntFMyajk7vnyOtzjGkDi
aKXAgP3PNJXVYS5fyMa8+EkbkVhWe1qxWJOg4hGg3/8BYGRxZY+JfQMydqsAyastwfp/WpZasaoK
GgPsLaQWMnDCG4pEgYHC0KHpAfLr7NymRJ52o+VrsrwGyrElQvV/W4qLO3glzurMeBI+xlwNi7Ka
NPCRRlNq+tgE8ud9SMyoPNCEW6XXaa64/QWa8sR6vqOsZZf4AeVX6j49Suo35DSAxH2dwNEXq+Vr
I7uZKfAn9G7m32NKfOCTLWfV1R3xSYYGH2T4R1TwwHMB9PGuwCNF3CAD7FlbYA4b1Frpi0hGvccz
WX5C2AbDKdLF1bjn5d7mxHzpq5hsy5nRDBOq5mukIeC864Ng7gcoWVzeiG3AWrMuP88KSpVg7sbU
f9vDEF8h9Wj6SAYWpqoB/2AP5vgSGUgDrixjoSlZf/igc5Gu/e4yfOTFUVkCzDzzsXTRLRGPnZAk
zyGlarMR+5g0lQ2RWvYLSEdPJlUnhYK8l8VFWyuw5THIwMT7Ox4MM1l9yIQKcLqFh4nFfKq91gdH
vn+jeyXzkjBDcnXqm6yKskQota3B+RSS0XDgLkF/nNbtJngze4rw8ZwY9TDqVjc58ZpyMRgN2orD
9vhNrqCxhln8pLBPawLPwxPBeC62tjec6RN0SKpyyXBDdE7goFYnUxcmIFurLh1e7lFeFSR9BDPG
nBwVmyvMl8a3p3/x4XongfEcZEknA8FEg+Xof+Y+ajNxTcLhJWnAFbLuTZC6zv7ISUq+3PUcWGa+
iXgd+X+kFqP7faESVgdlAwzXtIbst0LQPc6f+JXnYPZ626xAw9vVqFoCD5I0OeEqyhtqE0nWT2y3
nCBTYG4nsT1OFpkOhbKtnTcPS3isha7kQYWw7uGhTopdf6DEvWeQPoEyEiHDbHVX0yiKIty2PWct
p4X6v6oGBoABl3nmRu0JzP4PHaYCmyBYatQ0ZNS6k/xAFbpN5vcOPAhdwnvWdiWYhY0h23mqzAti
oSopTAPKKvvsSh006wlAL3kuOz3cv5w4ABzke5Syr7XCKInHAFr9gS9m6dlm02HsHWF8iQ==
`protect end_protected
